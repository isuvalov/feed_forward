--
--  Copyright (c) 2003 Launchbird Design Systems, Inc.
--  All rights reserved.
--  
--  Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
--    Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
--    Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES,
--  INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
--  IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--  OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
--  OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--  (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--  
--  Overview:
--  
--    Cordics (COordinate Rotation DIgital Computers) are used to calculate
--    trigonometric functions and complex plane phase rotations.
--    This rotation mode cordic rotates a complex vector by the initial angle.
--    If the rotation will transition through +-PI/2 then the "flip_i" control
--    input must be set.
--  
--  Interface:
--  
--    Synchronization:
--      clock_c  : Clock input.
--      enable_i : Synchronous enable.
--      reset_i  : Synchronous reset.
--  
--    Inputs:
--      flip_i   : Set to perform initial rotation if rotation will transition through +-PI/2
--      real_i   : Initial real component (signed).
--      imag_i   : Initial imaginary component (signed).
--      angle_i  : Initial angle (modulo 2PI).
--  
--    Outputs:
--      real_o   : Resulting real component (signed).
--      imag_o   : Resulting imaginary component (signed).
--      angle_o  : Resulting angle (modulo 2PI).
--  
--  Built In Parameters:
--  
--    Cordic Mode    = Rotation
--    Vector Width   = 18
--    Angle Width    = 18
--    Cordic Stages  = 18
--  
--  Resulting Pipeline Latency is 20 clock cycles.
--  
--  
--  
--  Generated by Confluence 0.6.3  --  Launchbird Design Systems, Inc.  --  www.launchbird.com
--  
--  Build Date : Fri Aug 22 09:44:26 CDT 2003
--  
--  Interface
--  
--    Build Name    : cf_cordic_r_18_18_18
--    Clock Domains : clock_c  
--    Vector Input  : enable_i(1)
--    Vector Input  : reset_i(1)
--    Vector Input  : flip_i(1)
--    Vector Input  : real_i(18)
--    Vector Input  : imag_i(18)
--    Vector Input  : ang_i(18)
--    Vector Output : real_o(18)
--    Vector Output : imag_o(18)
--    Vector Output : ang_o(18)
--  
--  
--  

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_cordic_r_18_18_18_31;
architecture rtl of cf_cordic_r_18_18_18_31 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(16 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(18 downto 0);
signal n7 : unsigned(18 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(18 downto 0);
begin
n1 <= i1(17 downto 17);
n2 <= not n1;
n3 <= i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n4 <= n2 & n3;
n5 <= "0";
n6 <= n5 & n4;
n7 <= n6 - n9;
n8 <= n7(18 downto 18);
n9 <= "0100000000000000000";
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_30;
architecture rtl of cf_cordic_r_18_18_18_30 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(1 downto 0);
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0);
signal n17 : unsigned(17 downto 0) := "000000000000000000";
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0);
signal n22 : unsigned(17 downto 0) := "000000000000000000";
signal s23_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= n1 & n1;
n3 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3) &
  i4(2 downto 2);
n4 <= n2 & n3;
n5 <= i3 + n4;
n6 <= i3 - n4;
n7 <= n5 when s23_1 = "1" else n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n8 <= "000000000000000000";
    elsif i1 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
n9 <= not s23_1;
n10 <= i3(17 downto 17);
n11 <= n10 & n10;
n12 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2);
n13 <= n11 & n12;
n14 <= i4 + n13;
n15 <= i4 - n13;
n16 <= n14 when n9 = "1" else n15;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n17 <= "000000000000000000";
    elsif i1 = "1" then
      n17 <= n16;
    end if;
  end if;
end process;
n18 <= "000010011111101101";
n19 <= i5 + n18;
n20 <= i5 - n18;
n21 <= n19 when s23_1 = "1" else n20;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n22 <= "000000000000000000";
    elsif i1 = "1" then
      n22 <= n21;
    end if;
  end if;
end process;
s23 : cf_cordic_r_18_18_18_31 port map (i5, s23_1);
o3 <= n22;
o2 <= n17;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end entity cf_cordic_r_18_18_18_29;
architecture rtl of cf_cordic_r_18_18_18_29 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(4 downto 0);
signal n5 : unsigned(5 downto 0);
signal n6 : unsigned(6 downto 0);
signal n7 : unsigned(7 downto 0);
signal n8 : unsigned(8 downto 0);
begin
n1 <= i1 & i1;
n2 <= i1 & n1;
n3 <= i1 & n2;
n4 <= i1 & n3;
n5 <= i1 & n4;
n6 <= i1 & n5;
n7 <= i1 & n6;
n8 <= i1 & n7;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_28;
architecture rtl of cf_cordic_r_18_18_18_28 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(8 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0);
signal n15 : unsigned(17 downto 0) := "000000000000000000";
signal n16 : unsigned(17 downto 0);
signal n17 : unsigned(17 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0) := "000000000000000000";
signal s21_1 : unsigned(8 downto 0);
signal s22_1 : unsigned(8 downto 0);
signal s23_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_r_18_18_18_29;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9);
n3 <= s21_1 & n2;
n4 <= i3 + n3;
n5 <= i3 - n3;
n6 <= n4 when s23_1 = "1" else n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= not s23_1;
n9 <= i3(17 downto 17);
n10 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9);
n11 <= s22_1 & n10;
n12 <= i4 + n11;
n13 <= i4 - n11;
n14 <= n12 when n8 = "1" else n13;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n15 <= "000000000000000000";
    elsif i1 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
n16 <= "000000000001010001";
n17 <= i5 + n16;
n18 <= i5 - n16;
n19 <= n17 when s23_1 = "1" else n18;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n20 <= "000000000000000000";
    elsif i1 = "1" then
      n20 <= n19;
    end if;
  end if;
end process;
s21 : cf_cordic_r_18_18_18_29 port map (n1, s21_1);
s22 : cf_cordic_r_18_18_18_29 port map (n9, s22_1);
s23 : cf_cordic_r_18_18_18_31 port map (i5, s23_1);
o3 <= n20;
o2 <= n15;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_27 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_cordic_r_18_18_18_27;
architecture rtl of cf_cordic_r_18_18_18_27 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(10 downto 0);
signal n3 : unsigned(11 downto 0);
signal n4 : unsigned(12 downto 0);
signal n5 : unsigned(13 downto 0);
signal n6 : unsigned(14 downto 0);
signal n7 : unsigned(15 downto 0);
signal s8_1 : unsigned(8 downto 0);
component cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_r_18_18_18_29;
begin
n1 <= i1 & s8_1;
n2 <= i1 & n1;
n3 <= i1 & n2;
n4 <= i1 & n3;
n5 <= i1 & n4;
n6 <= i1 & n5;
n7 <= i1 & n6;
s8 : cf_cordic_r_18_18_18_29 port map (i1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_26;
architecture rtl of cf_cordic_r_18_18_18_26 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(16 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(16 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0);
signal n17 : unsigned(17 downto 0) := "000000000000000000";
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0);
signal n22 : unsigned(17 downto 0) := "000000000000000000";
signal s23_1 : unsigned(15 downto 0);
signal s24_1 : unsigned(15 downto 0);
signal s25_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_27 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_r_18_18_18_27;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= n1 & s23_1;
n3 <= i4(17 downto 17);
n4 <= n2 & n3;
n5 <= i3 + n4;
n6 <= i3 - n4;
n7 <= n5 when s25_1 = "1" else n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n8 <= "000000000000000000";
    elsif i1 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
n9 <= not s25_1;
n10 <= i3(17 downto 17);
n11 <= n10 & s24_1;
n12 <= i3(17 downto 17);
n13 <= n11 & n12;
n14 <= i4 + n13;
n15 <= i4 - n13;
n16 <= n14 when n9 = "1" else n15;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n17 <= "000000000000000000";
    elsif i1 = "1" then
      n17 <= n16;
    end if;
  end if;
end process;
n18 <= "000000000000000000";
n19 <= i5 + n18;
n20 <= i5 - n18;
n21 <= n19 when s25_1 = "1" else n20;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n22 <= "000000000000000000";
    elsif i1 = "1" then
      n22 <= n21;
    end if;
  end if;
end process;
s23 : cf_cordic_r_18_18_18_27 port map (n1, s23_1);
s24 : cf_cordic_r_18_18_18_27 port map (n10, s24_1);
s25 : cf_cordic_r_18_18_18_31 port map (i5, s25_1);
o3 <= n22;
o2 <= n17;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_25;
architecture rtl of cf_cordic_r_18_18_18_25 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(1 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0);
signal n15 : unsigned(17 downto 0) := "000000000000000000";
signal n16 : unsigned(17 downto 0);
signal n17 : unsigned(17 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0) := "000000000000000000";
signal s21_1 : unsigned(15 downto 0);
signal s22_1 : unsigned(15 downto 0);
signal s23_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_27 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_r_18_18_18_27;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= i4(17 downto 17) &
  i4(16 downto 16);
n3 <= s21_1 & n2;
n4 <= i3 + n3;
n5 <= i3 - n3;
n6 <= n4 when s23_1 = "1" else n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= not s23_1;
n9 <= i3(17 downto 17);
n10 <= i3(17 downto 17) &
  i3(16 downto 16);
n11 <= s22_1 & n10;
n12 <= i4 + n11;
n13 <= i4 - n11;
n14 <= n12 when n8 = "1" else n13;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n15 <= "000000000000000000";
    elsif i1 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
n16 <= "000000000000000001";
n17 <= i5 + n16;
n18 <= i5 - n16;
n19 <= n17 when s23_1 = "1" else n18;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n20 <= "000000000000000000";
    elsif i1 = "1" then
      n20 <= n19;
    end if;
  end if;
end process;
s21 : cf_cordic_r_18_18_18_27 port map (n1, s21_1);
s22 : cf_cordic_r_18_18_18_27 port map (n9, s22_1);
s23 : cf_cordic_r_18_18_18_31 port map (i5, s23_1);
o3 <= n20;
o2 <= n15;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_24 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_24;
architecture rtl of cf_cordic_r_18_18_18_24 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(12 downto 0);
signal n6 : unsigned(13 downto 0);
signal n7 : unsigned(14 downto 0);
signal n8 : unsigned(2 downto 0);
signal n9 : unsigned(17 downto 0);
signal s10_1 : unsigned(8 downto 0);
component cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_r_18_18_18_29;
begin
n1 <= i1(17 downto 17);
n2 <= n1 & s10_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= n1 & n6;
n8 <= i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15);
n9 <= n7 & n8;
s10 : cf_cordic_r_18_18_18_29 port map (n1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_23 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_23;
architecture rtl of cf_cordic_r_18_18_18_23 is
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0) := "000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0) := "000000000000000000";
signal s15_1 : unsigned(17 downto 0);
signal s16_1 : unsigned(17 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_24 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_24;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "000000000000000001";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_r_18_18_18_24 port map (i3, s15_1);
s16 : cf_cordic_r_18_18_18_24 port map (i4, s16_1);
s17 : cf_cordic_r_18_18_18_31 port map (i5, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_22 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_22;
architecture rtl of cf_cordic_r_18_18_18_22 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(12 downto 0);
signal n6 : unsigned(13 downto 0);
signal n7 : unsigned(3 downto 0);
signal n8 : unsigned(17 downto 0);
signal s9_1 : unsigned(8 downto 0);
component cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_r_18_18_18_29;
begin
n1 <= i1(17 downto 17);
n2 <= n1 & s9_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14);
n8 <= n6 & n7;
s9 : cf_cordic_r_18_18_18_29 port map (n1, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_21;
architecture rtl of cf_cordic_r_18_18_18_21 is
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0) := "000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0) := "000000000000000000";
signal s15_1 : unsigned(17 downto 0);
signal s16_1 : unsigned(17 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_22 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_22;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "000000000000000011";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_r_18_18_18_22 port map (i3, s15_1);
s16 : cf_cordic_r_18_18_18_22 port map (i4, s16_1);
s17 : cf_cordic_r_18_18_18_31 port map (i5, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_20 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_20;
architecture rtl of cf_cordic_r_18_18_18_20 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(12 downto 0);
signal n6 : unsigned(4 downto 0);
signal n7 : unsigned(17 downto 0);
signal s8_1 : unsigned(8 downto 0);
component cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_r_18_18_18_29;
begin
n1 <= i1(17 downto 17);
n2 <= n1 & s8_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13);
n7 <= n5 & n6;
s8 : cf_cordic_r_18_18_18_29 port map (n1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_19;
architecture rtl of cf_cordic_r_18_18_18_19 is
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0) := "000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0) := "000000000000000000";
signal s15_1 : unsigned(17 downto 0);
signal s16_1 : unsigned(17 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_20 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_20;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "000000000000000101";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_r_18_18_18_20 port map (i3, s15_1);
s16 : cf_cordic_r_18_18_18_20 port map (i4, s16_1);
s17 : cf_cordic_r_18_18_18_31 port map (i5, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_18;
architecture rtl of cf_cordic_r_18_18_18_18 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(5 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0);
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(9 downto 0);
signal n14 : unsigned(10 downto 0);
signal n15 : unsigned(11 downto 0);
signal n16 : unsigned(5 downto 0);
signal n17 : unsigned(17 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(17 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0);
signal n25 : unsigned(17 downto 0);
signal n26 : unsigned(17 downto 0) := "000000000000000000";
signal s27_1 : unsigned(8 downto 0);
signal s28_1 : unsigned(8 downto 0);
signal s29_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_r_18_18_18_29;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= n1 & s27_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12);
n6 <= n4 & n5;
n7 <= i3 + n6;
n8 <= i3 - n6;
n9 <= n7 when s29_1 = "1" else n8;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n10 <= "000000000000000000";
    elsif i1 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
n11 <= not s29_1;
n12 <= i3(17 downto 17);
n13 <= n12 & s28_1;
n14 <= n12 & n13;
n15 <= n12 & n14;
n16 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12);
n17 <= n15 & n16;
n18 <= i4 + n17;
n19 <= i4 - n17;
n20 <= n18 when n11 = "1" else n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n21 <= "000000000000000000";
    elsif i1 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= "000000000000001010";
n23 <= i5 + n22;
n24 <= i5 - n22;
n25 <= n23 when s29_1 = "1" else n24;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n26 <= "000000000000000000";
    elsif i1 = "1" then
      n26 <= n25;
    end if;
  end if;
end process;
s27 : cf_cordic_r_18_18_18_29 port map (n1, s27_1);
s28 : cf_cordic_r_18_18_18_29 port map (n12, s28_1);
s29 : cf_cordic_r_18_18_18_31 port map (i5, s29_1);
o3 <= n26;
o2 <= n21;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_17;
architecture rtl of cf_cordic_r_18_18_18_17 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(6 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(9 downto 0);
signal n13 : unsigned(10 downto 0);
signal n14 : unsigned(6 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0);
signal n17 : unsigned(17 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0);
signal n22 : unsigned(17 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal s25_1 : unsigned(8 downto 0);
signal s26_1 : unsigned(8 downto 0);
signal s27_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_r_18_18_18_29;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= n1 & s25_1;
n3 <= n1 & n2;
n4 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11);
n5 <= n3 & n4;
n6 <= i3 + n5;
n7 <= i3 - n5;
n8 <= n6 when s27_1 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= not s27_1;
n11 <= i3(17 downto 17);
n12 <= n11 & s26_1;
n13 <= n11 & n12;
n14 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11);
n15 <= n13 & n14;
n16 <= i4 + n15;
n17 <= i4 - n15;
n18 <= n16 when n10 = "1" else n17;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n19 <= "000000000000000000";
    elsif i1 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= "000000000000010100";
n21 <= i5 + n20;
n22 <= i5 - n20;
n23 <= n21 when s27_1 = "1" else n22;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n24 <= "000000000000000000";
    elsif i1 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
s25 : cf_cordic_r_18_18_18_29 port map (n1, s25_1);
s26 : cf_cordic_r_18_18_18_29 port map (n11, s26_1);
s27 : cf_cordic_r_18_18_18_31 port map (i5, s27_1);
o3 <= n24;
o2 <= n19;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_16;
architecture rtl of cf_cordic_r_18_18_18_16 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(9 downto 0);
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0);
signal n17 : unsigned(17 downto 0) := "000000000000000000";
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0);
signal n22 : unsigned(17 downto 0) := "000000000000000000";
signal s23_1 : unsigned(8 downto 0);
signal s24_1 : unsigned(8 downto 0);
signal s25_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_29 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_r_18_18_18_29;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= n1 & s23_1;
n3 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10);
n4 <= n2 & n3;
n5 <= i3 + n4;
n6 <= i3 - n4;
n7 <= n5 when s25_1 = "1" else n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n8 <= "000000000000000000";
    elsif i1 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
n9 <= not s25_1;
n10 <= i3(17 downto 17);
n11 <= n10 & s24_1;
n12 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10);
n13 <= n11 & n12;
n14 <= i4 + n13;
n15 <= i4 - n13;
n16 <= n14 when n9 = "1" else n15;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n17 <= "000000000000000000";
    elsif i1 = "1" then
      n17 <= n16;
    end if;
  end if;
end process;
n18 <= "000000000000101001";
n19 <= i5 + n18;
n20 <= i5 - n18;
n21 <= n19 when s25_1 = "1" else n20;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n22 <= "000000000000000000";
    elsif i1 = "1" then
      n22 <= n21;
    end if;
  end if;
end process;
s23 : cf_cordic_r_18_18_18_29 port map (n1, s23_1);
s24 : cf_cordic_r_18_18_18_29 port map (n10, s24_1);
s25 : cf_cordic_r_18_18_18_31 port map (i5, s25_1);
o3 <= n22;
o2 <= n17;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_15;
architecture rtl of cf_cordic_r_18_18_18_15 is
signal s1_1 : unsigned(17 downto 0);
signal s1_2 : unsigned(17 downto 0);
signal s1_3 : unsigned(17 downto 0);
signal s2_1 : unsigned(17 downto 0);
signal s2_2 : unsigned(17 downto 0);
signal s2_3 : unsigned(17 downto 0);
signal s3_1 : unsigned(17 downto 0);
signal s3_2 : unsigned(17 downto 0);
signal s3_3 : unsigned(17 downto 0);
signal s4_1 : unsigned(17 downto 0);
signal s4_2 : unsigned(17 downto 0);
signal s4_3 : unsigned(17 downto 0);
signal s5_1 : unsigned(17 downto 0);
signal s5_2 : unsigned(17 downto 0);
signal s5_3 : unsigned(17 downto 0);
signal s6_1 : unsigned(17 downto 0);
signal s6_2 : unsigned(17 downto 0);
signal s6_3 : unsigned(17 downto 0);
signal s7_1 : unsigned(17 downto 0);
signal s7_2 : unsigned(17 downto 0);
signal s7_3 : unsigned(17 downto 0);
signal s8_1 : unsigned(17 downto 0);
signal s8_2 : unsigned(17 downto 0);
signal s8_3 : unsigned(17 downto 0);
component cf_cordic_r_18_18_18_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_26;
component cf_cordic_r_18_18_18_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_25;
component cf_cordic_r_18_18_18_23 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_23;
component cf_cordic_r_18_18_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_21;
component cf_cordic_r_18_18_18_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_19;
component cf_cordic_r_18_18_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_18;
component cf_cordic_r_18_18_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_17;
component cf_cordic_r_18_18_18_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_16;
begin
s1 : cf_cordic_r_18_18_18_26 port map (clock_c, i1, i2, s2_1, s2_2, s2_3, s1_1, s1_2, s1_3);
s2 : cf_cordic_r_18_18_18_25 port map (clock_c, i1, i2, s3_1, s3_2, s3_3, s2_1, s2_2, s2_3);
s3 : cf_cordic_r_18_18_18_23 port map (clock_c, i1, i2, s4_1, s4_2, s4_3, s3_1, s3_2, s3_3);
s4 : cf_cordic_r_18_18_18_21 port map (clock_c, i1, i2, s5_1, s5_2, s5_3, s4_1, s4_2, s4_3);
s5 : cf_cordic_r_18_18_18_19 port map (clock_c, i1, i2, s6_1, s6_2, s6_3, s5_1, s5_2, s5_3);
s6 : cf_cordic_r_18_18_18_18 port map (clock_c, i1, i2, s7_1, s7_2, s7_3, s6_1, s6_2, s6_3);
s7 : cf_cordic_r_18_18_18_17 port map (clock_c, i1, i2, s8_1, s8_2, s8_3, s7_1, s7_2, s7_3);
s8 : cf_cordic_r_18_18_18_16 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s1_3;
o2 <= s1_2;
o1 <= s1_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_14 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_14;
architecture rtl of cf_cordic_r_18_18_18_14 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(6 downto 0);
signal n8 : unsigned(7 downto 0);
signal n9 : unsigned(9 downto 0);
signal n10 : unsigned(17 downto 0);
begin
n1 <= i1(17 downto 17);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= n1 & n6;
n8 <= n1 & n7;
n9 <= i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8);
n10 <= n8 & n9;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_13;
architecture rtl of cf_cordic_r_18_18_18_13 is
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0) := "000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0) := "000000000000000000";
signal s15_1 : unsigned(17 downto 0);
signal s16_1 : unsigned(17 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_14 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_14;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "000000000010100011";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_r_18_18_18_14 port map (i3, s15_1);
s16 : cf_cordic_r_18_18_18_14 port map (i4, s16_1);
s17 : cf_cordic_r_18_18_18_31 port map (i5, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_12 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_12;
architecture rtl of cf_cordic_r_18_18_18_12 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(6 downto 0);
signal n8 : unsigned(10 downto 0);
signal n9 : unsigned(17 downto 0);
begin
n1 <= i1(17 downto 17);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= n1 & n6;
n8 <= i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7);
n9 <= n7 & n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_11;
architecture rtl of cf_cordic_r_18_18_18_11 is
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0) := "000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0) := "000000000000000000";
signal s15_1 : unsigned(17 downto 0);
signal s16_1 : unsigned(17 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_12 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_12;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "000000000101000110";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_r_18_18_18_12 port map (i3, s15_1);
s16 : cf_cordic_r_18_18_18_12 port map (i4, s16_1);
s17 : cf_cordic_r_18_18_18_31 port map (i5, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_10 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_10;
architecture rtl of cf_cordic_r_18_18_18_10 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(11 downto 0);
signal n8 : unsigned(17 downto 0);
begin
n1 <= i1(17 downto 17);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6);
n8 <= n6 & n7;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_9;
architecture rtl of cf_cordic_r_18_18_18_9 is
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0) := "000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0) := "000000000000000000";
signal s15_1 : unsigned(17 downto 0);
signal s16_1 : unsigned(17 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_10 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_10;
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "000000001010001100";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_r_18_18_18_10 port map (i3, s15_1);
s16 : cf_cordic_r_18_18_18_10 port map (i4, s16_1);
s17 : cf_cordic_r_18_18_18_31 port map (i5, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_8;
architecture rtl of cf_cordic_r_18_18_18_8 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(12 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0);
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0) := "000000000000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(1 downto 0);
signal n15 : unsigned(2 downto 0);
signal n16 : unsigned(3 downto 0);
signal n17 : unsigned(4 downto 0);
signal n18 : unsigned(12 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0);
signal n22 : unsigned(17 downto 0);
signal n23 : unsigned(17 downto 0) := "000000000000000000";
signal n24 : unsigned(17 downto 0);
signal n25 : unsigned(17 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0);
signal n28 : unsigned(17 downto 0) := "000000000000000000";
signal s29_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5);
n7 <= n5 & n6;
n8 <= i3 + n7;
n9 <= i3 - n7;
n10 <= n8 when s29_1 = "1" else n9;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n11 <= "000000000000000000";
    elsif i1 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= not s29_1;
n13 <= i3(17 downto 17);
n14 <= n13 & n13;
n15 <= n13 & n14;
n16 <= n13 & n15;
n17 <= n13 & n16;
n18 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5);
n19 <= n17 & n18;
n20 <= i4 + n19;
n21 <= i4 - n19;
n22 <= n20 when n12 = "1" else n21;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n23 <= "000000000000000000";
    elsif i1 = "1" then
      n23 <= n22;
    end if;
  end if;
end process;
n24 <= "000000010100010111";
n25 <= i5 + n24;
n26 <= i5 - n24;
n27 <= n25 when s29_1 = "1" else n26;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n28 <= "000000000000000000";
    elsif i1 = "1" then
      n28 <= n27;
    end if;
  end if;
end process;
s29 : cf_cordic_r_18_18_18_31 port map (i5, s29_1);
o3 <= n28;
o2 <= n23;
o1 <= n11;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_7;
architecture rtl of cf_cordic_r_18_18_18_7 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(13 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0);
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(1 downto 0);
signal n14 : unsigned(2 downto 0);
signal n15 : unsigned(3 downto 0);
signal n16 : unsigned(13 downto 0);
signal n17 : unsigned(17 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(17 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0);
signal n25 : unsigned(17 downto 0);
signal n26 : unsigned(17 downto 0) := "000000000000000000";
signal s27_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4);
n6 <= n4 & n5;
n7 <= i3 + n6;
n8 <= i3 - n6;
n9 <= n7 when s27_1 = "1" else n8;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n10 <= "000000000000000000";
    elsif i1 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
n11 <= not s27_1;
n12 <= i3(17 downto 17);
n13 <= n12 & n12;
n14 <= n12 & n13;
n15 <= n12 & n14;
n16 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4);
n17 <= n15 & n16;
n18 <= i4 + n17;
n19 <= i4 - n17;
n20 <= n18 when n11 = "1" else n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n21 <= "000000000000000000";
    elsif i1 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= "000000101000101100";
n23 <= i5 + n22;
n24 <= i5 - n22;
n25 <= n23 when s27_1 = "1" else n24;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n26 <= "000000000000000000";
    elsif i1 = "1" then
      n26 <= n25;
    end if;
  end if;
end process;
s27 : cf_cordic_r_18_18_18_31 port map (i5, s27_1);
o3 <= n26;
o2 <= n21;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_6;
architecture rtl of cf_cordic_r_18_18_18_6 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(14 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(1 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(14 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0);
signal n17 : unsigned(17 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0);
signal n22 : unsigned(17 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal s25_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3);
n5 <= n3 & n4;
n6 <= i3 + n5;
n7 <= i3 - n5;
n8 <= n6 when s25_1 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= not s25_1;
n11 <= i3(17 downto 17);
n12 <= n11 & n11;
n13 <= n11 & n12;
n14 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3);
n15 <= n13 & n14;
n16 <= i4 + n15;
n17 <= i4 - n15;
n18 <= n16 when n10 = "1" else n17;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n19 <= "000000000000000000";
    elsif i1 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= "000001010001000100";
n21 <= i5 + n20;
n22 <= i5 - n20;
n23 <= n21 when s25_1 = "1" else n22;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n24 <= "000000000000000000";
    elsif i1 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
s25 : cf_cordic_r_18_18_18_31 port map (i5, s25_1);
o3 <= n24;
o2 <= n19;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_5;
architecture rtl of cf_cordic_r_18_18_18_5 is
signal s1_1 : unsigned(17 downto 0);
signal s1_2 : unsigned(17 downto 0);
signal s1_3 : unsigned(17 downto 0);
signal s2_1 : unsigned(17 downto 0);
signal s2_2 : unsigned(17 downto 0);
signal s2_3 : unsigned(17 downto 0);
signal s3_1 : unsigned(17 downto 0);
signal s3_2 : unsigned(17 downto 0);
signal s3_3 : unsigned(17 downto 0);
signal s4_1 : unsigned(17 downto 0);
signal s4_2 : unsigned(17 downto 0);
signal s4_3 : unsigned(17 downto 0);
signal s5_1 : unsigned(17 downto 0);
signal s5_2 : unsigned(17 downto 0);
signal s5_3 : unsigned(17 downto 0);
signal s6_1 : unsigned(17 downto 0);
signal s6_2 : unsigned(17 downto 0);
signal s6_3 : unsigned(17 downto 0);
signal s7_1 : unsigned(17 downto 0);
signal s7_2 : unsigned(17 downto 0);
signal s7_3 : unsigned(17 downto 0);
signal s8_1 : unsigned(17 downto 0);
signal s8_2 : unsigned(17 downto 0);
signal s8_3 : unsigned(17 downto 0);
component cf_cordic_r_18_18_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_28;
component cf_cordic_r_18_18_18_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_15;
component cf_cordic_r_18_18_18_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_13;
component cf_cordic_r_18_18_18_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_11;
component cf_cordic_r_18_18_18_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_9;
component cf_cordic_r_18_18_18_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_8;
component cf_cordic_r_18_18_18_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_7;
component cf_cordic_r_18_18_18_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_6;
begin
s1 : cf_cordic_r_18_18_18_28 port map (clock_c, i1, i2, s3_1, s3_2, s3_3, s1_1, s1_2, s1_3);
s2 : cf_cordic_r_18_18_18_15 port map (clock_c, i1, i2, s1_1, s1_2, s1_3, s2_1, s2_2, s2_3);
s3 : cf_cordic_r_18_18_18_13 port map (clock_c, i1, i2, s4_1, s4_2, s4_3, s3_1, s3_2, s3_3);
s4 : cf_cordic_r_18_18_18_11 port map (clock_c, i1, i2, s5_1, s5_2, s5_3, s4_1, s4_2, s4_3);
s5 : cf_cordic_r_18_18_18_9 port map (clock_c, i1, i2, s6_1, s6_2, s6_3, s5_1, s5_2, s5_3);
s6 : cf_cordic_r_18_18_18_8 port map (clock_c, i1, i2, s7_1, s7_2, s7_3, s6_1, s6_2, s6_3);
s7 : cf_cordic_r_18_18_18_7 port map (clock_c, i1, i2, s8_1, s8_2, s8_3, s7_1, s7_2, s7_3);
s8 : cf_cordic_r_18_18_18_6 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_4;
architecture rtl of cf_cordic_r_18_18_18_4 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(16 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(16 downto 0);
signal n11 : unsigned(17 downto 0);
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0);
signal n15 : unsigned(17 downto 0) := "000000000000000000";
signal n16 : unsigned(17 downto 0);
signal n17 : unsigned(17 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0);
signal n20 : unsigned(17 downto 0) := "000000000000000000";
signal s21_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17);
n2 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3) &
  i4(2 downto 2) &
  i4(1 downto 1);
n3 <= n1 & n2;
n4 <= i3 + n3;
n5 <= i3 - n3;
n6 <= n4 when s21_1 = "1" else n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= not s21_1;
n9 <= i3(17 downto 17);
n10 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1);
n11 <= n9 & n10;
n12 <= i4 + n11;
n13 <= i4 - n11;
n14 <= n12 when n8 = "1" else n13;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n15 <= "000000000000000000";
    elsif i1 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
n16 <= "000100101110010000";
n17 <= i5 + n16;
n18 <= i5 - n16;
n19 <= n17 when s21_1 = "1" else n18;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n20 <= "000000000000000000";
    elsif i1 = "1" then
      n20 <= n19;
    end if;
  end if;
end process;
s21 : cf_cordic_r_18_18_18_31 port map (i5, s21_1);
o3 <= n20;
o2 <= n15;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_3;
architecture rtl of cf_cordic_r_18_18_18_3 is
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(17 downto 0) := "000000000000000000";
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0);
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0) := "000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(17 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_r_18_18_18_31 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_r_18_18_18_31;
begin
n1 <= i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3) &
  i4(2 downto 2) &
  i4(1 downto 1) &
  i4(0 downto 0);
n2 <= i3 + n1;
n3 <= i3 - n1;
n4 <= n2 when s17_1 = "1" else n3;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n5 <= "000000000000000000";
    elsif i1 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
n6 <= not s17_1;
n7 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= i4 + n7;
n9 <= i4 - n7;
n10 <= n8 when n6 = "1" else n9;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n11 <= "000000000000000000";
    elsif i1 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= "001000000000000000";
n13 <= i5 + n12;
n14 <= i5 - n12;
n15 <= n13 when s17_1 = "1" else n14;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n16 <= "000000000000000000";
    elsif i1 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
s17 : cf_cordic_r_18_18_18_31 port map (i5, s17_1);
o3 <= n16;
o2 <= n11;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
i6 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_2;
architecture rtl of cf_cordic_r_18_18_18_2 is
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(17 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0);
signal n11 : unsigned(17 downto 0) := "000000000000000000";
signal n12 : unsigned(17 downto 0);
begin
n1 <= "000000000000000000";
n2 <= n1 - i4;
n3 <= "000000000000000000";
n4 <= n3 - i5;
n5 <= i6 - n12;
n6 <= n2 when i3 = "1" else i4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= n4 when i3 = "1" else i5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= n5 when i3 = "1" else i6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n11 <= "000000000000000000";
    elsif i1 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= "100000000000000000";
o3 <= n11;
o2 <= n9;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
i6 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18_1;
architecture rtl of cf_cordic_r_18_18_18_1 is
signal n1 : unsigned(0 downto 0) := "0";
signal n2 : unsigned(17 downto 0) := "000000000000000000";
signal n3 : unsigned(17 downto 0) := "000000000000000000";
signal n4 : unsigned(17 downto 0) := "000000000000000000";
signal s5_1 : unsigned(17 downto 0);
signal s5_2 : unsigned(17 downto 0);
signal s5_3 : unsigned(17 downto 0);
signal s6_1 : unsigned(17 downto 0);
signal s6_2 : unsigned(17 downto 0);
signal s6_3 : unsigned(17 downto 0);
signal s7_1 : unsigned(17 downto 0);
signal s7_2 : unsigned(17 downto 0);
signal s7_3 : unsigned(17 downto 0);
signal s8_1 : unsigned(17 downto 0);
signal s8_2 : unsigned(17 downto 0);
signal s8_3 : unsigned(17 downto 0);
signal s9_1 : unsigned(17 downto 0);
signal s9_2 : unsigned(17 downto 0);
signal s9_3 : unsigned(17 downto 0);
component cf_cordic_r_18_18_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_30;
component cf_cordic_r_18_18_18_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_5;
component cf_cordic_r_18_18_18_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_4;
component cf_cordic_r_18_18_18_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_3;
component cf_cordic_r_18_18_18_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
i6 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_2;
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n1 <= "0";
    elsif i1 = "1" then
      n1 <= i3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n2 <= "000000000000000000";
    elsif i1 = "1" then
      n2 <= i4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n3 <= "000000000000000000";
    elsif i1 = "1" then
      n3 <= i5;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "000000000000000000";
    elsif i1 = "1" then
      n4 <= i6;
    end if;
  end if;
end process;
s5 : cf_cordic_r_18_18_18_30 port map (clock_c, i1, i2, s7_1, s7_2, s7_3, s5_1, s5_2, s5_3);
s6 : cf_cordic_r_18_18_18_5 port map (clock_c, i1, i2, s5_1, s5_2, s5_3, s6_1, s6_2, s6_3);
s7 : cf_cordic_r_18_18_18_4 port map (clock_c, i1, i2, s8_1, s8_2, s8_3, s7_1, s7_2, s7_3);
s8 : cf_cordic_r_18_18_18_3 port map (clock_c, i1, i2, s9_1, s9_2, s9_3, s8_1, s8_2, s8_3);
s9 : cf_cordic_r_18_18_18_2 port map (clock_c, i1, i2, n1, n2, n3, n4, s9_1, s9_2, s9_3);
o3 <= s6_3;
o2 <= s6_2;
o1 <= s6_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_r_18_18_18 is
port(
signal clock_c : in std_logic;
signal enable_i : in unsigned(0 downto 0);
signal reset_i : in unsigned(0 downto 0);
signal flip_i : in unsigned(0 downto 0);
signal real_i : in unsigned(17 downto 0);
signal imag_i : in unsigned(17 downto 0);
signal ang_i : in unsigned(17 downto 0);
signal real_o : out unsigned(17 downto 0);
signal imag_o : out unsigned(17 downto 0);
signal ang_o : out unsigned(17 downto 0));
end entity cf_cordic_r_18_18_18;
architecture rtl of cf_cordic_r_18_18_18 is
component cf_cordic_r_18_18_18_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(17 downto 0);
i5 : in  unsigned(17 downto 0);
i6 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0);
o3 : out unsigned(17 downto 0));
end component cf_cordic_r_18_18_18_1;
signal n1 : unsigned(17 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
begin
s1 : cf_cordic_r_18_18_18_1 port map (clock_c, enable_i, reset_i, flip_i, real_i, imag_i, ang_i, n1, n2, n3);
real_o <= n1;
imag_o <= n2;
ang_o <= n3;
end architecture rtl;


