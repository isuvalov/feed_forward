library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
library work;
use work.feedf_consts_pack.all;
use work.assert_pack.all;
use work.math_real.all;

USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

entity average_itertive_demod is
	generic(
		SIMULATION:integer:=1
	);
	port(
		clk : in STD_LOGIC;
		reset : in std_logic;
		after_pilot_start: in std_logic; --# �� ������ ���� ��� ������ i_ce
		i_ce : in std_logic;		
		i_samplesI: in std_logic_vector(15 downto 0);
		i_samplesQ: in std_logic_vector(15 downto 0);

		i_init_phaseI: in std_logic_vector(15 downto 0);
		i_init_phaseQ: in std_logic_vector(15 downto 0);

		o_samplesI: out std_logic_vector(15 downto 0);
		o_samplesQ: out std_logic_vector(15 downto 0);

		out_ce: out std_logic
		);
end average_itertive_demod;



architecture average_itertive_demod of average_itertive_demod is

function norming (val,x,y: std_logic_vector; rval:real) return std_logic_vector is
--# rval - future vector size
--# val - value that will be normalizate (or x or y)
--# x,y - input complex value
	variable abs_v:real;
	variable rett:std_logic_vector(val'Length-1 downto 0);
begin
	abs_v:=sqrt(real(conv_integer(signed(x)))*real(conv_integer(signed(x)))+real(conv_integer(signed(y)))*real(conv_integer(signed(y))) );
	if abs_v=0.0 then
		rett:=conv_std_logic_vector(0,val'Length);
	else
		rett:=conv_std_logic_vector(integer( rval*real(conv_integer(signed(val)))/abs_v ),val'Length);
	end if;
	return rett;
end norming;



function signed_abs (L: std_logic_vector) return std_logic_vector is
-- pragma label_applies_to abs
  
variable result : std_logic_vector(L'range) ;
--attribute IS_SIGNED of L:constant is TRUE ;
--attribute SYNTHESIS_RETURN of result:variable is "ABS" ;
begin
if (L(L'left) = '0' or L(L'left) = 'L') then
    result := L;
else
    result := 0 - signed(L);
end if;
    return result ;
end signed_abs;



function int_abs (L: integer) return integer is
	variable result : integer;
begin
	if (L>0) then
    	result := L;
	else
    	result := 0 - L;
	end if;
    return result ;
end int_abs;


constant NORMBIT:natural:=6;
constant NORMBITOUT:natural:=12;


type Tnorm_mem is array (0 to 4095) of std_logic_vector(11 downto 0);
constant norm_mem:Tnorm_mem:=  (
"111111111111", "100000000000", "010000000000", "001010101011", "001000000000", "000110011010", "000101010101", "000100100101", "000100000000", "000011100100", 
"000011001101", "000010111010", "000010101011", "000010011110", "000010010010", "000010001001", "000010000000", "000001111000", "000001110010", "000001101100", 
"000001100110", "000001100010", "000001011101", "000001011001", "000001010101", "000001010010", "000001001111", "000001001100", "000001001001", "000001000111", 
"000001000100", "000001000010", "000001000000", "000001000010", "000001000100", "000001000111", "000001001001", "000001001100", "000001001111", "000001010010", 
"000001010101", "000001011001", "000001011101", "000001100010", "000001100110", "000001101100", "000001110010", "000001111000", "000010000000", "000010001001", 
"000010010010", "000010011110", "000010101011", "000010111010", "000011001101", "000011100100", "000100000000", "000100100101", "000101010101", "000110011010", 
"001000000000", "001010101011", "010000000000", "100000000000", "100000000000", "010110101000", "001110010100", "001010000111", "000111110001", "000110010010", 
"000101010001", "000100100010", "000011111110", "000011100010", "000011001100", "000010111001", "000010101010", "000010011101", "000010010010", "000010001000", 
"000010000000", "000001111000", "000001110010", "000001101100", "000001100110", "000001100001", "000001011101", "000001011001", "000001010101", "000001010010", 
"000001001111", "000001001100", "000001001001", "000001000111", "000001000100", "000001000010", "000001000000", "000001000010", "000001000100", "000001000111", 
"000001001001", "000001001100", "000001001111", "000001010010", "000001010101", "000001011001", "000001011101", "000001100001", "000001100110", "000001101100", 
"000001110010", "000001111000", "000010000000", "000010001000", "000010010010", "000010011101", "000010101010", "000010111001", "000011001100", "000011100010", 
"000011111110", "000100100010", "000101010001", "000110010010", "000111110001", "001010000111", "001110010100", "010110101000", "010000000000", "001110010100", 
"001011010100", "001000111000", "000111001010", "000101111100", "000101000100", "000100011001", "000011111000", "000011011110", "000011001001", "000010110111", 
"000010101000", "000010011100", "000010010001", "000010000111", "000001111111", "000001111000", "000001110001", "000001101011", "000001100110", "000001100001", 
"000001011101", "000001011001", "000001010101", "000001010010", "000001001111", "000001001100", "000001001001", "000001000110", "000001000100", "000001000010", 
"000001000000", "000001000010", "000001000100", "000001000110", "000001001001", "000001001100", "000001001111", "000001010010", "000001010101", "000001011001", 
"000001011101", "000001100001", "000001100110", "000001101011", "000001110001", "000001111000", "000001111111", "000010000111", "000010010001", "000010011100", 
"000010101000", "000010110111", "000011001001", "000011011110", "000011111000", "000100011001", "000101000100", "000101111100", "000111001010", "001000111000", 
"001011010100", "001110010100", "001010101011", "001010000111", "001000111000", "000111100011", "000110011010", "000101011111", "000100110001", "000100001101", 
"000011110000", "000011011000", "000011000100", "000010110100", "000010100110", "000010011001", "000010001111", "000010000110", "000001111110", "000001110111", 
"000001110000", "000001101010", "000001100101", "000001100001", "000001011100", "000001011000", "000001010101", "000001010001", "000001001110", "000001001011", 
"000001001001", "000001000110", "000001000100", "000001000010", "000001000000", "000001000010", "000001000100", "000001000110", "000001001001", "000001001011", 
"000001001110", "000001010001", "000001010101", "000001011000", "000001011100", "000001100001", "000001100101", "000001101010", "000001110000", "000001110111", 
"000001111110", "000010000110", "000010001111", "000010011001", "000010100110", "000010110100", "000011000100", "000011011000", "000011110000", "000100001101", 
"000100110001", "000101011111", "000110011010", "000111100011", "001000111000", "001010000111", "001000000000", "000111110001", "000111001010", "000110011010", 
"000101101010", "000101000000", "000100011100", "000011111110", "000011100101", "000011010000", "000010111110", "000010101111", "000010100010", "000010010111", 
"000010001101", "000010000100", "000001111100", "000001110101", "000001101111", "000001101001", "000001100100", "000001100000", "000001011100", "000001011000", 
"000001010100", "000001010001", "000001001110", "000001001011", "000001001000", "000001000110", "000001000100", "000001000010", "000000111111", "000001000010", 
"000001000100", "000001000110", "000001001000", "000001001011", "000001001110", "000001010001", "000001010100", "000001011000", "000001011100", "000001100000", 
"000001100100", "000001101001", "000001101111", "000001110101", "000001111100", "000010000100", "000010001101", "000010010111", "000010100010", "000010101111", 
"000010111110", "000011010000", "000011100101", "000011111110", "000100011100", "000101000000", "000101101010", "000110011010", "000111001010", "000111110001", 
"000110011010", "000110010010", "000101111100", "000101011111", "000101000000", "000100100010", "000100000110", "000011101110", "000011011001", "000011000111", 
"000010110111", "000010101001", "000010011110", "000010010011", "000010001010", "000010000001", "000001111010", "000001110100", "000001101110", "000001101000", 
"000001100011", "000001011111", "000001011011", "000001010111", "000001010100", "000001010000", "000001001101", "000001001011", "000001001000", "000001000110", 
"000001000011", "000001000001", "000000111111", "000001000001", "000001000011", "000001000110", "000001001000", "000001001011", "000001001101", "000001010000", 
"000001010100", "000001010111", "000001011011", "000001011111", "000001100011", "000001101000", "000001101110", "000001110100", "000001111010", "000010000001", 
"000010001010", "000010010011", "000010011110", "000010101001", "000010110111", "000011000111", "000011011001", "000011101110", "000100000110", "000100100010", 
"000101000000", "000101011111", "000101111100", "000110010010", "000101010101", "000101010001", "000101000100", "000100110001", "000100011100", "000100000110", 
"000011110001", "000011011110", "000011001101", "000010111101", "000010110000", "000010100011", "000010011001", "000010001111", "000010000110", "000001111111", 
"000001111000", "000001110010", "000001101100", "000001100111", "000001100010", "000001011110", "000001011010", "000001010110", "000001010011", "000001010000", 
"000001001101", "000001001010", "000001001000", "000001000101", "000001000011", "000001000001", "000000111111", "000001000001", "000001000011", "000001000101", 
"000001001000", "000001001010", "000001001101", "000001010000", "000001010011", "000001010110", "000001011010", "000001011110", "000001100010", "000001100111", 
"000001101100", "000001110010", "000001111000", "000001111111", "000010000110", "000010001111", "000010011001", "000010100011", "000010110000", "000010111101", 
"000011001101", "000011011110", "000011110001", "000100000110", "000100011100", "000100110001", "000101000100", "000101010001", "000100100101", "000100100010", 
"000100011001", "000100001101", "000011111110", "000011101110", "000011011110", "000011001111", "000011000001", "000010110100", "000010101000", "000010011101", 
"000010010011", "000010001011", "000010000011", "000001111100", "000001110101", "000001101111", "000001101010", "000001100101", "000001100001", "000001011100", 
"000001011001", "000001010101", "000001010010", "000001001111", "000001001100", "000001001001", "000001000111", "000001000101", "000001000010", "000001000000", 
"000000111111", "000001000000", "000001000010", "000001000101", "000001000111", "000001001001", "000001001100", "000001001111", "000001010010", "000001010101", 
"000001011001", "000001011100", "000001100001", "000001100101", "000001101010", "000001101111", "000001110101", "000001111100", "000010000011", "000010001011", 
"000010010011", "000010011101", "000010101000", "000010110100", "000011000001", "000011001111", "000011011110", "000011101110", "000011111110", "000100001101", 
"000100011001", "000100100010", "000100000000", "000011111110", "000011111000", "000011110000", "000011100101", "000011011001", "000011001101", "000011000001", 
"000010110101", "000010101010", "000010100000", "000010010111", "000010001110", "000010000110", "000001111111", "000001111000", "000001110010", "000001101101", 
"000001101000", "000001100011", "000001011111", "000001011011", "000001010111", "000001010100", "000001010001", "000001001110", "000001001011", "000001001001", 
"000001000110", "000001000100", "000001000010", "000001000000", "000000111110", "000001000000", "000001000010", "000001000100", "000001000110", "000001001001", 
"000001001011", "000001001110", "000001010001", "000001010100", "000001010111", "000001011011", "000001011111", "000001100011", "000001101000", "000001101101", 
"000001110010", "000001111000", "000001111111", "000010000110", "000010001110", "000010010111", "000010100000", "000010101010", "000010110101", "000011000001", 
"000011001101", "000011011001", "000011100101", "000011110000", "000011111000", "000011111110", "000011100100", "000011100010", "000011011110", "000011011000", 
"000011010000", "000011000111", "000010111101", "000010110100", "000010101010", "000010100001", "000010011000", "000010010000", "000010001001", "000010000001", 
"000001111011", "000001110101", "000001110000", "000001101010", "000001100110", "000001100001", "000001011101", "000001011010", "000001010110", "000001010011", 
"000001010000", "000001001101", "000001001010", "000001001000", "000001000110", "000001000011", "000001000001", "000000111111", "000000111110", "000000111111", 
"000001000001", "000001000011", "000001000110", "000001001000", "000001001010", "000001001101", "000001010000", "000001010011", "000001010110", "000001011010", 
"000001011101", "000001100001", "000001100110", "000001101010", "000001110000", "000001110101", "000001111011", "000010000001", "000010001001", "000010010000", 
"000010011000", "000010100001", "000010101010", "000010110100", "000010111101", "000011000111", "000011010000", "000011011000", "000011011110", "000011100010", 
"000011001101", "000011001100", "000011001001", "000011000100", "000010111110", "000010110111", "000010110000", "000010101000", "000010100000", "000010011000", 
"000010010001", "000010001010", "000010000011", "000001111101", "000001110111", "000001110010", "000001101101", "000001101000", "000001100011", "000001011111", 
"000001011100", "000001011000", "000001010101", "000001010010", "000001001111", "000001001100", "000001001010", "000001000111", "000001000101", "000001000011", 
"000001000001", "000000111111", "000000111101", "000000111111", "000001000001", "000001000011", "000001000101", "000001000111", "000001001010", "000001001100", 
"000001001111", "000001010010", "000001010101", "000001011000", "000001011100", "000001011111", "000001100011", "000001101000", "000001101101", "000001110010", 
"000001110111", "000001111101", "000010000011", "000010001010", "000010010001", "000010011000", "000010100000", "000010101000", "000010110000", "000010110111", 
"000010111110", "000011000100", "000011001001", "000011001100", "000010111010", "000010111001", "000010110111", "000010110100", "000010101111", "000010101001", 
"000010100011", "000010011101", "000010010111", "000010010000", "000010001010", "000010000100", "000001111110", "000001111000", "000001110011", "000001101110", 
"000001101001", "000001100101", "000001100001", "000001011101", "000001011010", "000001010110", "000001010011", "000001010000", "000001001110", "000001001011", 
"000001001001", "000001000110", "000001000100", "000001000010", "000001000000", "000000111110", "000000111101", "000000111110", "000001000000", "000001000010", 
"000001000100", "000001000110", "000001001001", "000001001011", "000001001110", "000001010000", "000001010011", "000001010110", "000001011010", "000001011101", 
"000001100001", "000001100101", "000001101001", "000001101110", "000001110011", "000001111000", "000001111110", "000010000100", "000010001010", "000010010000", 
"000010010111", "000010011101", "000010100011", "000010101001", "000010101111", "000010110100", "000010110111", "000010111001", "000010101011", "000010101010", 
"000010101000", "000010100110", "000010100010", "000010011110", "000010011001", "000010010011", "000010001110", "000010001001", "000010000011", "000001111110", 
"000001111001", "000001110100", "000001101111", "000001101011", "000001100110", "000001100010", "000001011111", "000001011011", "000001011000", "000001010101", 
"000001010010", "000001001111", "000001001100", "000001001010", "000001001000", "000001000101", "000001000011", "000001000001", "000000111111", "000000111110", 
"000000111100", "000000111110", "000000111111", "000001000001", "000001000011", "000001000101", "000001001000", "000001001010", "000001001100", "000001001111", 
"000001010010", "000001010101", "000001011000", "000001011011", "000001011111", "000001100010", "000001100110", "000001101011", "000001101111", "000001110100", 
"000001111001", "000001111110", "000010000011", "000010001001", "000010001110", "000010010011", "000010011001", "000010011110", "000010100010", "000010100110", 
"000010101000", "000010101010", "000010011110", "000010011101", "000010011100", "000010011001", "000010010111", "000010010011", "000010001111", "000010001011", 
"000010000110", "000010000001", "000001111101", "000001111000", "000001110100", "000001101111", "000001101011", "000001100111", "000001100011", "000001100000", 
"000001011100", "000001011001", "000001010110", "000001010011", "000001010000", "000001001101", "000001001011", "000001001001", "000001000110", "000001000100", 
"000001000010", "000001000000", "000000111111", "000000111101", "000000111011", "000000111101", "000000111111", "000001000000", "000001000010", "000001000100", 
"000001000110", "000001001001", "000001001011", "000001001101", "000001010000", "000001010011", "000001010110", "000001011001", "000001011100", "000001100000", 
"000001100011", "000001100111", "000001101011", "000001101111", "000001110100", "000001111000", "000001111101", "000010000001", "000010000110", "000010001011", 
"000010001111", "000010010011", "000010010111", "000010011001", "000010011100", "000010011101", "000010010010", "000010010010", "000010010001", "000010001111", 
"000010001101", "000010001010", "000010000110", "000010000011", "000001111111", "000001111011", "000001110111", "000001110011", "000001101111", "000001101011", 
"000001100111", "000001100100", "000001100000", "000001011101", "000001011010", "000001010111", "000001010100", "000001010001", "000001001111", "000001001100", 
"000001001010", "000001000111", "000001000101", "000001000011", "000001000001", "000001000000", "000000111110", "000000111100", "000000111011", "000000111100", 
"000000111110", "000001000000", "000001000001", "000001000011", "000001000101", "000001000111", "000001001010", "000001001100", "000001001111", "000001010001", 
"000001010100", "000001010111", "000001011010", "000001011101", "000001100000", "000001100100", "000001100111", "000001101011", "000001101111", "000001110011", 
"000001110111", "000001111011", "000001111111", "000010000011", "000010000110", "000010001010", "000010001101", "000010001111", "000010010001", "000010010010", 
"000010001001", "000010001000", "000010000111", "000010000110", "000010000100", "000010000001", "000001111111", "000001111100", "000001111000", "000001110101", 
"000001110010", "000001101110", "000001101011", "000001100111", "000001100100", "000001100001", "000001011101", "000001011010", "000001010111", "000001010101", 
"000001010010", "000001001111", "000001001101", "000001001011", "000001001000", "000001000110", "000001000100", "000001000010", "000001000000", "000000111111", 
"000000111101", "000000111011", "000000111010", "000000111011", "000000111101", "000000111111", "000001000000", "000001000010", "000001000100", "000001000110", 
"000001001000", "000001001011", "000001001101", "000001001111", "000001010010", "000001010101", "000001010111", "000001011010", "000001011101", "000001100001", 
"000001100100", "000001100111", "000001101011", "000001101110", "000001110010", "000001110101", "000001111000", "000001111100", "000001111111", "000010000001", 
"000010000100", "000010000110", "000010000111", "000010001000", "000010000000", "000010000000", "000001111111", "000001111110", "000001111100", "000001111010", 
"000001111000", "000001110101", "000001110010", "000001110000", "000001101101", "000001101001", "000001100110", "000001100011", "000001100000", "000001011101", 
"000001011010", "000001011000", "000001010101", "000001010010", "000001010000", "000001001110", "000001001011", "000001001001", "000001000111", "000001000101", 
"000001000011", "000001000001", "000000111111", "000000111110", "000000111100", "000000111011", "000000111001", "000000111011", "000000111100", "000000111110", 
"000000111111", "000001000001", "000001000011", "000001000101", "000001000111", "000001001001", "000001001011", "000001001110", "000001010000", "000001010010", 
"000001010101", "000001011000", "000001011010", "000001011101", "000001100000", "000001100011", "000001100110", "000001101001", "000001101101", "000001110000", 
"000001110010", "000001110101", "000001111000", "000001111010", "000001111100", "000001111110", "000001111111", "000010000000", "000001111000", "000001111000", 
"000001111000", "000001110111", "000001110101", "000001110100", "000001110010", "000001101111", "000001101101", "000001101010", "000001101000", "000001100101", 
"000001100010", "000001100000", "000001011101", "000001011010", "000001011000", "000001010101", "000001010011", "000001010000", "000001001110", "000001001100", 
"000001001010", "000001001000", "000001000110", "000001000100", "000001000010", "000001000000", "000000111111", "000000111101", "000000111011", "000000111010", 
"000000111001", "000000111010", "000000111011", "000000111101", "000000111111", "000001000000", "000001000010", "000001000100", "000001000110", "000001001000", 
"000001001010", "000001001100", "000001001110", "000001010000", "000001010011", "000001010101", "000001011000", "000001011010", "000001011101", "000001100000", 
"000001100010", "000001100101", "000001101000", "000001101010", "000001101101", "000001101111", "000001110010", "000001110100", "000001110101", "000001110111", 
"000001111000", "000001111000", "000001110010", "000001110010", "000001110001", "000001110000", "000001101111", "000001101110", "000001101100", "000001101010", 
"000001101000", "000001100110", "000001100011", "000001100001", "000001011111", "000001011100", "000001011010", "000001010111", "000001010101", "000001010011", 
"000001010000", "000001001110", "000001001100", "000001001010", "000001001000", "000001000110", "000001000100", "000001000010", "000001000001", "000000111111", 
"000000111110", "000000111100", "000000111011", "000000111001", "000000111000", "000000111001", "000000111011", "000000111100", "000000111110", "000000111111", 
"000001000001", "000001000010", "000001000100", "000001000110", "000001001000", "000001001010", "000001001100", "000001001110", "000001010000", "000001010011", 
"000001010101", "000001010111", "000001011010", "000001011100", "000001011111", "000001100001", "000001100011", "000001100110", "000001101000", "000001101010", 
"000001101100", "000001101110", "000001101111", "000001110000", "000001110001", "000001110010", "000001101100", "000001101100", "000001101011", "000001101010", 
"000001101001", "000001101000", "000001100111", "000001100101", "000001100011", "000001100001", "000001011111", "000001011101", "000001011011", "000001011001", 
"000001010111", "000001010101", "000001010010", "000001010000", "000001001110", "000001001100", "000001001010", "000001001000", "000001000110", "000001000101", 
"000001000011", "000001000001", "000001000000", "000000111110", "000000111101", "000000111011", "000000111010", "000000111000", "000000110111", "000000111000", 
"000000111010", "000000111011", "000000111101", "000000111110", "000001000000", "000001000001", "000001000011", "000001000101", "000001000110", "000001001000", 
"000001001010", "000001001100", "000001001110", "000001010000", "000001010010", "000001010101", "000001010111", "000001011001", "000001011011", "000001011101", 
"000001011111", "000001100001", "000001100011", "000001100101", "000001100111", "000001101000", "000001101001", "000001101010", "000001101011", "000001101100", 
"000001100110", "000001100110", "000001100110", "000001100101", "000001100100", "000001100011", "000001100010", "000001100001", "000001011111", "000001011101", 
"000001011100", "000001011010", "000001011000", "000001010110", "000001010100", "000001010010", "000001010000", "000001001110", "000001001100", "000001001010", 
"000001001000", "000001000111", "000001000101", "000001000011", "000001000010", "000001000000", "000000111110", "000000111101", "000000111100", "000000111010", 
"000000111001", "000000111000", "000000110110", "000000111000", "000000111001", "000000111010", "000000111100", "000000111101", "000000111110", "000001000000", 
"000001000010", "000001000011", "000001000101", "000001000111", "000001001000", "000001001010", "000001001100", "000001001110", "000001010000", "000001010010", 
"000001010100", "000001010110", "000001011000", "000001011010", "000001011100", "000001011101", "000001011111", "000001100001", "000001100010", "000001100011", 
"000001100100", "000001100101", "000001100110", "000001100110", "000001100010", "000001100001", "000001100001", "000001100001", "000001100000", "000001011111", 
"000001011110", "000001011100", "000001011011", "000001011010", "000001011000", "000001010110", "000001010101", "000001010011", "000001010001", "000001001111", 
"000001001110", "000001001100", "000001001010", "000001001000", "000001000111", "000001000101", "000001000011", "000001000010", "000001000000", "000000111111", 
"000000111101", "000000111100", "000000111011", "000000111001", "000000111000", "000000110111", "000000110101", "000000110111", "000000111000", "000000111001", 
"000000111011", "000000111100", "000000111101", "000000111111", "000001000000", "000001000010", "000001000011", "000001000101", "000001000111", "000001001000", 
"000001001010", "000001001100", "000001001110", "000001001111", "000001010001", "000001010011", "000001010101", "000001010110", "000001011000", "000001011010", 
"000001011011", "000001011100", "000001011110", "000001011111", "000001100000", "000001100001", "000001100001", "000001100001", "000001011101", "000001011101", 
"000001011101", "000001011100", "000001011100", "000001011011", "000001011010", "000001011001", "000001010111", "000001010110", "000001010101", "000001010011", 
"000001010010", "000001010000", "000001001111", "000001001101", "000001001011", "000001001010", "000001001000", "000001000110", "000001000101", "000001000011", 
"000001000010", "000001000000", "000000111111", "000000111101", "000000111100", "000000111011", "000000111001", "000000111000", "000000110111", "000000110110", 
"000000110101", "000000110110", "000000110111", "000000111000", "000000111001", "000000111011", "000000111100", "000000111101", "000000111111", "000001000000", 
"000001000010", "000001000011", "000001000101", "000001000110", "000001001000", "000001001010", "000001001011", "000001001101", "000001001111", "000001010000", 
"000001010010", "000001010011", "000001010101", "000001010110", "000001010111", "000001011001", "000001011010", "000001011011", "000001011100", "000001011100", 
"000001011101", "000001011101", "000001011001", "000001011001", "000001011001", "000001011000", "000001011000", "000001010111", "000001010110", "000001010101", 
"000001010100", "000001010011", "000001010010", "000001010000", "000001001111", "000001001101", "000001001100", "000001001011", "000001001001", "000001001000", 
"000001000110", "000001000101", "000001000011", "000001000010", "000001000000", "000000111111", "000000111110", "000000111100", "000000111011", "000000111010", 
"000000111001", "000000110111", "000000110110", "000000110101", "000000110100", "000000110101", "000000110110", "000000110111", "000000111001", "000000111010", 
"000000111011", "000000111100", "000000111110", "000000111111", "000001000000", "000001000010", "000001000011", "000001000101", "000001000110", "000001001000", 
"000001001001", "000001001011", "000001001100", "000001001101", "000001001111", "000001010000", "000001010010", "000001010011", "000001010100", "000001010101", 
"000001010110", "000001010111", "000001011000", "000001011000", "000001011001", "000001011001", "000001010101", "000001010101", "000001010101", "000001010101", 
"000001010100", "000001010100", "000001010011", "000001010010", "000001010001", "000001010000", "000001001111", "000001001110", "000001001100", "000001001011", 
"000001001010", "000001001000", "000001000111", "000001000110", "000001000100", "000001000011", "000001000010", "000001000000", "000000111111", "000000111110", 
"000000111100", "000000111011", "000000111010", "000000111001", "000000111000", "000000110110", "000000110101", "000000110100", "000000110011", "000000110100", 
"000000110101", "000000110110", "000000111000", "000000111001", "000000111010", "000000111011", "000000111100", "000000111110", "000000111111", "000001000000", 
"000001000010", "000001000011", "000001000100", "000001000110", "000001000111", "000001001000", "000001001010", "000001001011", "000001001100", "000001001110", 
"000001001111", "000001010000", "000001010001", "000001010010", "000001010011", "000001010100", "000001010100", "000001010101", "000001010101", "000001010101", 
"000001010010", "000001010010", "000001010010", "000001010001", "000001010001", "000001010000", "000001010000", "000001001111", "000001001110", "000001001101", 
"000001001100", "000001001011", "000001001010", "000001001001", "000001000111", "000001000110", "000001000101", "000001000100", "000001000010", "000001000001", 
"000001000000", "000000111111", "000000111101", "000000111100", "000000111011", "000000111010", "000000111001", "000000111000", "000000110111", "000000110101", 
"000000110100", "000000110011", "000000110010", "000000110011", "000000110100", "000000110101", "000000110111", "000000111000", "000000111001", "000000111010", 
"000000111011", "000000111100", "000000111101", "000000111111", "000001000000", "000001000001", "000001000010", "000001000100", "000001000101", "000001000110", 
"000001000111", "000001001001", "000001001010", "000001001011", "000001001100", "000001001101", "000001001110", "000001001111", "000001010000", "000001010000", 
"000001010001", "000001010001", "000001010010", "000001010010", "000001001111", "000001001111", "000001001111", "000001001110", "000001001110", "000001001101", 
"000001001101", "000001001100", "000001001011", "000001001010", "000001001010", "000001001001", "000001001000", "000001000110", "000001000101", "000001000100", 
"000001000011", "000001000010", "000001000001", "000001000000", "000000111110", "000000111101", "000000111100", "000000111011", "000000111010", "000000111001", 
"000000111000", "000000110111", "000000110110", "000000110101", "000000110100", "000000110011", "000000110010", "000000110011", "000000110100", "000000110101", 
"000000110110", "000000110111", "000000111000", "000000111001", "000000111010", "000000111011", "000000111100", "000000111101", "000000111110", "000001000000", 
"000001000001", "000001000010", "000001000011", "000001000100", "000001000101", "000001000110", "000001001000", "000001001001", "000001001010", "000001001010", 
"000001001011", "000001001100", "000001001101", "000001001101", "000001001110", "000001001110", "000001001111", "000001001111", "000001001100", "000001001100", 
"000001001100", "000001001011", "000001001011", "000001001011", "000001001010", "000001001001", "000001001001", "000001001000", "000001000111", "000001000110", 
"000001000101", "000001000100", "000001000011", "000001000010", "000001000001", "000001000000", "000000111111", "000000111110", "000000111101", "000000111100", 
"000000111011", "000000111010", "000000111001", "000000111000", "000000110111", "000000110110", "000000110101", "000000110100", "000000110011", "000000110010", 
"000000110001", "000000110010", "000000110011", "000000110100", "000000110101", "000000110110", "000000110111", "000000111000", "000000111001", "000000111010", 
"000000111011", "000000111100", "000000111101", "000000111110", "000000111111", "000001000000", "000001000001", "000001000010", "000001000011", "000001000100", 
"000001000101", "000001000110", "000001000111", "000001001000", "000001001001", "000001001001", "000001001010", "000001001011", "000001001011", "000001001011", 
"000001001100", "000001001100", "000001001001", "000001001001", "000001001001", "000001001001", "000001001000", "000001001000", "000001001000", "000001000111", 
"000001000110", "000001000110", "000001000101", "000001000100", "000001000011", "000001000010", "000001000001", "000001000000", "000000111111", "000000111111", 
"000000111110", "000000111101", "000000111100", "000000111011", "000000111001", "000000111001", "000000111000", "000000110111", "000000110110", "000000110101", 
"000000110100", "000000110011", "000000110010", "000000110001", "000000110000", "000000110001", "000000110010", "000000110011", "000000110100", "000000110101", 
"000000110110", "000000110111", "000000111000", "000000111001", "000000111001", "000000111011", "000000111100", "000000111101", "000000111110", "000000111111", 
"000000111111", "000001000000", "000001000001", "000001000010", "000001000011", "000001000100", "000001000101", "000001000110", "000001000110", "000001000111", 
"000001001000", "000001001000", "000001001000", "000001001001", "000001001001", "000001001001", "000001000111", "000001000111", "000001000110", "000001000110", 
"000001000110", "000001000110", "000001000101", "000001000101", "000001000100", "000001000011", "000001000011", "000001000010", "000001000001", "000001000000", 
"000001000000", "000000111111", "000000111110", "000000111101", "000000111100", "000000111011", "000000111010", "000000111001", "000000111000", "000000110111", 
"000000110110", "000000110101", "000000110101", "000000110100", "000000110011", "000000110010", "000000110001", "000000110000", "000000101111", "000000110000", 
"000000110001", "000000110010", "000000110011", "000000110100", "000000110101", "000000110101", "000000110110", "000000110111", "000000111000", "000000111001", 
"000000111010", "000000111011", "000000111100", "000000111101", "000000111110", "000000111111", "000001000000", "000001000000", "000001000001", "000001000010", 
"000001000011", "000001000011", "000001000100", "000001000101", "000001000101", "000001000110", "000001000110", "000001000110", "000001000110", "000001000111", 
"000001000100", "000001000100", "000001000100", "000001000100", "000001000100", "000001000011", "000001000011", "000001000010", "000001000010", "000001000001", 
"000001000001", "000001000000", "000000111111", "000000111111", "000000111110", "000000111101", "000000111100", "000000111011", "000000111011", "000000111010", 
"000000111001", "000000111000", "000000110111", "000000110110", "000000110101", "000000110100", "000000110100", "000000110011", "000000110010", "000000110001", 
"000000110000", "000000101111", "000000101111", "000000101111", "000000110000", "000000110001", "000000110010", "000000110011", "000000110100", "000000110100", 
"000000110101", "000000110110", "000000110111", "000000111000", "000000111001", "000000111010", "000000111011", "000000111011", "000000111100", "000000111101", 
"000000111110", "000000111111", "000000111111", "000001000000", "000001000001", "000001000001", "000001000010", "000001000010", "000001000011", "000001000011", 
"000001000100", "000001000100", "000001000100", "000001000100", "000001000010", "000001000010", "000001000010", "000001000010", "000001000010", "000001000001", 
"000001000001", "000001000000", "000001000000", "000000111111", "000000111111", "000000111110", "000000111110", "000000111101", "000000111100", "000000111011", 
"000000111011", "000000111010", "000000111001", "000000111000", "000000111000", "000000110111", "000000110110", "000000110101", "000000110100", "000000110011", 
"000000110011", "000000110010", "000000110001", "000000110000", "000000101111", "000000101111", "000000101110", "000000101111", "000000101111", "000000110000", 
"000000110001", "000000110010", "000000110011", "000000110011", "000000110100", "000000110101", "000000110110", "000000110111", "000000111000", "000000111000", 
"000000111001", "000000111010", "000000111011", "000000111011", "000000111100", "000000111101", "000000111110", "000000111110", "000000111111", "000000111111", 
"000001000000", "000001000000", "000001000001", "000001000001", "000001000010", "000001000010", "000001000010", "000001000010", "000001000000", "000001000000", 
"000001000000", "000001000000", "000000111111", "000000111111", "000000111111", "000000111111", "000000111110", "000000111110", "000000111101", "000000111101", 
"000000111100", "000000111011", "000000111011", "000000111010", "000000111001", "000000111001", "000000111000", "000000110111", "000000110110", "000000110101", 
"000000110101", "000000110100", "000000110011", "000000110010", "000000110010", "000000110001", "000000110000", "000000101111", "000000101111", "000000101110", 
"000000101101", "000000101110", "000000101111", "000000101111", "000000110000", "000000110001", "000000110010", "000000110010", "000000110011", "000000110100", 
"000000110101", "000000110101", "000000110110", "000000110111", "000000111000", "000000111001", "000000111001", "000000111010", "000000111011", "000000111011", 
"000000111100", "000000111101", "000000111101", "000000111110", "000000111110", "000000111111", "000000111111", "000000111111", "000000111111", "000001000000", 
"000001000000", "000001000000", "000001000010", "000001000010", "000001000010", "000001000010", "000001000010", "000001000001", "000001000001", "000001000000", 
"000001000000", "000000111111", "000000111111", "000000111110", "000000111110", "000000111101", "000000111100", "000000111011", "000000111011", "000000111010", 
"000000111001", "000000111000", "000000111000", "000000110111", "000000110110", "000000110101", "000000110100", "000000110011", "000000110011", "000000110010", 
"000000110001", "000000110000", "000000101111", "000000101111", "000000101110", "000000101111", "000000101111", "000000110000", "000000110001", "000000110010", 
"000000110011", "000000110011", "000000110100", "000000110101", "000000110110", "000000110111", "000000111000", "000000111000", "000000111001", "000000111010", 
"000000111011", "000000111011", "000000111100", "000000111101", "000000111110", "000000111110", "000000111111", "000000111111", "000001000000", "000001000000", 
"000001000001", "000001000001", "000001000010", "000001000010", "000001000010", "000001000010", "000001000100", "000001000100", "000001000100", "000001000100", 
"000001000100", "000001000011", "000001000011", "000001000010", "000001000010", "000001000001", "000001000001", "000001000000", "000000111111", "000000111111", 
"000000111110", "000000111101", "000000111100", "000000111011", "000000111011", "000000111010", "000000111001", "000000111000", "000000110111", "000000110110", 
"000000110101", "000000110100", "000000110100", "000000110011", "000000110010", "000000110001", "000000110000", "000000101111", "000000101111", "000000101111", 
"000000110000", "000000110001", "000000110010", "000000110011", "000000110100", "000000110100", "000000110101", "000000110110", "000000110111", "000000111000", 
"000000111001", "000000111010", "000000111011", "000000111011", "000000111100", "000000111101", "000000111110", "000000111111", "000000111111", "000001000000", 
"000001000001", "000001000001", "000001000010", "000001000010", "000001000011", "000001000011", "000001000100", "000001000100", "000001000100", "000001000100", 
"000001000111", "000001000111", "000001000110", "000001000110", "000001000110", "000001000110", "000001000101", "000001000101", "000001000100", "000001000011", 
"000001000011", "000001000010", "000001000001", "000001000000", "000001000000", "000000111111", "000000111110", "000000111101", "000000111100", "000000111011", 
"000000111010", "000000111001", "000000111000", "000000110111", "000000110110", "000000110101", "000000110101", "000000110100", "000000110011", "000000110010", 
"000000110001", "000000110000", "000000101111", "000000110000", "000000110001", "000000110010", "000000110011", "000000110100", "000000110101", "000000110101", 
"000000110110", "000000110111", "000000111000", "000000111001", "000000111010", "000000111011", "000000111100", "000000111101", "000000111110", "000000111111", 
"000001000000", "000001000000", "000001000001", "000001000010", "000001000011", "000001000011", "000001000100", "000001000101", "000001000101", "000001000110", 
"000001000110", "000001000110", "000001000110", "000001000111", "000001001001", "000001001001", "000001001001", "000001001001", "000001001000", "000001001000", 
"000001001000", "000001000111", "000001000110", "000001000110", "000001000101", "000001000100", "000001000011", "000001000010", "000001000001", "000001000000", 
"000000111111", "000000111111", "000000111110", "000000111101", "000000111100", "000000111011", "000000111001", "000000111001", "000000111000", "000000110111", 
"000000110110", "000000110101", "000000110100", "000000110011", "000000110010", "000000110001", "000000110000", "000000110001", "000000110010", "000000110011", 
"000000110100", "000000110101", "000000110110", "000000110111", "000000111000", "000000111001", "000000111001", "000000111011", "000000111100", "000000111101", 
"000000111110", "000000111111", "000000111111", "000001000000", "000001000001", "000001000010", "000001000011", "000001000100", "000001000101", "000001000110", 
"000001000110", "000001000111", "000001001000", "000001001000", "000001001000", "000001001001", "000001001001", "000001001001", "000001001100", "000001001100", 
"000001001100", "000001001011", "000001001011", "000001001011", "000001001010", "000001001001", "000001001001", "000001001000", "000001000111", "000001000110", 
"000001000101", "000001000100", "000001000011", "000001000010", "000001000001", "000001000000", "000000111111", "000000111110", "000000111101", "000000111100", 
"000000111011", "000000111010", "000000111001", "000000111000", "000000110111", "000000110110", "000000110101", "000000110100", "000000110011", "000000110010", 
"000000110001", "000000110010", "000000110011", "000000110100", "000000110101", "000000110110", "000000110111", "000000111000", "000000111001", "000000111010", 
"000000111011", "000000111100", "000000111101", "000000111110", "000000111111", "000001000000", "000001000001", "000001000010", "000001000011", "000001000100", 
"000001000101", "000001000110", "000001000111", "000001001000", "000001001001", "000001001001", "000001001010", "000001001011", "000001001011", "000001001011", 
"000001001100", "000001001100", "000001001111", "000001001111", "000001001111", "000001001110", "000001001110", "000001001101", "000001001101", "000001001100", 
"000001001011", "000001001010", "000001001010", "000001001001", "000001001000", "000001000110", "000001000101", "000001000100", "000001000011", "000001000010", 
"000001000001", "000001000000", "000000111110", "000000111101", "000000111100", "000000111011", "000000111010", "000000111001", "000000111000", "000000110111", 
"000000110110", "000000110101", "000000110100", "000000110011", "000000110010", "000000110011", "000000110100", "000000110101", "000000110110", "000000110111", 
"000000111000", "000000111001", "000000111010", "000000111011", "000000111100", "000000111101", "000000111110", "000001000000", "000001000001", "000001000010", 
"000001000011", "000001000100", "000001000101", "000001000110", "000001001000", "000001001001", "000001001010", "000001001010", "000001001011", "000001001100", 
"000001001101", "000001001101", "000001001110", "000001001110", "000001001111", "000001001111", "000001010010", "000001010010", "000001010010", "000001010001", 
"000001010001", "000001010000", "000001010000", "000001001111", "000001001110", "000001001101", "000001001100", "000001001011", "000001001010", "000001001001", 
"000001000111", "000001000110", "000001000101", "000001000100", "000001000010", "000001000001", "000001000000", "000000111111", "000000111101", "000000111100", 
"000000111011", "000000111010", "000000111001", "000000111000", "000000110111", "000000110101", "000000110100", "000000110011", "000000110010", "000000110011", 
"000000110100", "000000110101", "000000110111", "000000111000", "000000111001", "000000111010", "000000111011", "000000111100", "000000111101", "000000111111", 
"000001000000", "000001000001", "000001000010", "000001000100", "000001000101", "000001000110", "000001000111", "000001001001", "000001001010", "000001001011", 
"000001001100", "000001001101", "000001001110", "000001001111", "000001010000", "000001010000", "000001010001", "000001010001", "000001010010", "000001010010", 
"000001010101", "000001010101", "000001010101", "000001010101", "000001010100", "000001010100", "000001010011", "000001010010", "000001010001", "000001010000", 
"000001001111", "000001001110", "000001001100", "000001001011", "000001001010", "000001001000", "000001000111", "000001000110", "000001000100", "000001000011", 
"000001000010", "000001000000", "000000111111", "000000111110", "000000111100", "000000111011", "000000111010", "000000111001", "000000111000", "000000110110", 
"000000110101", "000000110100", "000000110011", "000000110100", "000000110101", "000000110110", "000000111000", "000000111001", "000000111010", "000000111011", 
"000000111100", "000000111110", "000000111111", "000001000000", "000001000010", "000001000011", "000001000100", "000001000110", "000001000111", "000001001000", 
"000001001010", "000001001011", "000001001100", "000001001110", "000001001111", "000001010000", "000001010001", "000001010010", "000001010011", "000001010100", 
"000001010100", "000001010101", "000001010101", "000001010101", "000001011001", "000001011001", "000001011001", "000001011000", "000001011000", "000001010111", 
"000001010110", "000001010101", "000001010100", "000001010011", "000001010010", "000001010000", "000001001111", "000001001101", "000001001100", "000001001011", 
"000001001001", "000001001000", "000001000110", "000001000101", "000001000011", "000001000010", "000001000000", "000000111111", "000000111110", "000000111100", 
"000000111011", "000000111010", "000000111001", "000000110111", "000000110110", "000000110101", "000000110100", "000000110101", "000000110110", "000000110111", 
"000000111001", "000000111010", "000000111011", "000000111100", "000000111110", "000000111111", "000001000000", "000001000010", "000001000011", "000001000101", 
"000001000110", "000001001000", "000001001001", "000001001011", "000001001100", "000001001101", "000001001111", "000001010000", "000001010010", "000001010011", 
"000001010100", "000001010101", "000001010110", "000001010111", "000001011000", "000001011000", "000001011001", "000001011001", "000001011101", "000001011101", 
"000001011101", "000001011100", "000001011100", "000001011011", "000001011010", "000001011001", "000001010111", "000001010110", "000001010101", "000001010011", 
"000001010010", "000001010000", "000001001111", "000001001101", "000001001011", "000001001010", "000001001000", "000001000110", "000001000101", "000001000011", 
"000001000010", "000001000000", "000000111111", "000000111101", "000000111100", "000000111011", "000000111001", "000000111000", "000000110111", "000000110110", 
"000000110101", "000000110110", "000000110111", "000000111000", "000000111001", "000000111011", "000000111100", "000000111101", "000000111111", "000001000000", 
"000001000010", "000001000011", "000001000101", "000001000110", "000001001000", "000001001010", "000001001011", "000001001101", "000001001111", "000001010000", 
"000001010010", "000001010011", "000001010101", "000001010110", "000001010111", "000001011001", "000001011010", "000001011011", "000001011100", "000001011100", 
"000001011101", "000001011101", "000001100010", "000001100001", "000001100001", "000001100001", "000001100000", "000001011111", "000001011110", "000001011100", 
"000001011011", "000001011010", "000001011000", "000001010110", "000001010101", "000001010011", "000001010001", "000001001111", "000001001110", "000001001100", 
"000001001010", "000001001000", "000001000111", "000001000101", "000001000011", "000001000010", "000001000000", "000000111111", "000000111101", "000000111100", 
"000000111011", "000000111001", "000000111000", "000000110111", "000000110101", "000000110111", "000000111000", "000000111001", "000000111011", "000000111100", 
"000000111101", "000000111111", "000001000000", "000001000010", "000001000011", "000001000101", "000001000111", "000001001000", "000001001010", "000001001100", 
"000001001110", "000001001111", "000001010001", "000001010011", "000001010101", "000001010110", "000001011000", "000001011010", "000001011011", "000001011100", 
"000001011110", "000001011111", "000001100000", "000001100001", "000001100001", "000001100001", "000001100110", "000001100110", "000001100110", "000001100101", 
"000001100100", "000001100011", "000001100010", "000001100001", "000001011111", "000001011101", "000001011100", "000001011010", "000001011000", "000001010110", 
"000001010100", "000001010010", "000001010000", "000001001110", "000001001100", "000001001010", "000001001000", "000001000111", "000001000101", "000001000011", 
"000001000010", "000001000000", "000000111110", "000000111101", "000000111100", "000000111010", "000000111001", "000000111000", "000000110110", "000000111000", 
"000000111001", "000000111010", "000000111100", "000000111101", "000000111110", "000001000000", "000001000010", "000001000011", "000001000101", "000001000111", 
"000001001000", "000001001010", "000001001100", "000001001110", "000001010000", "000001010010", "000001010100", "000001010110", "000001011000", "000001011010", 
"000001011100", "000001011101", "000001011111", "000001100001", "000001100010", "000001100011", "000001100100", "000001100101", "000001100110", "000001100110", 
"000001101100", "000001101100", "000001101011", "000001101010", "000001101001", "000001101000", "000001100111", "000001100101", "000001100011", "000001100001", 
"000001011111", "000001011101", "000001011011", "000001011001", "000001010111", "000001010101", "000001010010", "000001010000", "000001001110", "000001001100", 
"000001001010", "000001001000", "000001000110", "000001000101", "000001000011", "000001000001", "000001000000", "000000111110", "000000111101", "000000111011", 
"000000111010", "000000111000", "000000110111", "000000111000", "000000111010", "000000111011", "000000111101", "000000111110", "000001000000", "000001000001", 
"000001000011", "000001000101", "000001000110", "000001001000", "000001001010", "000001001100", "000001001110", "000001010000", "000001010010", "000001010101", 
"000001010111", "000001011001", "000001011011", "000001011101", "000001011111", "000001100001", "000001100011", "000001100101", "000001100111", "000001101000", 
"000001101001", "000001101010", "000001101011", "000001101100", "000001110010", "000001110010", "000001110001", "000001110000", "000001101111", "000001101110", 
"000001101100", "000001101010", "000001101000", "000001100110", "000001100011", "000001100001", "000001011111", "000001011100", "000001011010", "000001010111", 
"000001010101", "000001010011", "000001010000", "000001001110", "000001001100", "000001001010", "000001001000", "000001000110", "000001000100", "000001000010", 
"000001000001", "000000111111", "000000111110", "000000111100", "000000111011", "000000111001", "000000111000", "000000111001", "000000111011", "000000111100", 
"000000111110", "000000111111", "000001000001", "000001000010", "000001000100", "000001000110", "000001001000", "000001001010", "000001001100", "000001001110", 
"000001010000", "000001010011", "000001010101", "000001010111", "000001011010", "000001011100", "000001011111", "000001100001", "000001100011", "000001100110", 
"000001101000", "000001101010", "000001101100", "000001101110", "000001101111", "000001110000", "000001110001", "000001110010", "000001111000", "000001111000", 
"000001111000", "000001110111", "000001110101", "000001110100", "000001110010", "000001101111", "000001101101", "000001101010", "000001101000", "000001100101", 
"000001100010", "000001100000", "000001011101", "000001011010", "000001011000", "000001010101", "000001010011", "000001010000", "000001001110", "000001001100", 
"000001001010", "000001001000", "000001000110", "000001000100", "000001000010", "000001000000", "000000111111", "000000111101", "000000111011", "000000111010", 
"000000111001", "000000111010", "000000111011", "000000111101", "000000111111", "000001000000", "000001000010", "000001000100", "000001000110", "000001001000", 
"000001001010", "000001001100", "000001001110", "000001010000", "000001010011", "000001010101", "000001011000", "000001011010", "000001011101", "000001100000", 
"000001100010", "000001100101", "000001101000", "000001101010", "000001101101", "000001101111", "000001110010", "000001110100", "000001110101", "000001110111", 
"000001111000", "000001111000", "000010000000", "000010000000", "000001111111", "000001111110", "000001111100", "000001111010", "000001111000", "000001110101", 
"000001110010", "000001110000", "000001101101", "000001101001", "000001100110", "000001100011", "000001100000", "000001011101", "000001011010", "000001011000", 
"000001010101", "000001010010", "000001010000", "000001001110", "000001001011", "000001001001", "000001000111", "000001000101", "000001000011", "000001000001", 
"000000111111", "000000111110", "000000111100", "000000111011", "000000111001", "000000111011", "000000111100", "000000111110", "000000111111", "000001000001", 
"000001000011", "000001000101", "000001000111", "000001001001", "000001001011", "000001001110", "000001010000", "000001010010", "000001010101", "000001011000", 
"000001011010", "000001011101", "000001100000", "000001100011", "000001100110", "000001101001", "000001101101", "000001110000", "000001110010", "000001110101", 
"000001111000", "000001111010", "000001111100", "000001111110", "000001111111", "000010000000", "000010001001", "000010001000", "000010000111", "000010000110", 
"000010000100", "000010000001", "000001111111", "000001111100", "000001111000", "000001110101", "000001110010", "000001101110", "000001101011", "000001100111", 
"000001100100", "000001100001", "000001011101", "000001011010", "000001010111", "000001010101", "000001010010", "000001001111", "000001001101", "000001001011", 
"000001001000", "000001000110", "000001000100", "000001000010", "000001000000", "000000111111", "000000111101", "000000111011", "000000111010", "000000111011", 
"000000111101", "000000111111", "000001000000", "000001000010", "000001000100", "000001000110", "000001001000", "000001001011", "000001001101", "000001001111", 
"000001010010", "000001010101", "000001010111", "000001011010", "000001011101", "000001100001", "000001100100", "000001100111", "000001101011", "000001101110", 
"000001110010", "000001110101", "000001111000", "000001111100", "000001111111", "000010000001", "000010000100", "000010000110", "000010000111", "000010001000", 
"000010010010", "000010010010", "000010010001", "000010001111", "000010001101", "000010001010", "000010000110", "000010000011", "000001111111", "000001111011", 
"000001110111", "000001110011", "000001101111", "000001101011", "000001100111", "000001100100", "000001100000", "000001011101", "000001011010", "000001010111", 
"000001010100", "000001010001", "000001001111", "000001001100", "000001001010", "000001000111", "000001000101", "000001000011", "000001000001", "000001000000", 
"000000111110", "000000111100", "000000111011", "000000111100", "000000111110", "000001000000", "000001000001", "000001000011", "000001000101", "000001000111", 
"000001001010", "000001001100", "000001001111", "000001010001", "000001010100", "000001010111", "000001011010", "000001011101", "000001100000", "000001100100", 
"000001100111", "000001101011", "000001101111", "000001110011", "000001110111", "000001111011", "000001111111", "000010000011", "000010000110", "000010001010", 
"000010001101", "000010001111", "000010010001", "000010010010", "000010011110", "000010011101", "000010011100", "000010011001", "000010010111", "000010010011", 
"000010001111", "000010001011", "000010000110", "000010000001", "000001111101", "000001111000", "000001110100", "000001101111", "000001101011", "000001100111", 
"000001100011", "000001100000", "000001011100", "000001011001", "000001010110", "000001010011", "000001010000", "000001001101", "000001001011", "000001001001", 
"000001000110", "000001000100", "000001000010", "000001000000", "000000111111", "000000111101", "000000111011", "000000111101", "000000111111", "000001000000", 
"000001000010", "000001000100", "000001000110", "000001001001", "000001001011", "000001001101", "000001010000", "000001010011", "000001010110", "000001011001", 
"000001011100", "000001100000", "000001100011", "000001100111", "000001101011", "000001101111", "000001110100", "000001111000", "000001111101", "000010000001", 
"000010000110", "000010001011", "000010001111", "000010010011", "000010010111", "000010011001", "000010011100", "000010011101", "000010101011", "000010101010", 
"000010101000", "000010100110", "000010100010", "000010011110", "000010011001", "000010010011", "000010001110", "000010001001", "000010000011", "000001111110", 
"000001111001", "000001110100", "000001101111", "000001101011", "000001100110", "000001100010", "000001011111", "000001011011", "000001011000", "000001010101", 
"000001010010", "000001001111", "000001001100", "000001001010", "000001001000", "000001000101", "000001000011", "000001000001", "000000111111", "000000111110", 
"000000111100", "000000111110", "000000111111", "000001000001", "000001000011", "000001000101", "000001001000", "000001001010", "000001001100", "000001001111", 
"000001010010", "000001010101", "000001011000", "000001011011", "000001011111", "000001100010", "000001100110", "000001101011", "000001101111", "000001110100", 
"000001111001", "000001111110", "000010000011", "000010001001", "000010001110", "000010010011", "000010011001", "000010011110", "000010100010", "000010100110", 
"000010101000", "000010101010", "000010111010", "000010111001", "000010110111", "000010110100", "000010101111", "000010101001", "000010100011", "000010011101", 
"000010010111", "000010010000", "000010001010", "000010000100", "000001111110", "000001111000", "000001110011", "000001101110", "000001101001", "000001100101", 
"000001100001", "000001011101", "000001011010", "000001010110", "000001010011", "000001010000", "000001001110", "000001001011", "000001001001", "000001000110", 
"000001000100", "000001000010", "000001000000", "000000111110", "000000111101", "000000111110", "000001000000", "000001000010", "000001000100", "000001000110", 
"000001001001", "000001001011", "000001001110", "000001010000", "000001010011", "000001010110", "000001011010", "000001011101", "000001100001", "000001100101", 
"000001101001", "000001101110", "000001110011", "000001111000", "000001111110", "000010000100", "000010001010", "000010010000", "000010010111", "000010011101", 
"000010100011", "000010101001", "000010101111", "000010110100", "000010110111", "000010111001", "000011001101", "000011001100", "000011001001", "000011000100", 
"000010111110", "000010110111", "000010110000", "000010101000", "000010100000", "000010011000", "000010010001", "000010001010", "000010000011", "000001111101", 
"000001110111", "000001110010", "000001101101", "000001101000", "000001100011", "000001011111", "000001011100", "000001011000", "000001010101", "000001010010", 
"000001001111", "000001001100", "000001001010", "000001000111", "000001000101", "000001000011", "000001000001", "000000111111", "000000111101", "000000111111", 
"000001000001", "000001000011", "000001000101", "000001000111", "000001001010", "000001001100", "000001001111", "000001010010", "000001010101", "000001011000", 
"000001011100", "000001011111", "000001100011", "000001101000", "000001101101", "000001110010", "000001110111", "000001111101", "000010000011", "000010001010", 
"000010010001", "000010011000", "000010100000", "000010101000", "000010110000", "000010110111", "000010111110", "000011000100", "000011001001", "000011001100", 
"000011100100", "000011100010", "000011011110", "000011011000", "000011010000", "000011000111", "000010111101", "000010110100", "000010101010", "000010100001", 
"000010011000", "000010010000", "000010001001", "000010000001", "000001111011", "000001110101", "000001110000", "000001101010", "000001100110", "000001100001", 
"000001011101", "000001011010", "000001010110", "000001010011", "000001010000", "000001001101", "000001001010", "000001001000", "000001000110", "000001000011", 
"000001000001", "000000111111", "000000111110", "000000111111", "000001000001", "000001000011", "000001000110", "000001001000", "000001001010", "000001001101", 
"000001010000", "000001010011", "000001010110", "000001011010", "000001011101", "000001100001", "000001100110", "000001101010", "000001110000", "000001110101", 
"000001111011", "000010000001", "000010001001", "000010010000", "000010011000", "000010100001", "000010101010", "000010110100", "000010111101", "000011000111", 
"000011010000", "000011011000", "000011011110", "000011100010", "000100000000", "000011111110", "000011111000", "000011110000", "000011100101", "000011011001", 
"000011001101", "000011000001", "000010110101", "000010101010", "000010100000", "000010010111", "000010001110", "000010000110", "000001111111", "000001111000", 
"000001110010", "000001101101", "000001101000", "000001100011", "000001011111", "000001011011", "000001010111", "000001010100", "000001010001", "000001001110", 
"000001001011", "000001001001", "000001000110", "000001000100", "000001000010", "000001000000", "000000111110", "000001000000", "000001000010", "000001000100", 
"000001000110", "000001001001", "000001001011", "000001001110", "000001010001", "000001010100", "000001010111", "000001011011", "000001011111", "000001100011", 
"000001101000", "000001101101", "000001110010", "000001111000", "000001111111", "000010000110", "000010001110", "000010010111", "000010100000", "000010101010", 
"000010110101", "000011000001", "000011001101", "000011011001", "000011100101", "000011110000", "000011111000", "000011111110", "000100100101", "000100100010", 
"000100011001", "000100001101", "000011111110", "000011101110", "000011011110", "000011001111", "000011000001", "000010110100", "000010101000", "000010011101", 
"000010010011", "000010001011", "000010000011", "000001111100", "000001110101", "000001101111", "000001101010", "000001100101", "000001100001", "000001011100", 
"000001011001", "000001010101", "000001010010", "000001001111", "000001001100", "000001001001", "000001000111", "000001000101", "000001000010", "000001000000", 
"000000111111", "000001000000", "000001000010", "000001000101", "000001000111", "000001001001", "000001001100", "000001001111", "000001010010", "000001010101", 
"000001011001", "000001011100", "000001100001", "000001100101", "000001101010", "000001101111", "000001110101", "000001111100", "000010000011", "000010001011", 
"000010010011", "000010011101", "000010101000", "000010110100", "000011000001", "000011001111", "000011011110", "000011101110", "000011111110", "000100001101", 
"000100011001", "000100100010", "000101010101", "000101010001", "000101000100", "000100110001", "000100011100", "000100000110", "000011110001", "000011011110", 
"000011001101", "000010111101", "000010110000", "000010100011", "000010011001", "000010001111", "000010000110", "000001111111", "000001111000", "000001110010", 
"000001101100", "000001100111", "000001100010", "000001011110", "000001011010", "000001010110", "000001010011", "000001010000", "000001001101", "000001001010", 
"000001001000", "000001000101", "000001000011", "000001000001", "000000111111", "000001000001", "000001000011", "000001000101", "000001001000", "000001001010", 
"000001001101", "000001010000", "000001010011", "000001010110", "000001011010", "000001011110", "000001100010", "000001100111", "000001101100", "000001110010", 
"000001111000", "000001111111", "000010000110", "000010001111", "000010011001", "000010100011", "000010110000", "000010111101", "000011001101", "000011011110", 
"000011110001", "000100000110", "000100011100", "000100110001", "000101000100", "000101010001", "000110011010", "000110010010", "000101111100", "000101011111", 
"000101000000", "000100100010", "000100000110", "000011101110", "000011011001", "000011000111", "000010110111", "000010101001", "000010011110", "000010010011", 
"000010001010", "000010000001", "000001111010", "000001110100", "000001101110", "000001101000", "000001100011", "000001011111", "000001011011", "000001010111", 
"000001010100", "000001010000", "000001001101", "000001001011", "000001001000", "000001000110", "000001000011", "000001000001", "000000111111", "000001000001", 
"000001000011", "000001000110", "000001001000", "000001001011", "000001001101", "000001010000", "000001010100", "000001010111", "000001011011", "000001011111", 
"000001100011", "000001101000", "000001101110", "000001110100", "000001111010", "000010000001", "000010001010", "000010010011", "000010011110", "000010101001", 
"000010110111", "000011000111", "000011011001", "000011101110", "000100000110", "000100100010", "000101000000", "000101011111", "000101111100", "000110010010", 
"001000000000", "000111110001", "000111001010", "000110011010", "000101101010", "000101000000", "000100011100", "000011111110", "000011100101", "000011010000", 
"000010111110", "000010101111", "000010100010", "000010010111", "000010001101", "000010000100", "000001111100", "000001110101", "000001101111", "000001101001", 
"000001100100", "000001100000", "000001011100", "000001011000", "000001010100", "000001010001", "000001001110", "000001001011", "000001001000", "000001000110", 
"000001000100", "000001000010", "000000111111", "000001000010", "000001000100", "000001000110", "000001001000", "000001001011", "000001001110", "000001010001", 
"000001010100", "000001011000", "000001011100", "000001100000", "000001100100", "000001101001", "000001101111", "000001110101", "000001111100", "000010000100", 
"000010001101", "000010010111", "000010100010", "000010101111", "000010111110", "000011010000", "000011100101", "000011111110", "000100011100", "000101000000", 
"000101101010", "000110011010", "000111001010", "000111110001", "001010101011", "001010000111", "001000111000", "000111100011", "000110011010", "000101011111", 
"000100110001", "000100001101", "000011110000", "000011011000", "000011000100", "000010110100", "000010100110", "000010011001", "000010001111", "000010000110", 
"000001111110", "000001110111", "000001110000", "000001101010", "000001100101", "000001100001", "000001011100", "000001011000", "000001010101", "000001010001", 
"000001001110", "000001001011", "000001001001", "000001000110", "000001000100", "000001000010", "000001000000", "000001000010", "000001000100", "000001000110", 
"000001001001", "000001001011", "000001001110", "000001010001", "000001010101", "000001011000", "000001011100", "000001100001", "000001100101", "000001101010", 
"000001110000", "000001110111", "000001111110", "000010000110", "000010001111", "000010011001", "000010100110", "000010110100", "000011000100", "000011011000", 
"000011110000", "000100001101", "000100110001", "000101011111", "000110011010", "000111100011", "001000111000", "001010000111", "010000000000", "001110010100", 
"001011010100", "001000111000", "000111001010", "000101111100", "000101000100", "000100011001", "000011111000", "000011011110", "000011001001", "000010110111", 
"000010101000", "000010011100", "000010010001", "000010000111", "000001111111", "000001111000", "000001110001", "000001101011", "000001100110", "000001100001", 
"000001011101", "000001011001", "000001010101", "000001010010", "000001001111", "000001001100", "000001001001", "000001000110", "000001000100", "000001000010", 
"000001000000", "000001000010", "000001000100", "000001000110", "000001001001", "000001001100", "000001001111", "000001010010", "000001010101", "000001011001", 
"000001011101", "000001100001", "000001100110", "000001101011", "000001110001", "000001111000", "000001111111", "000010000111", "000010010001", "000010011100", 
"000010101000", "000010110111", "000011001001", "000011011110", "000011111000", "000100011001", "000101000100", "000101111100", "000111001010", "001000111000", 
"001011010100", "001110010100", "100000000000", "010110101000", "001110010100", "001010000111", "000111110001", "000110010010", "000101010001", "000100100010", 
"000011111110", "000011100010", "000011001100", "000010111001", "000010101010", "000010011101", "000010010010", "000010001000", "000010000000", "000001111000", 
"000001110010", "000001101100", "000001100110", "000001100001", "000001011101", "000001011001", "000001010101", "000001010010", "000001001111", "000001001100", 
"000001001001", "000001000111", "000001000100", "000001000010", "000001000000", "000001000010", "000001000100", "000001000111", "000001001001", "000001001100", 
"000001001111", "000001010010", "000001010101", "000001011001", "000001011101", "000001100001", "000001100110", "000001101100", "000001110010", "000001111000", 
"000010000000", "000010001000", "000010010010", "000010011101", "000010101010", "000010111001", "000011001100", "000011100010", "000011111110", "000100100010", 
"000101010001", "000110010010", "000111110001", "001010000111", "001110010100", "010110101000" );




constant BITSIZE:integer:=8;
constant SH:integer:=3;

signal mulval_a:std_logic_vector(NORMBITOUT-1 downto 0):=(others=>'0');
signal acum_re_1w,acum_im_1w,acum_re_new,acum_im_new,acum_re,acum_im,sample_rotI,sample_rotQ:std_logic_vector(15 downto 0);
signal acum_re_mula,acum_im_mula:std_logic_vector(15+NORMBITOUT+1 downto 0):=(others=>'0');
signal table_re,table_im,to_tab_re,to_tab_im:std_logic_vector(BITSIZE-1 downto 0);
signal table_reE,table_imE:std_logic_vector(15 downto 0);
signal ce_1w,ce_table,ce_acum,shift1,shift2:std_logic;
signal poval:std_logic_vector(NORMBIT*2-1 downto 0);


--signal poval:std_logic_vector(NORM_LEN-1 downto 0);

signal povval_x,povval_y:std_logic_vector(NORMBIT-1 downto 0);

begin

SIM01: if SIMULATION=1 generate
--	save_complexdata_i: entity work.save_complexdata
--		port map(
--		clk =>clk,
--		i_ce =>i_ce,
--		i_samplesI=>i_samplesI,
--		i_samplesQ=>i_samplesQ,
--
--		i_ce2 =>after_pilot_start,
--		i_samplesI2=>i_init_phaseI,
--		i_samplesQ2=>i_init_phaseQ
--		);
end generate;


table_reE<=table_re&EXT("0",16-BITSIZE);
table_imE<=table_im&EXT("0",16-BITSIZE);

complex_mult_q_i: entity work.complex_mult_q
	generic map(
		SHIFT_MUL=>1,
		CONJUGATION=>'1' --# ��������� �� ����������� �����, ���� '1' - �� ���������
	)
	port map(
		clk =>clk,
		i_ce =>i_ce,

		A_I=>i_samplesI,
		B_Q=>i_samplesQ,

		C_I=>acum_re,
		D_Q=>acum_im,

		o_I=>sample_rotI,
		o_Q=>sample_rotQ,
		out_ce=>open
		);

complex_mult_q_ii: entity work.complex_mult_qr
	generic map(
		SHIFT_MUL=>3, --# (����� ������� ��� 3)
		CONJUGATION=>'0' --# ��������� �� ����������� �����, ���� '1' - �� ���������
	)
	port map(
		clk =>clk,

		load =>after_pilot_start,

		init_I=>i_init_phaseI,
		init_Q=>i_init_phaseQ,

		i_ce =>ce_table,
		A_I=>acum_re_1w,       --# 6101+1i*1157  (�����)
		B_Q=>acum_im_1w,


		C_I=>table_reE,        --# 32256-1i*4352 (�����)
		D_Q=>table_imE,

		o_I=>acum_re_new, --# ��� ���������� ������������ ������ ���� 12318+1i*656
		o_Q=>acum_im_new,
		out_ce=>ce_acum
		);

shift1<='1' when unsigned(signed_abs(sample_rotI(sample_rotI'Length-1 downto 6)))>127 or unsigned(signed_abs(sample_rotQ(sample_rotQ'Length-1 downto 6)))>127  else '0';

--to_tab_re<=SXT(sample_rotI(sample_rotI'Length-1 downto 9),BITSIZE) when 
--	unsigned(signed_abs(sample_rotI(sample_rotI'Length-1 downto 6)))>127 or unsigned(signed_abs(sample_rotQ(sample_rotQ'Length-1 downto 6)))>127 
--	else sample_rotI(6+BITSIZE-1 downto 6);

--to_tab_im<=SXT(sample_rotQ(sample_rotQ'Length-1 downto 9),BITSIZE) when 
--	unsigned(signed_abs(sample_rotI(sample_rotI'Length-1 downto 6)))>127 or unsigned(signed_abs(sample_rotQ(sample_rotQ'Length-1 downto 6)))>127 
--	else sample_rotQ(6+BITSIZE-1 downto 6);

--to_tab_re<=sample_rotI(5+BITSIZE-1 downto 5); --# !!!was
--to_tab_im<=sample_rotQ(5+BITSIZE-1 downto 5);


to_tab_re<=sample_rotI(sample_rotI'Length-1 downto sample_rotI'Length-BITSIZE);
to_tab_im<=sample_rotQ(sample_rotI'Length-1 downto sample_rotI'Length-BITSIZE);


--to_tab_re<=norming(sample_rotI(5+BITSIZE-1 downto 5),sample_rotI(5+BITSIZE-1 downto 5),sample_rotQ(5+BITSIZE-1 downto 5),8192.0);
--to_tab_im<=norming(sample_rotQ(5+BITSIZE-1 downto 5),sample_rotI(5+BITSIZE-1 downto 5),sample_rotQ(5+BITSIZE-1 downto 5),8192.0);


table_demod_i:entity work.table_demod
	generic map(
		BIT_IN=>BITSIZE,
		BIT_OUT=>BITSIZE
	)
	 port map(
		  clk =>clk,
		  i_ce=>ce_1w,
	      sample_in_re=>to_tab_re,
	      sample_in_im=>to_tab_im,
		  o_ce=>ce_table,
	      sample_out_re=>table_re,
	      sample_out_im=>table_im
		 );
		




povval_x<=acum_re_new(acum_re_new'Length-1 downto acum_re_new'Length-NORMBIT);  --# was
povval_y<=acum_im_new(acum_re_new'Length-1 downto acum_re_new'Length-NORMBIT);





--poval<=acum_im_new(acum_re_new'Length-1-1 downto acum_re_new'Length-NORMBIT-1)&acum_re_new(acum_re_new'Length-1-1 downto acum_re_new'Length-NORMBIT-1);
poval<=acum_im_new(acum_re_new'Length-1 downto acum_re_new'Length-NORMBIT)&acum_re_new(acum_re_new'Length-1 downto acum_re_new'Length-NORMBIT);
mulval_a<=norm_mem(conv_integer(acum_im_new(acum_re_new'Length-1 downto acum_re_new'Length-NORMBIT)&acum_re_new(acum_re_new'Length-1 downto acum_re_new'Length-NORMBIT)));

process(clk) is
variable v_acum_re_mula,v_acum_im_mula:std_logic_vector(acum_re_mula'Length-1 downto 0):=(others=>'0');

begin
	if rising_edge(clk) then
		ce_1w<=i_ce;
		out_ce<=i_ce;


--o_samplesI<=norming(sample_rotI,sample_rotI,sample_rotQ,8192.0);
--o_samplesQ<=norming(sample_rotQ,sample_rotI,sample_rotQ,8192.0);


--o_samplesI<=conv_std_logic_vector( integer(8192.0*real(conv_integer(signed(sample_rotI)))/sqrt(real(conv_integer(signed(sample_rotI)))*real(conv_integer(signed(sample_rotI)))+real(conv_integer(signed(sample_rotQ)))*real(conv_integer(signed(sample_rotQ))) )), o_samplesI'Length);
--o_samplesQ<=conv_std_logic_vector( integer(8192.0*real(conv_integer(signed(sample_rotQ)))/sqrt(real(conv_integer(signed(sample_rotI)))*real(conv_integer(signed(sample_rotI)))+real(conv_integer(signed(sample_rotQ)))*real(conv_integer(signed(sample_rotQ))) )), o_samplesI'Length);

		o_samplesI<=sample_rotI;
		o_samplesQ<=sample_rotQ;

--			acum_re_1w<=i_init_phaseI;
--			acum_im_1w<=i_init_phaseQ;

		if after_pilot_start='1' then
				acum_re_1w<=i_init_phaseI;
				acum_im_1w<=i_init_phaseQ;
--				acum_re_1w<=norming(i_init_phaseI,i_init_phaseI,i_init_phaseQ,8192.0);
--				acum_im_1w<=norming(i_init_phaseQ,i_init_phaseI,i_init_phaseQ,8192.0);

		else
				acum_re_1w<=acum_re;
				acum_im_1w<=acum_im;
		end if;

--		if after_pilot_start='1' then
--			acum_re<=(others=>'0');--i_init_phaseI;
--			acum_im<=(others=>'0');--i_init_phaseQ;
--		else        --# reset
--			if ce_acum='1' then



				v_acum_re_mula:=signed(acum_re_new)*unsigned(mulval_a);
				v_acum_im_mula:=signed(acum_im_new)*unsigned(mulval_a);

				acum_re_mula<=signed(acum_re_new)*unsigned(mulval_a);
				acum_im_mula<=signed(acum_im_new)*unsigned(mulval_a);

--# was
--				acum_re<=v_acum_re_mula(acum_re_mula'Length-1-(NORMBIT-1) downto acum_re_mula'Length-acum_re'Length-(NORMBIT-1));
--				acum_im<=v_acum_im_mula(acum_re_mula'Length-1-(NORMBIT-1) downto acum_re_mula'Length-acum_re'Length-(NORMBIT-1));

				acum_re<=SXT(v_acum_re_mula(acum_re_mula'Length-1-NORMBIT downto acum_re_mula'Length-acum_re'Length-NORMBIT+1),acum_re'Length);
				acum_im<=SXT(v_acum_im_mula(acum_re_mula'Length-1-NORMBIT downto acum_re_mula'Length-acum_re'Length-NORMBIT+1),acum_im'Length);



--				acum_re<=norming(acum_re_new,acum_re_new,acum_im_new,8192.0);
--				acum_im<=norming(acum_im_new,acum_re_new,acum_im_new,8192.0);


--				acum_re<=conv_std_logic_vector( integer(8192.0*real(conv_integer(signed(acum_re_new)))/sqrt(real(conv_integer(signed(acum_re_new)))*real(conv_integer(signed(acum_re_new)))+real(conv_integer(signed(acum_im_new)))*real(conv_integer(signed(acum_im_new))) )), acum_re'Length);
--				acum_im<=conv_std_logic_vector( integer(8192.0*real(conv_integer(signed(acum_im_new)))/sqrt(real(conv_integer(signed(acum_re_new)))*real(conv_integer(signed(acum_re_new)))+real(conv_integer(signed(acum_im_new)))*real(conv_integer(signed(acum_im_new))) )), acum_re'Length);



--			end if; --# i_ce
--		end if;     --# reset
	end if;
end process;



end average_itertive_demod;



