library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
library work;
use work.feedf_consts_pack.all;


entity qcomplex_norm is
	port(
		clk : in STD_LOGIC;
		i_ce : in std_logic;		
		i_samplesI: in std_logic_vector(15 downto 0);
		i_samplesQ: in std_logic_vector(15 downto 0);

		o_ce : out std_logic;		
		o_samplesI: out std_logic_vector(15 downto 0);
		o_samplesQ: out std_logic_vector(15 downto 0)
		);
end qcomplex_norm;



architecture qcomplex_norm of qcomplex_norm is

constant NORMBIT:natural:=5;
constant NORMBITOUT:natural:=8;

type Tnorm_mem is array (0 to 1023) of std_logic_vector(7 downto 0);
constant norm_mem:Tnorm_mem:=  (
"11111111", 
"11111111", "10000000", "01010101", "01000000", "00110011", "00101011", "00100100", "00100000", "00011100", "00011010", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00010001", "00010010", "00010100", "00010101", 
"00010111", "00011010", "00011100", "00100000", "00100100", "00101011", "00110011", "01000000", "01010101", "10000000", "11111111", "11111111", "10110100", "01110010", "01010001", "00111110", "00110010", "00101010", "00100100", "00100000", 
"00011100", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00010001", "00010010", "00010100", "00010101", "00010111", "00011001", "00011100", "00100000", "00100100", "00101010", "00110010", "00111110", 
"01010001", "01110010", "10110100", "10000000", "01110010", "01011010", "01000111", "00111001", "00101111", "00101000", "00100011", "00011111", "00011100", "00011001", "00010111", "00010101", "00010011", "00010010", "00010001", "00010000", 
"00010001", "00010010", "00010011", "00010101", "00010111", "00011001", "00011100", "00011111", "00100011", "00101000", "00101111", "00111001", "01000111", "01011010", "01110010", "01010101", "01010001", "01000111", "00111100", "00110011", 
"00101100", "00100110", "00100001", "00011110", "00011011", "00011000", "00010110", "00010101", "00010011", "00010010", "00010001", "00010000", "00010001", "00010010", "00010011", "00010101", "00010110", "00011000", "00011011", "00011110", 
"00100001", "00100110", "00101100", "00110011", "00111100", "01000111", "01010001", "01000000", "00111110", "00111001", "00110011", "00101101", "00101000", "00100011", "00100000", "00011101", "00011010", "00011000", "00010110", "00010100", 
"00010011", "00010010", "00010000", "00001111", "00010000", "00010010", "00010011", "00010100", "00010110", "00011000", "00011010", "00011101", "00100000", "00100011", "00101000", "00101101", "00110011", "00111001", "00111110", "00110011", 
"00110010", "00101111", "00101100", "00101000", "00100100", "00100001", "00011110", "00011011", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", "00010000", "00010001", "00010010", "00010100", 
"00010101", "00010111", "00011001", "00011011", "00011110", "00100001", "00100100", "00101000", "00101100", "00101111", "00110010", "00101011", "00101010", "00101000", "00100110", "00100011", "00100001", "00011110", "00011100", "00011010", 
"00011000", "00010110", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010110", "00011000", "00011010", "00011100", "00011110", "00100001", "00100011", 
"00100110", "00101000", "00101010", "00100100", "00100100", "00100011", "00100001", "00100000", "00011110", "00011100", "00011010", "00011000", "00010110", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", "00001111", 
"00001111", "00010000", "00010001", "00010010", "00010100", "00010101", "00010110", "00011000", "00011010", "00011100", "00011110", "00100000", "00100001", "00100011", "00100100", "00100000", "00100000", "00011111", "00011110", "00011101", 
"00011011", "00011010", "00011000", "00010111", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010111", 
"00011000", "00011010", "00011011", "00011101", "00011110", "00011111", "00100000", "00011100", "00011100", "00011100", "00011011", "00011010", "00011001", "00011000", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", 
"00010000", "00001111", "00001111", "00001110", "00001111", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00011000", "00011001", "00011010", "00011011", "00011100", "00011100", "00011010", 
"00011001", "00011001", "00011000", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001110", "00001111", "00010000", "00010000", 
"00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011000", "00011001", "00011001", "00010111", "00010111", "00010111", "00010110", "00010110", "00010101", "00010100", "00010100", "00010011", 
"00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", "00010010", "00010011", "00010100", "00010100", "00010101", "00010110", 
"00010110", "00010111", "00010111", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", "00010011", "00010010", "00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001101", 
"00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", "00010010", "00010010", "00010011", "00010100", "00010100", "00010101", "00010101", "00010101", "00010100", "00010100", "00010011", "00010011", "00010011", 
"00010010", "00010010", "00010001", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", 
"00010001", "00010010", "00010010", "00010011", "00010011", "00010011", "00010100", "00010010", "00010010", "00010010", "00010010", "00010010", "00010001", "00010001", "00010000", "00010000", "00001111", "00001111", "00001110", "00001110", 
"00001101", "00001101", "00001100", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00001111", "00010000", "00010000", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010001", 
"00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001100", "00001100", "00001100", "00001101", "00001101", 
"00001110", "00001110", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001111", "00001110", 
"00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001100", "00001011", "00001100", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", 
"00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001100", 
"00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010010", 
"00010001", "00010001", "00010000", "00010000", "00001111", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00001111", "00010000", 
"00010000", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010100", "00010100", "00010011", "00010011", "00010011", "00010010", "00010010", "00010001", "00010001", "00010000", "00010000", "00001111", "00001110", 
"00001110", "00001101", "00001101", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", "00010001", "00010010", "00010010", "00010011", "00010011", "00010011", "00010100", "00010101", 
"00010101", "00010101", "00010101", "00010100", "00010100", "00010011", "00010010", "00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001101", "00001101", "00001110", "00001110", "00001111", 
"00010000", "00010000", "00010001", "00010010", "00010010", "00010011", "00010100", "00010100", "00010101", "00010101", "00010101", "00010111", "00010111", "00010111", "00010110", "00010110", "00010101", "00010100", "00010100", "00010011", 
"00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", "00010010", "00010011", "00010100", "00010100", "00010101", "00010110", 
"00010110", "00010111", "00010111", "00011010", "00011001", "00011001", "00011000", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", 
"00001110", "00001111", "00010000", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011000", "00011001", "00011001", "00011100", "00011100", "00011100", "00011011", "00011010", 
"00011001", "00011000", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001111", "00001110", "00001111", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", 
"00010110", "00011000", "00011001", "00011010", "00011011", "00011100", "00011100", "00100000", "00100000", "00011111", "00011110", "00011101", "00011011", "00011010", "00011000", "00010111", "00010101", "00010100", "00010011", "00010010", 
"00010001", "00010000", "00001111", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010111", "00011000", "00011010", "00011011", "00011101", "00011110", "00011111", "00100000", "00100100", 
"00100100", "00100011", "00100001", "00100000", "00011110", "00011100", "00011010", "00011000", "00010110", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", "00001111", "00001111", "00010000", "00010001", "00010010", 
"00010100", "00010101", "00010110", "00011000", "00011010", "00011100", "00011110", "00100000", "00100001", "00100011", "00100100", "00101011", "00101010", "00101000", "00100110", "00100011", "00100001", "00011110", "00011100", "00011010", 
"00011000", "00010110", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010110", "00011000", "00011010", "00011100", "00011110", "00100001", "00100011", 
"00100110", "00101000", "00101010", "00110011", "00110010", "00101111", "00101100", "00101000", "00100100", "00100001", "00011110", "00011011", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", 
"00010000", "00010001", "00010010", "00010100", "00010101", "00010111", "00011001", "00011011", "00011110", "00100001", "00100100", "00101000", "00101100", "00101111", "00110010", "01000000", "00111110", "00111001", "00110011", "00101101", 
"00101000", "00100011", "00100000", "00011101", "00011010", "00011000", "00010110", "00010100", "00010011", "00010010", "00010000", "00001111", "00010000", "00010010", "00010011", "00010100", "00010110", "00011000", "00011010", "00011101", 
"00100000", "00100011", "00101000", "00101101", "00110011", "00111001", "00111110", "01010101", "01010001", "01000111", "00111100", "00110011", "00101100", "00100110", "00100001", "00011110", "00011011", "00011000", "00010110", "00010101", 
"00010011", "00010010", "00010001", "00010000", "00010001", "00010010", "00010011", "00010101", "00010110", "00011000", "00011011", "00011110", "00100001", "00100110", "00101100", "00110011", "00111100", "01000111", "01010001", "10000000", 
"01110010", "01011010", "01000111", "00111001", "00101111", "00101000", "00100011", "00011111", "00011100", "00011001", "00010111", "00010101", "00010011", "00010010", "00010001", "00010000", "00010001", "00010010", "00010011", "00010101", 
"00010111", "00011001", "00011100", "00011111", "00100011", "00101000", "00101111", "00111001", "01000111", "01011010", "01110010", "11111111", "10110100", "01110010", "01010001", "00111110", "00110010", "00101010", "00100100", "00100000", 
"00011100", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00010001", "00010010", "00010100", "00010101", "00010111", "00011001", "00011100", "00100000", "00100100", "00101010", "00110010", "00111110", 
"01010001", "01110010", "10110100" );


signal ce_1w,ce_2w:std_logic;
signal mulval_a:std_logic_vector(NORMBITOUT-1 downto 0):=(others=>'0');
signal samplesI_1w,samplesQ_1w:std_logic_vector(i_samplesI'Length-1 downto 0);
signal acum_re_mula,acum_im_mula:std_logic_vector(15+NORMBITOUT+1 downto 0):=(others=>'0');

begin

process (clk) is
begin		
	if rising_edge(clk) then

		ce_1w<=i_ce;
		ce_2w<=ce_1w;

		if i_ce='1' then
		    mulval_a<=norm_mem(conv_integer(i_samplesI(i_samplesI'Length-1-1 downto i_samplesI'Length-NORMBIT-1)&i_samplesQ(i_samplesQ'Length-1-1 downto i_samplesQ'Length-NORMBIT-1)));
			samplesI_1w<=i_samplesI;
			samplesQ_1w<=i_samplesQ;
		end if;
		
		if ce_1w='1' then
			acum_re_mula<=signed(samplesI_1w)*unsigned(mulval_a);
			acum_im_mula<=signed(samplesQ_1w)*unsigned(mulval_a);
		end if;

		o_ce<=ce_2w;
		o_samplesI<=acum_re_mula(acum_re_mula'Length-1-NORMBIT downto acum_re_mula'Length-o_samplesI'Length-NORMBIT);
		o_samplesQ<=acum_im_mula(acum_re_mula'Length-1-NORMBIT downto acum_re_mula'Length-o_samplesQ'Length-NORMBIT);


	end if;
end process;


end qcomplex_norm;


