core_phaseerrors_mif_inst : core_phaseerrors_mif PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
