library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
library work;
use work.feedf_consts_pack.all;
use work.assert_pack.all;
use work.math_real.all;

USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

entity average_itertive_demod is
	generic(
		SIMULATION:integer:=1
	);
	port(
		clk : in STD_LOGIC;
		reset : in std_logic;
		after_pilot_start: in std_logic; --# �� ������ ���� ��� ������ i_ce
		i_ce : in std_logic;		
		i_samplesI: in std_logic_vector(15 downto 0);
		i_samplesQ: in std_logic_vector(15 downto 0);

		i_init_phaseI: in std_logic_vector(15 downto 0);
		i_init_phaseQ: in std_logic_vector(15 downto 0);

		o_samplesI: out std_logic_vector(15 downto 0);
		o_samplesQ: out std_logic_vector(15 downto 0);

		out_ce: out std_logic
		);
end average_itertive_demod;



architecture average_itertive_demod of average_itertive_demod is

function norming (val,x,y: std_logic_vector; rval:real) return std_logic_vector is
--# rval - future vector size
--# val - value that will be normalizate (or x or y)
--# x,y - input complex value
	variable abs_v:real;
	variable rett:std_logic_vector(val'Length-1 downto 0);
begin
	abs_v:=sqrt(real(conv_integer(signed(x)))*real(conv_integer(signed(x)))+real(conv_integer(signed(y)))*real(conv_integer(signed(y))) );
	if abs_v=0.0 then
		rett:=conv_std_logic_vector(0,val'Length);
	else
		rett:=conv_std_logic_vector(integer( rval*real(conv_integer(signed(val)))/abs_v ),val'Length);
	end if;
	return rett;
end norming;



function signed_abs (L: std_logic_vector) return std_logic_vector is
-- pragma label_applies_to abs
  
variable result : std_logic_vector(L'range) ;
--attribute IS_SIGNED of L:constant is TRUE ;
--attribute SYNTHESIS_RETURN of result:variable is "ABS" ;
begin
if (L(L'left) = '0' or L(L'left) = 'L') then
    result := L;
else
    result := 0 - signed(L);
end if;
    return result ;
end signed_abs;



function int_abs (L: integer) return integer is
	variable result : integer;
begin
	if (L>0) then
    	result := L;
	else
    	result := 0 - L;
	end if;
    return result ;
end int_abs;


constant NORMBIT:natural:=5;
constant NORMBITOUT:natural:=8;

type Tnorm_mem is array (0 to 1023) of std_logic_vector(7 downto 0);
constant norm_mem:Tnorm_mem:=  (
"11111111", 
"11111111", "10000000", "01010101", "01000000", "00110011", "00101011", "00100100", "00100000", "00011100", "00011010", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00010001", "00010010", "00010100", "00010101", 
"00010111", "00011010", "00011100", "00100000", "00100100", "00101011", "00110011", "01000000", "01010101", "10000000", "11111111", "11111111", "10110100", "01110010", "01010001", "00111110", "00110010", "00101010", "00100100", "00100000", 
"00011100", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00010001", "00010010", "00010100", "00010101", "00010111", "00011001", "00011100", "00100000", "00100100", "00101010", "00110010", "00111110", 
"01010001", "01110010", "10110100", "10000000", "01110010", "01011010", "01000111", "00111001", "00101111", "00101000", "00100011", "00011111", "00011100", "00011001", "00010111", "00010101", "00010011", "00010010", "00010001", "00010000", 
"00010001", "00010010", "00010011", "00010101", "00010111", "00011001", "00011100", "00011111", "00100011", "00101000", "00101111", "00111001", "01000111", "01011010", "01110010", "01010101", "01010001", "01000111", "00111100", "00110011", 
"00101100", "00100110", "00100001", "00011110", "00011011", "00011000", "00010110", "00010101", "00010011", "00010010", "00010001", "00010000", "00010001", "00010010", "00010011", "00010101", "00010110", "00011000", "00011011", "00011110", 
"00100001", "00100110", "00101100", "00110011", "00111100", "01000111", "01010001", "01000000", "00111110", "00111001", "00110011", "00101101", "00101000", "00100011", "00100000", "00011101", "00011010", "00011000", "00010110", "00010100", 
"00010011", "00010010", "00010000", "00001111", "00010000", "00010010", "00010011", "00010100", "00010110", "00011000", "00011010", "00011101", "00100000", "00100011", "00101000", "00101101", "00110011", "00111001", "00111110", "00110011", 
"00110010", "00101111", "00101100", "00101000", "00100100", "00100001", "00011110", "00011011", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", "00010000", "00010001", "00010010", "00010100", 
"00010101", "00010111", "00011001", "00011011", "00011110", "00100001", "00100100", "00101000", "00101100", "00101111", "00110010", "00101011", "00101010", "00101000", "00100110", "00100011", "00100001", "00011110", "00011100", "00011010", 
"00011000", "00010110", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010110", "00011000", "00011010", "00011100", "00011110", "00100001", "00100011", 
"00100110", "00101000", "00101010", "00100100", "00100100", "00100011", "00100001", "00100000", "00011110", "00011100", "00011010", "00011000", "00010110", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", "00001111", 
"00001111", "00010000", "00010001", "00010010", "00010100", "00010101", "00010110", "00011000", "00011010", "00011100", "00011110", "00100000", "00100001", "00100011", "00100100", "00100000", "00100000", "00011111", "00011110", "00011101", 
"00011011", "00011010", "00011000", "00010111", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010111", 
"00011000", "00011010", "00011011", "00011101", "00011110", "00011111", "00100000", "00011100", "00011100", "00011100", "00011011", "00011010", "00011001", "00011000", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", 
"00010000", "00001111", "00001111", "00001110", "00001111", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00011000", "00011001", "00011010", "00011011", "00011100", "00011100", "00011010", 
"00011001", "00011001", "00011000", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001110", "00001111", "00010000", "00010000", 
"00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011000", "00011001", "00011001", "00010111", "00010111", "00010111", "00010110", "00010110", "00010101", "00010100", "00010100", "00010011", 
"00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", "00010010", "00010011", "00010100", "00010100", "00010101", "00010110", 
"00010110", "00010111", "00010111", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", "00010011", "00010010", "00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001101", 
"00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", "00010010", "00010010", "00010011", "00010100", "00010100", "00010101", "00010101", "00010101", "00010100", "00010100", "00010011", "00010011", "00010011", 
"00010010", "00010010", "00010001", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", 
"00010001", "00010010", "00010010", "00010011", "00010011", "00010011", "00010100", "00010010", "00010010", "00010010", "00010010", "00010010", "00010001", "00010001", "00010000", "00010000", "00001111", "00001111", "00001110", "00001110", 
"00001101", "00001101", "00001100", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00001111", "00010000", "00010000", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010001", 
"00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001100", "00001100", "00001100", "00001101", "00001101", 
"00001110", "00001110", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001111", "00001110", 
"00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001100", "00001011", "00001100", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", 
"00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001100", 
"00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010010", 
"00010001", "00010001", "00010000", "00010000", "00001111", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00001111", "00010000", 
"00010000", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010100", "00010100", "00010011", "00010011", "00010011", "00010010", "00010010", "00010001", "00010001", "00010000", "00010000", "00001111", "00001110", 
"00001110", "00001101", "00001101", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", "00010001", "00010010", "00010010", "00010011", "00010011", "00010011", "00010100", "00010101", 
"00010101", "00010101", "00010101", "00010100", "00010100", "00010011", "00010010", "00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001101", "00001101", "00001110", "00001110", "00001111", 
"00010000", "00010000", "00010001", "00010010", "00010010", "00010011", "00010100", "00010100", "00010101", "00010101", "00010101", "00010111", "00010111", "00010111", "00010110", "00010110", "00010101", "00010100", "00010100", "00010011", 
"00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", "00001101", "00001110", "00001110", "00001111", "00010000", "00010000", "00010001", "00010010", "00010011", "00010100", "00010100", "00010101", "00010110", 
"00010110", "00010111", "00010111", "00011010", "00011001", "00011001", "00011000", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00010000", "00001111", "00001110", "00001110", 
"00001110", "00001111", "00010000", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011000", "00011001", "00011001", "00011100", "00011100", "00011100", "00011011", "00011010", 
"00011001", "00011000", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001111", "00001110", "00001111", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", 
"00010110", "00011000", "00011001", "00011010", "00011011", "00011100", "00011100", "00100000", "00100000", "00011111", "00011110", "00011101", "00011011", "00011010", "00011000", "00010111", "00010101", "00010100", "00010011", "00010010", 
"00010001", "00010000", "00001111", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010111", "00011000", "00011010", "00011011", "00011101", "00011110", "00011111", "00100000", "00100100", 
"00100100", "00100011", "00100001", "00100000", "00011110", "00011100", "00011010", "00011000", "00010110", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", "00001111", "00001111", "00010000", "00010001", "00010010", 
"00010100", "00010101", "00010110", "00011000", "00011010", "00011100", "00011110", "00100000", "00100001", "00100011", "00100100", "00101011", "00101010", "00101000", "00100110", "00100011", "00100001", "00011110", "00011100", "00011010", 
"00011000", "00010110", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010110", "00011000", "00011010", "00011100", "00011110", "00100001", "00100011", 
"00100110", "00101000", "00101010", "00110011", "00110010", "00101111", "00101100", "00101000", "00100100", "00100001", "00011110", "00011011", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", 
"00010000", "00010001", "00010010", "00010100", "00010101", "00010111", "00011001", "00011011", "00011110", "00100001", "00100100", "00101000", "00101100", "00101111", "00110010", "01000000", "00111110", "00111001", "00110011", "00101101", 
"00101000", "00100011", "00100000", "00011101", "00011010", "00011000", "00010110", "00010100", "00010011", "00010010", "00010000", "00001111", "00010000", "00010010", "00010011", "00010100", "00010110", "00011000", "00011010", "00011101", 
"00100000", "00100011", "00101000", "00101101", "00110011", "00111001", "00111110", "01010101", "01010001", "01000111", "00111100", "00110011", "00101100", "00100110", "00100001", "00011110", "00011011", "00011000", "00010110", "00010101", 
"00010011", "00010010", "00010001", "00010000", "00010001", "00010010", "00010011", "00010101", "00010110", "00011000", "00011011", "00011110", "00100001", "00100110", "00101100", "00110011", "00111100", "01000111", "01010001", "10000000", 
"01110010", "01011010", "01000111", "00111001", "00101111", "00101000", "00100011", "00011111", "00011100", "00011001", "00010111", "00010101", "00010011", "00010010", "00010001", "00010000", "00010001", "00010010", "00010011", "00010101", 
"00010111", "00011001", "00011100", "00011111", "00100011", "00101000", "00101111", "00111001", "01000111", "01011010", "01110010", "11111111", "10110100", "01110010", "01010001", "00111110", "00110010", "00101010", "00100100", "00100000", 
"00011100", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00010000", "00010001", "00010010", "00010100", "00010101", "00010111", "00011001", "00011100", "00100000", "00100100", "00101010", "00110010", "00111110", 
"01010001", "01110010", "10110100" );



constant BITSIZE:integer:=8;
constant SH:integer:=3;

signal mulval_a:std_logic_vector(NORMBITOUT-1 downto 0):=(others=>'0');
signal acum_re_1w,acum_im_1w,acum_re_new,acum_im_new,acum_re,acum_im,sample_rotI,sample_rotQ:std_logic_vector(15 downto 0);
signal acum_re_mula,acum_im_mula:std_logic_vector(15+NORMBITOUT+1 downto 0):=(others=>'0');
signal table_re,table_im,to_tab_re,to_tab_im:std_logic_vector(BITSIZE-1 downto 0);
signal table_reE,table_imE:std_logic_vector(15 downto 0);
signal ce_1w,ce_table,ce_acum,shift1,shift2:std_logic;
signal poval:std_logic_vector(NORMBIT*2-1 downto 0);
signal povval_x,povval_y:std_logic_vector(NORMBIT-1 downto 0);

begin

SIM01: if SIMULATION=1 generate
--	save_complexdata_i: entity work.save_complexdata
--		port map(
--		clk =>clk,
--		i_ce =>i_ce,
--		i_samplesI=>i_samplesI,
--		i_samplesQ=>i_samplesQ,
--
--		i_ce2 =>after_pilot_start,
--		i_samplesI2=>i_init_phaseI,
--		i_samplesQ2=>i_init_phaseQ
--		);
end generate;


table_reE<=table_re&EXT("0",16-BITSIZE);
table_imE<=table_im&EXT("0",16-BITSIZE);

complex_mult_q_i: entity work.complex_mult_q
	generic map(
		SHIFT_MUL=>1,
		CONJUGATION=>'1' --# ��������� �� ����������� �����, ���� '1' - �� ���������
	)
	port map(
		clk =>clk,
		i_ce =>i_ce,

		A_I=>i_samplesI,
		B_Q=>i_samplesQ,

		C_I=>acum_re,
		D_Q=>acum_im,

		o_I=>sample_rotI,
		o_Q=>sample_rotQ,
		out_ce=>open
		);

complex_mult_q_ii: entity work.complex_mult_qr
	generic map(
		SHIFT_MUL=>3, --# (����� ������� ��� 3)
		CONJUGATION=>'0' --# ��������� �� ����������� �����, ���� '1' - �� ���������
	)
	port map(
		clk =>clk,

		load =>after_pilot_start,

		init_I=>i_init_phaseI,
		init_Q=>i_init_phaseQ,

		i_ce =>ce_table,
		A_I=>acum_re_1w,       --# 6101+1i*1157  (�����)
		B_Q=>acum_im_1w,

		C_I=>table_reE,        --# 32256-1i*4352 (�����)
		D_Q=>table_imE,

		o_I=>acum_re_new, --# ��� ���������� ������������ ������ ���� 12318+1i*656
		o_Q=>acum_im_new,
		out_ce=>ce_acum
		);

shift1<='1' when unsigned(signed_abs(sample_rotI(sample_rotI'Length-1 downto 6)))>127 or unsigned(signed_abs(sample_rotQ(sample_rotQ'Length-1 downto 6)))>127  else '0';

--to_tab_re<=SXT(sample_rotI(sample_rotI'Length-1 downto 9),BITSIZE) when 
--	unsigned(signed_abs(sample_rotI(sample_rotI'Length-1 downto 6)))>127 or unsigned(signed_abs(sample_rotQ(sample_rotQ'Length-1 downto 6)))>127 
--	else sample_rotI(6+BITSIZE-1 downto 6);

--to_tab_im<=SXT(sample_rotQ(sample_rotQ'Length-1 downto 9),BITSIZE) when 
--	unsigned(signed_abs(sample_rotI(sample_rotI'Length-1 downto 6)))>127 or unsigned(signed_abs(sample_rotQ(sample_rotQ'Length-1 downto 6)))>127 
--	else sample_rotQ(6+BITSIZE-1 downto 6);

to_tab_re<=sample_rotI(5+BITSIZE-1 downto 5); --# !!!was
to_tab_im<=sample_rotQ(5+BITSIZE-1 downto 5);


--to_tab_re<=norming(sample_rotI(5+BITSIZE-1 downto 5),sample_rotI(5+BITSIZE-1 downto 5),sample_rotQ(5+BITSIZE-1 downto 5),8192.0);
--to_tab_im<=norming(sample_rotQ(5+BITSIZE-1 downto 5),sample_rotI(5+BITSIZE-1 downto 5),sample_rotQ(5+BITSIZE-1 downto 5),8192.0);


table_demod_i:entity work.table_demod
	generic map(
		BIT_IN=>BITSIZE,
		BIT_OUT=>BITSIZE
	)
	 port map(
		  clk =>clk,
		  i_ce=>ce_1w,
	      sample_in_re=>to_tab_re,
	      sample_in_im=>to_tab_im,
		  o_ce=>ce_table,
	      sample_out_re=>table_re,
	      sample_out_im=>table_im
		 );
		




povval_x<=acum_re_new(acum_re_new'Length-1-1 downto acum_re_new'Length-NORMBIT-1);  --# was
povval_y<=acum_im_new(acum_re_new'Length-1-1 downto acum_re_new'Length-NORMBIT-1);





poval<=acum_im_new(acum_re_new'Length-1-1 downto acum_re_new'Length-NORMBIT-1)&acum_re_new(acum_re_new'Length-1-1 downto acum_re_new'Length-NORMBIT-1);
mulval_a<=norm_mem(conv_integer(poval));

process(clk) is
variable v_acum_re_mula,v_acum_im_mula:std_logic_vector(acum_re_mula'Length-1 downto 0):=(others=>'0');

begin
	if rising_edge(clk) then
		ce_1w<=i_ce;
		out_ce<=i_ce;


o_samplesI<=norming(sample_rotI,sample_rotI,sample_rotQ,8192.0);
o_samplesQ<=norming(sample_rotQ,sample_rotI,sample_rotQ,8192.0);


--o_samplesI<=conv_std_logic_vector( integer(8192.0*real(conv_integer(signed(sample_rotI)))/sqrt(real(conv_integer(signed(sample_rotI)))*real(conv_integer(signed(sample_rotI)))+real(conv_integer(signed(sample_rotQ)))*real(conv_integer(signed(sample_rotQ))) )), o_samplesI'Length);
--o_samplesQ<=conv_std_logic_vector( integer(8192.0*real(conv_integer(signed(sample_rotQ)))/sqrt(real(conv_integer(signed(sample_rotI)))*real(conv_integer(signed(sample_rotI)))+real(conv_integer(signed(sample_rotQ)))*real(conv_integer(signed(sample_rotQ))) )), o_samplesI'Length);

--		o_samplesI<=sample_rotI;
--		o_samplesQ<=sample_rotQ;

--			acum_re_1w<=i_init_phaseI;
--			acum_im_1w<=i_init_phaseQ;

		if after_pilot_start='1' then
				acum_re_1w<=i_init_phaseI;
				acum_im_1w<=i_init_phaseQ;
		else
				acum_re_1w<=acum_re;
				acum_im_1w<=acum_im;
		end if;

--		if after_pilot_start='1' then
--			acum_re<=(others=>'0');--i_init_phaseI;
--			acum_im<=(others=>'0');--i_init_phaseQ;
--		else        --# reset
--			if ce_acum='1' then



				v_acum_re_mula:=signed(acum_re_new)*signed('0'&mulval_a);
				v_acum_im_mula:=signed(acum_im_new)*signed('0'&mulval_a);

				acum_re_mula<=signed(acum_re_new)*signed('0'&mulval_a);
				acum_im_mula<=signed(acum_im_new)*signed('0'&mulval_a);

--# was
--				acum_re<=v_acum_re_mula(acum_re_mula'Length-1-(NORMBIT-1) downto acum_re_mula'Length-acum_re'Length-(NORMBIT-1));
--				acum_im<=v_acum_im_mula(acum_re_mula'Length-1-(NORMBIT-1) downto acum_re_mula'Length-acum_re'Length-(NORMBIT-1));

				acum_re<=norming(acum_re_new,acum_re_new,acum_im_new,8192.0);
				acum_im<=norming(acum_im_new,acum_re_new,acum_im_new,8192.0);


--				acum_re<=conv_std_logic_vector( integer(8192.0*real(conv_integer(signed(acum_re_new)))/sqrt(real(conv_integer(signed(acum_re_new)))*real(conv_integer(signed(acum_re_new)))+real(conv_integer(signed(acum_im_new)))*real(conv_integer(signed(acum_im_new))) )), acum_re'Length);
--				acum_im<=conv_std_logic_vector( integer(8192.0*real(conv_integer(signed(acum_im_new)))/sqrt(real(conv_integer(signed(acum_re_new)))*real(conv_integer(signed(acum_re_new)))+real(conv_integer(signed(acum_im_new)))*real(conv_integer(signed(acum_im_new))) )), acum_re'Length);



--			end if; --# i_ce
--		end if;     --# reset
	end if;
end process;



end average_itertive_demod;



