sqrt32to16_altera_inst : sqrt32to16_altera PORT MAP (
		aclr	 => aclr_sig,
		clk	 => clk_sig,
		ena	 => ena_sig,
		radical	 => radical_sig,
		q	 => q_sig,
		remainder	 => remainder_sig
	);
