module table_phaseerrors
(
input wire clk,
input wire[8:0] input_angles,
input wire[8:0] phase_acum_mod,

output reg [8:0] phi_error,
output reg [9:0] val_engle
);
wire [15:0] test_pos;
reg [18:0] ram [65535:0];


initial begin
ram[0] = {9'd0,10'd0};
ram[1] = {9'd3,10'd3};
ram[2] = {9'd6,10'd6};
ram[3] = {9'd9,10'd9};
ram[4] = {9'd12,10'd12};
ram[5] = {9'd15,10'd15};
ram[6] = {9'd18,10'd18};
ram[7] = {9'd21,10'd21};
ram[8] = {9'd25,10'd25};
ram[9] = {9'd28,10'd28};
ram[10] = {9'd31,10'd31};
ram[11] = {9'd34,10'd34};
ram[12] = {9'd37,10'd37};
ram[13] = {9'd40,10'd40};
ram[14] = {9'd43,10'd43};
ram[15] = {9'd47,10'd47};
ram[16] = {9'd50,10'd50};
ram[17] = {9'd53,10'd53};
ram[18] = {9'd56,10'd56};
ram[19] = {9'd59,10'd59};
ram[20] = {9'd62,10'd62};
ram[21] = {9'd65,10'd65};
ram[22] = {9'd69,10'd69};
ram[23] = {9'd72,10'd72};
ram[24] = {9'd75,10'd75};
ram[25] = {9'd78,10'd78};
ram[26] = {9'd81,10'd81};
ram[27] = {9'd84,10'd84};
ram[28] = {9'd87,10'd87};
ram[29] = {9'd91,10'd91};
ram[30] = {9'd94,10'd94};
ram[31] = {9'd97,10'd97};
ram[32] = {-9'd100,10'd100};
ram[33] = {-9'd97,10'd103};
ram[34] = {-9'd94,10'd106};
ram[35] = {-9'd91,10'd109};
ram[36] = {-9'd88,10'd113};
ram[37] = {-9'd85,10'd116};
ram[38] = {-9'd81,10'd119};
ram[39] = {-9'd78,10'd122};
ram[40] = {-9'd75,10'd125};
ram[41] = {-9'd72,10'd128};
ram[42] = {-9'd69,10'd131};
ram[43] = {-9'd66,10'd135};
ram[44] = {-9'd63,10'd138};
ram[45] = {-9'd59,10'd141};
ram[46] = {-9'd56,10'd144};
ram[47] = {-9'd53,10'd147};
ram[48] = {-9'd50,10'd150};
ram[49] = {-9'd47,10'd153};
ram[50] = {-9'd44,10'd157};
ram[51] = {-9'd41,10'd160};
ram[52] = {-9'd37,10'd163};
ram[53] = {-9'd34,10'd166};
ram[54] = {-9'd31,10'd169};
ram[55] = {-9'd28,10'd172};
ram[56] = {-9'd25,10'd175};
ram[57] = {-9'd22,10'd179};
ram[58] = {-9'd19,10'd182};
ram[59] = {-9'd15,10'd185};
ram[60] = {-9'd12,10'd188};
ram[61] = {-9'd9,10'd191};
ram[62] = {-9'd6,10'd194};
ram[63] = {-9'd3,10'd197};
ram[64] = {9'd0,10'd201};
ram[65] = {9'd3,10'd204};
ram[66] = {9'd7,10'd207};
ram[67] = {9'd10,10'd210};
ram[68] = {9'd13,10'd213};
ram[69] = {9'd16,10'd216};
ram[70] = {9'd19,10'd219};
ram[71] = {9'd22,10'd223};
ram[72] = {9'd25,10'd226};
ram[73] = {9'd29,10'd229};
ram[74] = {9'd32,10'd232};
ram[75] = {9'd35,10'd235};
ram[76] = {9'd38,10'd238};
ram[77] = {9'd41,10'd241};
ram[78] = {9'd44,10'd245};
ram[79] = {9'd47,10'd248};
ram[80] = {9'd51,10'd251};
ram[81] = {9'd54,10'd254};
ram[82] = {9'd57,10'd257};
ram[83] = {9'd60,10'd260};
ram[84] = {9'd63,10'd263};
ram[85] = {9'd66,10'd267};
ram[86] = {9'd69,10'd270};
ram[87] = {9'd73,10'd273};
ram[88] = {9'd76,10'd276};
ram[89] = {9'd79,10'd279};
ram[90] = {9'd82,10'd282};
ram[91] = {9'd85,10'd285};
ram[92] = {9'd88,10'd289};
ram[93] = {9'd91,10'd292};
ram[94] = {9'd95,10'd295};
ram[95] = {9'd98,10'd298};
ram[96] = {-9'd99,10'd301};
ram[97] = {-9'd96,10'd304};
ram[98] = {-9'd93,10'd307};
ram[99] = {-9'd90,10'd311};
ram[100] = {-9'd87,10'd314};
ram[101] = {-9'd84,10'd317};
ram[102] = {-9'd81,10'd320};
ram[103] = {-9'd77,10'd323};
ram[104] = {-9'd74,10'd326};
ram[105] = {-9'd71,10'd329};
ram[106] = {-9'd68,10'd333};
ram[107] = {-9'd65,10'd336};
ram[108] = {-9'd62,10'd339};
ram[109] = {-9'd59,10'd342};
ram[110] = {-9'd55,10'd345};
ram[111] = {-9'd52,10'd348};
ram[112] = {-9'd49,10'd351};
ram[113] = {-9'd46,10'd354};
ram[114] = {-9'd43,10'd358};
ram[115] = {-9'd40,10'd361};
ram[116] = {-9'd37,10'd364};
ram[117] = {-9'd33,10'd367};
ram[118] = {-9'd30,10'd370};
ram[119] = {-9'd27,10'd373};
ram[120] = {-9'd24,10'd376};
ram[121] = {-9'd21,10'd380};
ram[122] = {-9'd18,10'd383};
ram[123] = {-9'd15,10'd386};
ram[124] = {-9'd11,10'd389};
ram[125] = {-9'd8,10'd392};
ram[126] = {-9'd5,10'd395};
ram[127] = {-9'd2,10'd398};
ram[128] = {-9'd2,10'd398};
ram[129] = {9'd1,-10'd399};
ram[130] = {9'd4,-10'd396};
ram[131] = {9'd7,-10'd393};
ram[132] = {9'd10,-10'd390};
ram[133] = {9'd14,-10'd387};
ram[134] = {9'd17,-10'd384};
ram[135] = {9'd20,-10'd381};
ram[136] = {9'd23,-10'd377};
ram[137] = {9'd26,-10'd374};
ram[138] = {9'd29,-10'd371};
ram[139] = {9'd32,-10'd368};
ram[140] = {9'd36,-10'd365};
ram[141] = {9'd39,-10'd362};
ram[142] = {9'd42,-10'd359};
ram[143] = {9'd45,-10'd355};
ram[144] = {9'd48,-10'd352};
ram[145] = {9'd51,-10'd349};
ram[146] = {9'd54,-10'd346};
ram[147] = {9'd58,-10'd343};
ram[148] = {9'd61,-10'd340};
ram[149] = {9'd64,-10'd337};
ram[150] = {9'd67,-10'd334};
ram[151] = {9'd70,-10'd330};
ram[152] = {9'd73,-10'd327};
ram[153] = {9'd76,-10'd324};
ram[154] = {9'd80,-10'd321};
ram[155] = {9'd83,-10'd318};
ram[156] = {9'd86,-10'd315};
ram[157] = {9'd89,-10'd312};
ram[158] = {9'd92,-10'd308};
ram[159] = {9'd95,-10'd305};
ram[160] = {9'd98,-10'd302};
ram[161] = {-9'd99,-10'd299};
ram[162] = {-9'd96,-10'd296};
ram[163] = {-9'd92,-10'd293};
ram[164] = {-9'd89,-10'd290};
ram[165] = {-9'd86,-10'd286};
ram[166] = {-9'd83,-10'd283};
ram[167] = {-9'd80,-10'd280};
ram[168] = {-9'd77,-10'd277};
ram[169] = {-9'd74,-10'd274};
ram[170] = {-9'd70,-10'd271};
ram[171] = {-9'd67,-10'd268};
ram[172] = {-9'd64,-10'd264};
ram[173] = {-9'd61,-10'd261};
ram[174] = {-9'd58,-10'd258};
ram[175] = {-9'd55,-10'd255};
ram[176] = {-9'd52,-10'd252};
ram[177] = {-9'd48,-10'd249};
ram[178] = {-9'd45,-10'd246};
ram[179] = {-9'd42,-10'd242};
ram[180] = {-9'd39,-10'd239};
ram[181] = {-9'd36,-10'd236};
ram[182] = {-9'd33,-10'd233};
ram[183] = {-9'd30,-10'd230};
ram[184] = {-9'd26,-10'd227};
ram[185] = {-9'd23,-10'd224};
ram[186] = {-9'd20,-10'd220};
ram[187] = {-9'd17,-10'd217};
ram[188] = {-9'd14,-10'd214};
ram[189] = {-9'd11,-10'd211};
ram[190] = {-9'd8,-10'd208};
ram[191] = {-9'd4,-10'd205};
ram[192] = {-9'd1,-10'd202};
ram[193] = {9'd2,-10'd198};
ram[194] = {9'd5,-10'd195};
ram[195] = {9'd8,-10'd192};
ram[196] = {9'd11,-10'd189};
ram[197] = {9'd14,-10'd186};
ram[198] = {9'd18,-10'd183};
ram[199] = {9'd21,-10'd180};
ram[200] = {9'd24,-10'd176};
ram[201] = {9'd27,-10'd173};
ram[202] = {9'd30,-10'd170};
ram[203] = {9'd33,-10'd167};
ram[204] = {9'd36,-10'd164};
ram[205] = {9'd40,-10'd161};
ram[206] = {9'd43,-10'd158};
ram[207] = {9'd46,-10'd154};
ram[208] = {9'd49,-10'd151};
ram[209] = {9'd52,-10'd148};
ram[210] = {9'd55,-10'd145};
ram[211] = {9'd58,-10'd142};
ram[212] = {9'd62,-10'd139};
ram[213] = {9'd65,-10'd136};
ram[214] = {9'd68,-10'd132};
ram[215] = {9'd71,-10'd129};
ram[216] = {9'd74,-10'd126};
ram[217] = {9'd77,-10'd123};
ram[218] = {9'd80,-10'd120};
ram[219] = {9'd84,-10'd117};
ram[220] = {9'd87,-10'd114};
ram[221] = {9'd90,-10'd110};
ram[222] = {9'd93,-10'd107};
ram[223] = {9'd96,-10'd104};
ram[224] = {9'd99,-10'd101};
ram[225] = {-9'd98,-10'd98};
ram[226] = {-9'd95,-10'd95};
ram[227] = {-9'd92,-10'd92};
ram[228] = {-9'd88,-10'd88};
ram[229] = {-9'd85,-10'd85};
ram[230] = {-9'd82,-10'd82};
ram[231] = {-9'd79,-10'd79};
ram[232] = {-9'd76,-10'd76};
ram[233] = {-9'd73,-10'd73};
ram[234] = {-9'd70,-10'd70};
ram[235] = {-9'd66,-10'd66};
ram[236] = {-9'd63,-10'd63};
ram[237] = {-9'd60,-10'd60};
ram[238] = {-9'd57,-10'd57};
ram[239] = {-9'd54,-10'd54};
ram[240] = {-9'd51,-10'd51};
ram[241] = {-9'd48,-10'd48};
ram[242] = {-9'd44,-10'd44};
ram[243] = {-9'd41,-10'd41};
ram[244] = {-9'd38,-10'd38};
ram[245] = {-9'd35,-10'd35};
ram[246] = {-9'd32,-10'd32};
ram[247] = {-9'd29,-10'd29};
ram[248] = {-9'd26,-10'd26};
ram[249] = {-9'd22,-10'd22};
ram[250] = {-9'd19,-10'd19};
ram[251] = {-9'd16,-10'd16};
ram[252] = {-9'd13,-10'd13};
ram[253] = {-9'd10,-10'd10};
ram[254] = {-9'd7,-10'd7};
ram[255] = {-9'd4,-10'd4};
ram[256] = {-9'd4,-10'd4};
ram[257] = {9'd0,10'd0};
ram[258] = {9'd3,10'd3};
ram[259] = {9'd6,10'd6};
ram[260] = {9'd9,10'd9};
ram[261] = {9'd12,10'd12};
ram[262] = {9'd15,10'd15};
ram[263] = {9'd18,10'd18};
ram[264] = {9'd21,10'd21};
ram[265] = {9'd25,10'd25};
ram[266] = {9'd28,10'd28};
ram[267] = {9'd31,10'd31};
ram[268] = {9'd34,10'd34};
ram[269] = {9'd37,10'd37};
ram[270] = {9'd40,10'd40};
ram[271] = {9'd43,10'd43};
ram[272] = {9'd47,10'd47};
ram[273] = {9'd50,10'd50};
ram[274] = {9'd53,10'd53};
ram[275] = {9'd56,10'd56};
ram[276] = {9'd59,10'd59};
ram[277] = {9'd62,10'd62};
ram[278] = {9'd65,10'd65};
ram[279] = {9'd69,10'd69};
ram[280] = {9'd72,10'd72};
ram[281] = {9'd75,10'd75};
ram[282] = {9'd78,10'd78};
ram[283] = {9'd81,10'd81};
ram[284] = {9'd84,10'd84};
ram[285] = {9'd87,10'd87};
ram[286] = {9'd91,10'd91};
ram[287] = {9'd94,10'd94};
ram[288] = {9'd97,10'd97};
ram[289] = {-9'd100,10'd100};
ram[290] = {-9'd97,10'd103};
ram[291] = {-9'd94,10'd106};
ram[292] = {-9'd91,10'd109};
ram[293] = {-9'd88,10'd113};
ram[294] = {-9'd85,10'd116};
ram[295] = {-9'd81,10'd119};
ram[296] = {-9'd78,10'd122};
ram[297] = {-9'd75,10'd125};
ram[298] = {-9'd72,10'd128};
ram[299] = {-9'd69,10'd131};
ram[300] = {-9'd66,10'd135};
ram[301] = {-9'd63,10'd138};
ram[302] = {-9'd59,10'd141};
ram[303] = {-9'd56,10'd144};
ram[304] = {-9'd53,10'd147};
ram[305] = {-9'd50,10'd150};
ram[306] = {-9'd47,10'd153};
ram[307] = {-9'd44,10'd157};
ram[308] = {-9'd41,10'd160};
ram[309] = {-9'd37,10'd163};
ram[310] = {-9'd34,10'd166};
ram[311] = {-9'd31,10'd169};
ram[312] = {-9'd28,10'd172};
ram[313] = {-9'd25,10'd175};
ram[314] = {-9'd22,10'd179};
ram[315] = {-9'd19,10'd182};
ram[316] = {-9'd15,10'd185};
ram[317] = {-9'd12,10'd188};
ram[318] = {-9'd9,10'd191};
ram[319] = {-9'd6,10'd194};
ram[320] = {-9'd3,10'd197};
ram[321] = {9'd0,10'd201};
ram[322] = {9'd3,10'd204};
ram[323] = {9'd7,10'd207};
ram[324] = {9'd10,10'd210};
ram[325] = {9'd13,10'd213};
ram[326] = {9'd16,10'd216};
ram[327] = {9'd19,10'd219};
ram[328] = {9'd22,10'd223};
ram[329] = {9'd25,10'd226};
ram[330] = {9'd29,10'd229};
ram[331] = {9'd32,10'd232};
ram[332] = {9'd35,10'd235};
ram[333] = {9'd38,10'd238};
ram[334] = {9'd41,10'd241};
ram[335] = {9'd44,10'd245};
ram[336] = {9'd47,10'd248};
ram[337] = {9'd51,10'd251};
ram[338] = {9'd54,10'd254};
ram[339] = {9'd57,10'd257};
ram[340] = {9'd60,10'd260};
ram[341] = {9'd63,10'd263};
ram[342] = {9'd66,10'd267};
ram[343] = {9'd69,10'd270};
ram[344] = {9'd73,10'd273};
ram[345] = {9'd76,10'd276};
ram[346] = {9'd79,10'd279};
ram[347] = {9'd82,10'd282};
ram[348] = {9'd85,10'd285};
ram[349] = {9'd88,10'd289};
ram[350] = {9'd91,10'd292};
ram[351] = {9'd95,10'd295};
ram[352] = {9'd98,10'd298};
ram[353] = {-9'd99,10'd301};
ram[354] = {-9'd96,10'd304};
ram[355] = {-9'd93,10'd307};
ram[356] = {-9'd90,10'd311};
ram[357] = {-9'd87,10'd314};
ram[358] = {-9'd84,10'd317};
ram[359] = {-9'd81,10'd320};
ram[360] = {-9'd77,10'd323};
ram[361] = {-9'd74,10'd326};
ram[362] = {-9'd71,10'd329};
ram[363] = {-9'd68,10'd333};
ram[364] = {-9'd65,10'd336};
ram[365] = {-9'd62,10'd339};
ram[366] = {-9'd59,10'd342};
ram[367] = {-9'd55,10'd345};
ram[368] = {-9'd52,10'd348};
ram[369] = {-9'd49,10'd351};
ram[370] = {-9'd46,10'd354};
ram[371] = {-9'd43,10'd358};
ram[372] = {-9'd40,10'd361};
ram[373] = {-9'd37,10'd364};
ram[374] = {-9'd33,10'd367};
ram[375] = {-9'd30,10'd370};
ram[376] = {-9'd27,10'd373};
ram[377] = {-9'd24,10'd376};
ram[378] = {-9'd21,10'd380};
ram[379] = {-9'd18,10'd383};
ram[380] = {-9'd15,10'd386};
ram[381] = {-9'd11,10'd389};
ram[382] = {-9'd8,10'd392};
ram[383] = {-9'd5,10'd395};
ram[384] = {-9'd5,10'd395};
ram[385] = {-9'd2,10'd398};
ram[386] = {9'd1,-10'd399};
ram[387] = {9'd4,-10'd396};
ram[388] = {9'd7,-10'd393};
ram[389] = {9'd10,-10'd390};
ram[390] = {9'd14,-10'd387};
ram[391] = {9'd17,-10'd384};
ram[392] = {9'd20,-10'd381};
ram[393] = {9'd23,-10'd377};
ram[394] = {9'd26,-10'd374};
ram[395] = {9'd29,-10'd371};
ram[396] = {9'd32,-10'd368};
ram[397] = {9'd36,-10'd365};
ram[398] = {9'd39,-10'd362};
ram[399] = {9'd42,-10'd359};
ram[400] = {9'd45,-10'd355};
ram[401] = {9'd48,-10'd352};
ram[402] = {9'd51,-10'd349};
ram[403] = {9'd54,-10'd346};
ram[404] = {9'd58,-10'd343};
ram[405] = {9'd61,-10'd340};
ram[406] = {9'd64,-10'd337};
ram[407] = {9'd67,-10'd334};
ram[408] = {9'd70,-10'd330};
ram[409] = {9'd73,-10'd327};
ram[410] = {9'd76,-10'd324};
ram[411] = {9'd80,-10'd321};
ram[412] = {9'd83,-10'd318};
ram[413] = {9'd86,-10'd315};
ram[414] = {9'd89,-10'd312};
ram[415] = {9'd92,-10'd308};
ram[416] = {9'd95,-10'd305};
ram[417] = {9'd98,-10'd302};
ram[418] = {-9'd99,-10'd299};
ram[419] = {-9'd96,-10'd296};
ram[420] = {-9'd92,-10'd293};
ram[421] = {-9'd89,-10'd290};
ram[422] = {-9'd86,-10'd286};
ram[423] = {-9'd83,-10'd283};
ram[424] = {-9'd80,-10'd280};
ram[425] = {-9'd77,-10'd277};
ram[426] = {-9'd74,-10'd274};
ram[427] = {-9'd70,-10'd271};
ram[428] = {-9'd67,-10'd268};
ram[429] = {-9'd64,-10'd264};
ram[430] = {-9'd61,-10'd261};
ram[431] = {-9'd58,-10'd258};
ram[432] = {-9'd55,-10'd255};
ram[433] = {-9'd52,-10'd252};
ram[434] = {-9'd48,-10'd249};
ram[435] = {-9'd45,-10'd246};
ram[436] = {-9'd42,-10'd242};
ram[437] = {-9'd39,-10'd239};
ram[438] = {-9'd36,-10'd236};
ram[439] = {-9'd33,-10'd233};
ram[440] = {-9'd30,-10'd230};
ram[441] = {-9'd26,-10'd227};
ram[442] = {-9'd23,-10'd224};
ram[443] = {-9'd20,-10'd220};
ram[444] = {-9'd17,-10'd217};
ram[445] = {-9'd14,-10'd214};
ram[446] = {-9'd11,-10'd211};
ram[447] = {-9'd8,-10'd208};
ram[448] = {-9'd4,-10'd205};
ram[449] = {-9'd1,-10'd202};
ram[450] = {9'd2,-10'd198};
ram[451] = {9'd5,-10'd195};
ram[452] = {9'd8,-10'd192};
ram[453] = {9'd11,-10'd189};
ram[454] = {9'd14,-10'd186};
ram[455] = {9'd18,-10'd183};
ram[456] = {9'd21,-10'd180};
ram[457] = {9'd24,-10'd176};
ram[458] = {9'd27,-10'd173};
ram[459] = {9'd30,-10'd170};
ram[460] = {9'd33,-10'd167};
ram[461] = {9'd36,-10'd164};
ram[462] = {9'd40,-10'd161};
ram[463] = {9'd43,-10'd158};
ram[464] = {9'd46,-10'd154};
ram[465] = {9'd49,-10'd151};
ram[466] = {9'd52,-10'd148};
ram[467] = {9'd55,-10'd145};
ram[468] = {9'd58,-10'd142};
ram[469] = {9'd62,-10'd139};
ram[470] = {9'd65,-10'd136};
ram[471] = {9'd68,-10'd132};
ram[472] = {9'd71,-10'd129};
ram[473] = {9'd74,-10'd126};
ram[474] = {9'd77,-10'd123};
ram[475] = {9'd80,-10'd120};
ram[476] = {9'd84,-10'd117};
ram[477] = {9'd87,-10'd114};
ram[478] = {9'd90,-10'd110};
ram[479] = {9'd93,-10'd107};
ram[480] = {9'd96,-10'd104};
ram[481] = {9'd99,-10'd101};
ram[482] = {-9'd98,-10'd98};
ram[483] = {-9'd95,-10'd95};
ram[484] = {-9'd92,-10'd92};
ram[485] = {-9'd88,-10'd88};
ram[486] = {-9'd85,-10'd85};
ram[487] = {-9'd82,-10'd82};
ram[488] = {-9'd79,-10'd79};
ram[489] = {-9'd76,-10'd76};
ram[490] = {-9'd73,-10'd73};
ram[491] = {-9'd70,-10'd70};
ram[492] = {-9'd66,-10'd66};
ram[493] = {-9'd63,-10'd63};
ram[494] = {-9'd60,-10'd60};
ram[495] = {-9'd57,-10'd57};
ram[496] = {-9'd54,-10'd54};
ram[497] = {-9'd51,-10'd51};
ram[498] = {-9'd48,-10'd48};
ram[499] = {-9'd44,-10'd44};
ram[500] = {-9'd41,-10'd41};
ram[501] = {-9'd38,-10'd38};
ram[502] = {-9'd35,-10'd35};
ram[503] = {-9'd32,-10'd32};
ram[504] = {-9'd29,-10'd29};
ram[505] = {-9'd26,-10'd26};
ram[506] = {-9'd22,-10'd22};
ram[507] = {-9'd19,-10'd19};
ram[508] = {-9'd16,-10'd16};
ram[509] = {-9'd13,-10'd13};
ram[510] = {-9'd10,-10'd10};
ram[511] = {-9'd7,-10'd7};
ram[512] = {-9'd7,-10'd7};
ram[513] = {-9'd4,-10'd4};
ram[514] = {9'd0,10'd0};
ram[515] = {9'd3,10'd3};
ram[516] = {9'd6,10'd6};
ram[517] = {9'd9,10'd9};
ram[518] = {9'd12,10'd12};
ram[519] = {9'd15,10'd15};
ram[520] = {9'd18,10'd18};
ram[521] = {9'd21,10'd21};
ram[522] = {9'd25,10'd25};
ram[523] = {9'd28,10'd28};
ram[524] = {9'd31,10'd31};
ram[525] = {9'd34,10'd34};
ram[526] = {9'd37,10'd37};
ram[527] = {9'd40,10'd40};
ram[528] = {9'd43,10'd43};
ram[529] = {9'd47,10'd47};
ram[530] = {9'd50,10'd50};
ram[531] = {9'd53,10'd53};
ram[532] = {9'd56,10'd56};
ram[533] = {9'd59,10'd59};
ram[534] = {9'd62,10'd62};
ram[535] = {9'd65,10'd65};
ram[536] = {9'd69,10'd69};
ram[537] = {9'd72,10'd72};
ram[538] = {9'd75,10'd75};
ram[539] = {9'd78,10'd78};
ram[540] = {9'd81,10'd81};
ram[541] = {9'd84,10'd84};
ram[542] = {9'd87,10'd87};
ram[543] = {9'd91,10'd91};
ram[544] = {9'd94,10'd94};
ram[545] = {9'd97,10'd97};
ram[546] = {-9'd100,10'd100};
ram[547] = {-9'd97,10'd103};
ram[548] = {-9'd94,10'd106};
ram[549] = {-9'd91,10'd109};
ram[550] = {-9'd88,10'd113};
ram[551] = {-9'd85,10'd116};
ram[552] = {-9'd81,10'd119};
ram[553] = {-9'd78,10'd122};
ram[554] = {-9'd75,10'd125};
ram[555] = {-9'd72,10'd128};
ram[556] = {-9'd69,10'd131};
ram[557] = {-9'd66,10'd135};
ram[558] = {-9'd63,10'd138};
ram[559] = {-9'd59,10'd141};
ram[560] = {-9'd56,10'd144};
ram[561] = {-9'd53,10'd147};
ram[562] = {-9'd50,10'd150};
ram[563] = {-9'd47,10'd153};
ram[564] = {-9'd44,10'd157};
ram[565] = {-9'd41,10'd160};
ram[566] = {-9'd37,10'd163};
ram[567] = {-9'd34,10'd166};
ram[568] = {-9'd31,10'd169};
ram[569] = {-9'd28,10'd172};
ram[570] = {-9'd25,10'd175};
ram[571] = {-9'd22,10'd179};
ram[572] = {-9'd19,10'd182};
ram[573] = {-9'd15,10'd185};
ram[574] = {-9'd12,10'd188};
ram[575] = {-9'd9,10'd191};
ram[576] = {-9'd6,10'd194};
ram[577] = {-9'd3,10'd197};
ram[578] = {9'd0,10'd201};
ram[579] = {9'd3,10'd204};
ram[580] = {9'd7,10'd207};
ram[581] = {9'd10,10'd210};
ram[582] = {9'd13,10'd213};
ram[583] = {9'd16,10'd216};
ram[584] = {9'd19,10'd219};
ram[585] = {9'd22,10'd223};
ram[586] = {9'd25,10'd226};
ram[587] = {9'd29,10'd229};
ram[588] = {9'd32,10'd232};
ram[589] = {9'd35,10'd235};
ram[590] = {9'd38,10'd238};
ram[591] = {9'd41,10'd241};
ram[592] = {9'd44,10'd245};
ram[593] = {9'd47,10'd248};
ram[594] = {9'd51,10'd251};
ram[595] = {9'd54,10'd254};
ram[596] = {9'd57,10'd257};
ram[597] = {9'd60,10'd260};
ram[598] = {9'd63,10'd263};
ram[599] = {9'd66,10'd267};
ram[600] = {9'd69,10'd270};
ram[601] = {9'd73,10'd273};
ram[602] = {9'd76,10'd276};
ram[603] = {9'd79,10'd279};
ram[604] = {9'd82,10'd282};
ram[605] = {9'd85,10'd285};
ram[606] = {9'd88,10'd289};
ram[607] = {9'd91,10'd292};
ram[608] = {9'd95,10'd295};
ram[609] = {9'd98,10'd298};
ram[610] = {-9'd99,10'd301};
ram[611] = {-9'd96,10'd304};
ram[612] = {-9'd93,10'd307};
ram[613] = {-9'd90,10'd311};
ram[614] = {-9'd87,10'd314};
ram[615] = {-9'd84,10'd317};
ram[616] = {-9'd81,10'd320};
ram[617] = {-9'd77,10'd323};
ram[618] = {-9'd74,10'd326};
ram[619] = {-9'd71,10'd329};
ram[620] = {-9'd68,10'd333};
ram[621] = {-9'd65,10'd336};
ram[622] = {-9'd62,10'd339};
ram[623] = {-9'd59,10'd342};
ram[624] = {-9'd55,10'd345};
ram[625] = {-9'd52,10'd348};
ram[626] = {-9'd49,10'd351};
ram[627] = {-9'd46,10'd354};
ram[628] = {-9'd43,10'd358};
ram[629] = {-9'd40,10'd361};
ram[630] = {-9'd37,10'd364};
ram[631] = {-9'd33,10'd367};
ram[632] = {-9'd30,10'd370};
ram[633] = {-9'd27,10'd373};
ram[634] = {-9'd24,10'd376};
ram[635] = {-9'd21,10'd380};
ram[636] = {-9'd18,10'd383};
ram[637] = {-9'd15,10'd386};
ram[638] = {-9'd11,10'd389};
ram[639] = {-9'd8,10'd392};
ram[640] = {-9'd8,10'd392};
ram[641] = {-9'd5,10'd395};
ram[642] = {-9'd2,10'd398};
ram[643] = {9'd1,-10'd399};
ram[644] = {9'd4,-10'd396};
ram[645] = {9'd7,-10'd393};
ram[646] = {9'd10,-10'd390};
ram[647] = {9'd14,-10'd387};
ram[648] = {9'd17,-10'd384};
ram[649] = {9'd20,-10'd381};
ram[650] = {9'd23,-10'd377};
ram[651] = {9'd26,-10'd374};
ram[652] = {9'd29,-10'd371};
ram[653] = {9'd32,-10'd368};
ram[654] = {9'd36,-10'd365};
ram[655] = {9'd39,-10'd362};
ram[656] = {9'd42,-10'd359};
ram[657] = {9'd45,-10'd355};
ram[658] = {9'd48,-10'd352};
ram[659] = {9'd51,-10'd349};
ram[660] = {9'd54,-10'd346};
ram[661] = {9'd58,-10'd343};
ram[662] = {9'd61,-10'd340};
ram[663] = {9'd64,-10'd337};
ram[664] = {9'd67,-10'd334};
ram[665] = {9'd70,-10'd330};
ram[666] = {9'd73,-10'd327};
ram[667] = {9'd76,-10'd324};
ram[668] = {9'd80,-10'd321};
ram[669] = {9'd83,-10'd318};
ram[670] = {9'd86,-10'd315};
ram[671] = {9'd89,-10'd312};
ram[672] = {9'd92,-10'd308};
ram[673] = {9'd95,-10'd305};
ram[674] = {9'd98,-10'd302};
ram[675] = {-9'd99,-10'd299};
ram[676] = {-9'd96,-10'd296};
ram[677] = {-9'd92,-10'd293};
ram[678] = {-9'd89,-10'd290};
ram[679] = {-9'd86,-10'd286};
ram[680] = {-9'd83,-10'd283};
ram[681] = {-9'd80,-10'd280};
ram[682] = {-9'd77,-10'd277};
ram[683] = {-9'd74,-10'd274};
ram[684] = {-9'd70,-10'd271};
ram[685] = {-9'd67,-10'd268};
ram[686] = {-9'd64,-10'd264};
ram[687] = {-9'd61,-10'd261};
ram[688] = {-9'd58,-10'd258};
ram[689] = {-9'd55,-10'd255};
ram[690] = {-9'd52,-10'd252};
ram[691] = {-9'd48,-10'd249};
ram[692] = {-9'd45,-10'd246};
ram[693] = {-9'd42,-10'd242};
ram[694] = {-9'd39,-10'd239};
ram[695] = {-9'd36,-10'd236};
ram[696] = {-9'd33,-10'd233};
ram[697] = {-9'd30,-10'd230};
ram[698] = {-9'd26,-10'd227};
ram[699] = {-9'd23,-10'd224};
ram[700] = {-9'd20,-10'd220};
ram[701] = {-9'd17,-10'd217};
ram[702] = {-9'd14,-10'd214};
ram[703] = {-9'd11,-10'd211};
ram[704] = {-9'd8,-10'd208};
ram[705] = {-9'd4,-10'd205};
ram[706] = {-9'd1,-10'd202};
ram[707] = {9'd2,-10'd198};
ram[708] = {9'd5,-10'd195};
ram[709] = {9'd8,-10'd192};
ram[710] = {9'd11,-10'd189};
ram[711] = {9'd14,-10'd186};
ram[712] = {9'd18,-10'd183};
ram[713] = {9'd21,-10'd180};
ram[714] = {9'd24,-10'd176};
ram[715] = {9'd27,-10'd173};
ram[716] = {9'd30,-10'd170};
ram[717] = {9'd33,-10'd167};
ram[718] = {9'd36,-10'd164};
ram[719] = {9'd40,-10'd161};
ram[720] = {9'd43,-10'd158};
ram[721] = {9'd46,-10'd154};
ram[722] = {9'd49,-10'd151};
ram[723] = {9'd52,-10'd148};
ram[724] = {9'd55,-10'd145};
ram[725] = {9'd58,-10'd142};
ram[726] = {9'd62,-10'd139};
ram[727] = {9'd65,-10'd136};
ram[728] = {9'd68,-10'd132};
ram[729] = {9'd71,-10'd129};
ram[730] = {9'd74,-10'd126};
ram[731] = {9'd77,-10'd123};
ram[732] = {9'd80,-10'd120};
ram[733] = {9'd84,-10'd117};
ram[734] = {9'd87,-10'd114};
ram[735] = {9'd90,-10'd110};
ram[736] = {9'd93,-10'd107};
ram[737] = {9'd96,-10'd104};
ram[738] = {9'd99,-10'd101};
ram[739] = {-9'd98,-10'd98};
ram[740] = {-9'd95,-10'd95};
ram[741] = {-9'd92,-10'd92};
ram[742] = {-9'd88,-10'd88};
ram[743] = {-9'd85,-10'd85};
ram[744] = {-9'd82,-10'd82};
ram[745] = {-9'd79,-10'd79};
ram[746] = {-9'd76,-10'd76};
ram[747] = {-9'd73,-10'd73};
ram[748] = {-9'd70,-10'd70};
ram[749] = {-9'd66,-10'd66};
ram[750] = {-9'd63,-10'd63};
ram[751] = {-9'd60,-10'd60};
ram[752] = {-9'd57,-10'd57};
ram[753] = {-9'd54,-10'd54};
ram[754] = {-9'd51,-10'd51};
ram[755] = {-9'd48,-10'd48};
ram[756] = {-9'd44,-10'd44};
ram[757] = {-9'd41,-10'd41};
ram[758] = {-9'd38,-10'd38};
ram[759] = {-9'd35,-10'd35};
ram[760] = {-9'd32,-10'd32};
ram[761] = {-9'd29,-10'd29};
ram[762] = {-9'd26,-10'd26};
ram[763] = {-9'd22,-10'd22};
ram[764] = {-9'd19,-10'd19};
ram[765] = {-9'd16,-10'd16};
ram[766] = {-9'd13,-10'd13};
ram[767] = {-9'd10,-10'd10};
ram[768] = {-9'd10,-10'd10};
ram[769] = {-9'd7,-10'd7};
ram[770] = {-9'd4,-10'd4};
ram[771] = {9'd0,10'd0};
ram[772] = {9'd3,10'd3};
ram[773] = {9'd6,10'd6};
ram[774] = {9'd9,10'd9};
ram[775] = {9'd12,10'd12};
ram[776] = {9'd15,10'd15};
ram[777] = {9'd18,10'd18};
ram[778] = {9'd21,10'd21};
ram[779] = {9'd25,10'd25};
ram[780] = {9'd28,10'd28};
ram[781] = {9'd31,10'd31};
ram[782] = {9'd34,10'd34};
ram[783] = {9'd37,10'd37};
ram[784] = {9'd40,10'd40};
ram[785] = {9'd43,10'd43};
ram[786] = {9'd47,10'd47};
ram[787] = {9'd50,10'd50};
ram[788] = {9'd53,10'd53};
ram[789] = {9'd56,10'd56};
ram[790] = {9'd59,10'd59};
ram[791] = {9'd62,10'd62};
ram[792] = {9'd65,10'd65};
ram[793] = {9'd69,10'd69};
ram[794] = {9'd72,10'd72};
ram[795] = {9'd75,10'd75};
ram[796] = {9'd78,10'd78};
ram[797] = {9'd81,10'd81};
ram[798] = {9'd84,10'd84};
ram[799] = {9'd87,10'd87};
ram[800] = {9'd91,10'd91};
ram[801] = {9'd94,10'd94};
ram[802] = {9'd97,10'd97};
ram[803] = {-9'd100,10'd100};
ram[804] = {-9'd97,10'd103};
ram[805] = {-9'd94,10'd106};
ram[806] = {-9'd91,10'd109};
ram[807] = {-9'd88,10'd113};
ram[808] = {-9'd85,10'd116};
ram[809] = {-9'd81,10'd119};
ram[810] = {-9'd78,10'd122};
ram[811] = {-9'd75,10'd125};
ram[812] = {-9'd72,10'd128};
ram[813] = {-9'd69,10'd131};
ram[814] = {-9'd66,10'd135};
ram[815] = {-9'd63,10'd138};
ram[816] = {-9'd59,10'd141};
ram[817] = {-9'd56,10'd144};
ram[818] = {-9'd53,10'd147};
ram[819] = {-9'd50,10'd150};
ram[820] = {-9'd47,10'd153};
ram[821] = {-9'd44,10'd157};
ram[822] = {-9'd41,10'd160};
ram[823] = {-9'd37,10'd163};
ram[824] = {-9'd34,10'd166};
ram[825] = {-9'd31,10'd169};
ram[826] = {-9'd28,10'd172};
ram[827] = {-9'd25,10'd175};
ram[828] = {-9'd22,10'd179};
ram[829] = {-9'd19,10'd182};
ram[830] = {-9'd15,10'd185};
ram[831] = {-9'd12,10'd188};
ram[832] = {-9'd9,10'd191};
ram[833] = {-9'd6,10'd194};
ram[834] = {-9'd3,10'd197};
ram[835] = {9'd0,10'd201};
ram[836] = {9'd3,10'd204};
ram[837] = {9'd7,10'd207};
ram[838] = {9'd10,10'd210};
ram[839] = {9'd13,10'd213};
ram[840] = {9'd16,10'd216};
ram[841] = {9'd19,10'd219};
ram[842] = {9'd22,10'd223};
ram[843] = {9'd25,10'd226};
ram[844] = {9'd29,10'd229};
ram[845] = {9'd32,10'd232};
ram[846] = {9'd35,10'd235};
ram[847] = {9'd38,10'd238};
ram[848] = {9'd41,10'd241};
ram[849] = {9'd44,10'd245};
ram[850] = {9'd47,10'd248};
ram[851] = {9'd51,10'd251};
ram[852] = {9'd54,10'd254};
ram[853] = {9'd57,10'd257};
ram[854] = {9'd60,10'd260};
ram[855] = {9'd63,10'd263};
ram[856] = {9'd66,10'd267};
ram[857] = {9'd69,10'd270};
ram[858] = {9'd73,10'd273};
ram[859] = {9'd76,10'd276};
ram[860] = {9'd79,10'd279};
ram[861] = {9'd82,10'd282};
ram[862] = {9'd85,10'd285};
ram[863] = {9'd88,10'd289};
ram[864] = {9'd91,10'd292};
ram[865] = {9'd95,10'd295};
ram[866] = {9'd98,10'd298};
ram[867] = {-9'd99,10'd301};
ram[868] = {-9'd96,10'd304};
ram[869] = {-9'd93,10'd307};
ram[870] = {-9'd90,10'd311};
ram[871] = {-9'd87,10'd314};
ram[872] = {-9'd84,10'd317};
ram[873] = {-9'd81,10'd320};
ram[874] = {-9'd77,10'd323};
ram[875] = {-9'd74,10'd326};
ram[876] = {-9'd71,10'd329};
ram[877] = {-9'd68,10'd333};
ram[878] = {-9'd65,10'd336};
ram[879] = {-9'd62,10'd339};
ram[880] = {-9'd59,10'd342};
ram[881] = {-9'd55,10'd345};
ram[882] = {-9'd52,10'd348};
ram[883] = {-9'd49,10'd351};
ram[884] = {-9'd46,10'd354};
ram[885] = {-9'd43,10'd358};
ram[886] = {-9'd40,10'd361};
ram[887] = {-9'd37,10'd364};
ram[888] = {-9'd33,10'd367};
ram[889] = {-9'd30,10'd370};
ram[890] = {-9'd27,10'd373};
ram[891] = {-9'd24,10'd376};
ram[892] = {-9'd21,10'd380};
ram[893] = {-9'd18,10'd383};
ram[894] = {-9'd15,10'd386};
ram[895] = {-9'd11,10'd389};
ram[896] = {-9'd11,10'd389};
ram[897] = {-9'd8,10'd392};
ram[898] = {-9'd5,10'd395};
ram[899] = {-9'd2,10'd398};
ram[900] = {9'd1,-10'd399};
ram[901] = {9'd4,-10'd396};
ram[902] = {9'd7,-10'd393};
ram[903] = {9'd10,-10'd390};
ram[904] = {9'd14,-10'd387};
ram[905] = {9'd17,-10'd384};
ram[906] = {9'd20,-10'd381};
ram[907] = {9'd23,-10'd377};
ram[908] = {9'd26,-10'd374};
ram[909] = {9'd29,-10'd371};
ram[910] = {9'd32,-10'd368};
ram[911] = {9'd36,-10'd365};
ram[912] = {9'd39,-10'd362};
ram[913] = {9'd42,-10'd359};
ram[914] = {9'd45,-10'd355};
ram[915] = {9'd48,-10'd352};
ram[916] = {9'd51,-10'd349};
ram[917] = {9'd54,-10'd346};
ram[918] = {9'd58,-10'd343};
ram[919] = {9'd61,-10'd340};
ram[920] = {9'd64,-10'd337};
ram[921] = {9'd67,-10'd334};
ram[922] = {9'd70,-10'd330};
ram[923] = {9'd73,-10'd327};
ram[924] = {9'd76,-10'd324};
ram[925] = {9'd80,-10'd321};
ram[926] = {9'd83,-10'd318};
ram[927] = {9'd86,-10'd315};
ram[928] = {9'd89,-10'd312};
ram[929] = {9'd92,-10'd308};
ram[930] = {9'd95,-10'd305};
ram[931] = {9'd98,-10'd302};
ram[932] = {-9'd99,-10'd299};
ram[933] = {-9'd96,-10'd296};
ram[934] = {-9'd92,-10'd293};
ram[935] = {-9'd89,-10'd290};
ram[936] = {-9'd86,-10'd286};
ram[937] = {-9'd83,-10'd283};
ram[938] = {-9'd80,-10'd280};
ram[939] = {-9'd77,-10'd277};
ram[940] = {-9'd74,-10'd274};
ram[941] = {-9'd70,-10'd271};
ram[942] = {-9'd67,-10'd268};
ram[943] = {-9'd64,-10'd264};
ram[944] = {-9'd61,-10'd261};
ram[945] = {-9'd58,-10'd258};
ram[946] = {-9'd55,-10'd255};
ram[947] = {-9'd52,-10'd252};
ram[948] = {-9'd48,-10'd249};
ram[949] = {-9'd45,-10'd246};
ram[950] = {-9'd42,-10'd242};
ram[951] = {-9'd39,-10'd239};
ram[952] = {-9'd36,-10'd236};
ram[953] = {-9'd33,-10'd233};
ram[954] = {-9'd30,-10'd230};
ram[955] = {-9'd26,-10'd227};
ram[956] = {-9'd23,-10'd224};
ram[957] = {-9'd20,-10'd220};
ram[958] = {-9'd17,-10'd217};
ram[959] = {-9'd14,-10'd214};
ram[960] = {-9'd11,-10'd211};
ram[961] = {-9'd8,-10'd208};
ram[962] = {-9'd4,-10'd205};
ram[963] = {-9'd1,-10'd202};
ram[964] = {9'd2,-10'd198};
ram[965] = {9'd5,-10'd195};
ram[966] = {9'd8,-10'd192};
ram[967] = {9'd11,-10'd189};
ram[968] = {9'd14,-10'd186};
ram[969] = {9'd18,-10'd183};
ram[970] = {9'd21,-10'd180};
ram[971] = {9'd24,-10'd176};
ram[972] = {9'd27,-10'd173};
ram[973] = {9'd30,-10'd170};
ram[974] = {9'd33,-10'd167};
ram[975] = {9'd36,-10'd164};
ram[976] = {9'd40,-10'd161};
ram[977] = {9'd43,-10'd158};
ram[978] = {9'd46,-10'd154};
ram[979] = {9'd49,-10'd151};
ram[980] = {9'd52,-10'd148};
ram[981] = {9'd55,-10'd145};
ram[982] = {9'd58,-10'd142};
ram[983] = {9'd62,-10'd139};
ram[984] = {9'd65,-10'd136};
ram[985] = {9'd68,-10'd132};
ram[986] = {9'd71,-10'd129};
ram[987] = {9'd74,-10'd126};
ram[988] = {9'd77,-10'd123};
ram[989] = {9'd80,-10'd120};
ram[990] = {9'd84,-10'd117};
ram[991] = {9'd87,-10'd114};
ram[992] = {9'd90,-10'd110};
ram[993] = {9'd93,-10'd107};
ram[994] = {9'd96,-10'd104};
ram[995] = {9'd99,-10'd101};
ram[996] = {-9'd98,-10'd98};
ram[997] = {-9'd95,-10'd95};
ram[998] = {-9'd92,-10'd92};
ram[999] = {-9'd88,-10'd88};
ram[1000] = {-9'd85,-10'd85};
ram[1001] = {-9'd82,-10'd82};
ram[1002] = {-9'd79,-10'd79};
ram[1003] = {-9'd76,-10'd76};
ram[1004] = {-9'd73,-10'd73};
ram[1005] = {-9'd70,-10'd70};
ram[1006] = {-9'd66,-10'd66};
ram[1007] = {-9'd63,-10'd63};
ram[1008] = {-9'd60,-10'd60};
ram[1009] = {-9'd57,-10'd57};
ram[1010] = {-9'd54,-10'd54};
ram[1011] = {-9'd51,-10'd51};
ram[1012] = {-9'd48,-10'd48};
ram[1013] = {-9'd44,-10'd44};
ram[1014] = {-9'd41,-10'd41};
ram[1015] = {-9'd38,-10'd38};
ram[1016] = {-9'd35,-10'd35};
ram[1017] = {-9'd32,-10'd32};
ram[1018] = {-9'd29,-10'd29};
ram[1019] = {-9'd26,-10'd26};
ram[1020] = {-9'd22,-10'd22};
ram[1021] = {-9'd19,-10'd19};
ram[1022] = {-9'd16,-10'd16};
ram[1023] = {-9'd13,-10'd13};
ram[1024] = {-9'd13,-10'd13};
ram[1025] = {-9'd10,-10'd10};
ram[1026] = {-9'd7,-10'd7};
ram[1027] = {-9'd4,-10'd4};
ram[1028] = {9'd0,10'd0};
ram[1029] = {9'd3,10'd3};
ram[1030] = {9'd6,10'd6};
ram[1031] = {9'd9,10'd9};
ram[1032] = {9'd12,10'd12};
ram[1033] = {9'd15,10'd15};
ram[1034] = {9'd18,10'd18};
ram[1035] = {9'd21,10'd21};
ram[1036] = {9'd25,10'd25};
ram[1037] = {9'd28,10'd28};
ram[1038] = {9'd31,10'd31};
ram[1039] = {9'd34,10'd34};
ram[1040] = {9'd37,10'd37};
ram[1041] = {9'd40,10'd40};
ram[1042] = {9'd43,10'd43};
ram[1043] = {9'd47,10'd47};
ram[1044] = {9'd50,10'd50};
ram[1045] = {9'd53,10'd53};
ram[1046] = {9'd56,10'd56};
ram[1047] = {9'd59,10'd59};
ram[1048] = {9'd62,10'd62};
ram[1049] = {9'd65,10'd65};
ram[1050] = {9'd69,10'd69};
ram[1051] = {9'd72,10'd72};
ram[1052] = {9'd75,10'd75};
ram[1053] = {9'd78,10'd78};
ram[1054] = {9'd81,10'd81};
ram[1055] = {9'd84,10'd84};
ram[1056] = {9'd87,10'd87};
ram[1057] = {9'd91,10'd91};
ram[1058] = {9'd94,10'd94};
ram[1059] = {9'd97,10'd97};
ram[1060] = {-9'd100,10'd100};
ram[1061] = {-9'd97,10'd103};
ram[1062] = {-9'd94,10'd106};
ram[1063] = {-9'd91,10'd109};
ram[1064] = {-9'd88,10'd113};
ram[1065] = {-9'd85,10'd116};
ram[1066] = {-9'd81,10'd119};
ram[1067] = {-9'd78,10'd122};
ram[1068] = {-9'd75,10'd125};
ram[1069] = {-9'd72,10'd128};
ram[1070] = {-9'd69,10'd131};
ram[1071] = {-9'd66,10'd135};
ram[1072] = {-9'd63,10'd138};
ram[1073] = {-9'd59,10'd141};
ram[1074] = {-9'd56,10'd144};
ram[1075] = {-9'd53,10'd147};
ram[1076] = {-9'd50,10'd150};
ram[1077] = {-9'd47,10'd153};
ram[1078] = {-9'd44,10'd157};
ram[1079] = {-9'd41,10'd160};
ram[1080] = {-9'd37,10'd163};
ram[1081] = {-9'd34,10'd166};
ram[1082] = {-9'd31,10'd169};
ram[1083] = {-9'd28,10'd172};
ram[1084] = {-9'd25,10'd175};
ram[1085] = {-9'd22,10'd179};
ram[1086] = {-9'd19,10'd182};
ram[1087] = {-9'd15,10'd185};
ram[1088] = {-9'd12,10'd188};
ram[1089] = {-9'd9,10'd191};
ram[1090] = {-9'd6,10'd194};
ram[1091] = {-9'd3,10'd197};
ram[1092] = {9'd0,10'd201};
ram[1093] = {9'd3,10'd204};
ram[1094] = {9'd7,10'd207};
ram[1095] = {9'd10,10'd210};
ram[1096] = {9'd13,10'd213};
ram[1097] = {9'd16,10'd216};
ram[1098] = {9'd19,10'd219};
ram[1099] = {9'd22,10'd223};
ram[1100] = {9'd25,10'd226};
ram[1101] = {9'd29,10'd229};
ram[1102] = {9'd32,10'd232};
ram[1103] = {9'd35,10'd235};
ram[1104] = {9'd38,10'd238};
ram[1105] = {9'd41,10'd241};
ram[1106] = {9'd44,10'd245};
ram[1107] = {9'd47,10'd248};
ram[1108] = {9'd51,10'd251};
ram[1109] = {9'd54,10'd254};
ram[1110] = {9'd57,10'd257};
ram[1111] = {9'd60,10'd260};
ram[1112] = {9'd63,10'd263};
ram[1113] = {9'd66,10'd267};
ram[1114] = {9'd69,10'd270};
ram[1115] = {9'd73,10'd273};
ram[1116] = {9'd76,10'd276};
ram[1117] = {9'd79,10'd279};
ram[1118] = {9'd82,10'd282};
ram[1119] = {9'd85,10'd285};
ram[1120] = {9'd88,10'd289};
ram[1121] = {9'd91,10'd292};
ram[1122] = {9'd95,10'd295};
ram[1123] = {9'd98,10'd298};
ram[1124] = {-9'd99,10'd301};
ram[1125] = {-9'd96,10'd304};
ram[1126] = {-9'd93,10'd307};
ram[1127] = {-9'd90,10'd311};
ram[1128] = {-9'd87,10'd314};
ram[1129] = {-9'd84,10'd317};
ram[1130] = {-9'd81,10'd320};
ram[1131] = {-9'd77,10'd323};
ram[1132] = {-9'd74,10'd326};
ram[1133] = {-9'd71,10'd329};
ram[1134] = {-9'd68,10'd333};
ram[1135] = {-9'd65,10'd336};
ram[1136] = {-9'd62,10'd339};
ram[1137] = {-9'd59,10'd342};
ram[1138] = {-9'd55,10'd345};
ram[1139] = {-9'd52,10'd348};
ram[1140] = {-9'd49,10'd351};
ram[1141] = {-9'd46,10'd354};
ram[1142] = {-9'd43,10'd358};
ram[1143] = {-9'd40,10'd361};
ram[1144] = {-9'd37,10'd364};
ram[1145] = {-9'd33,10'd367};
ram[1146] = {-9'd30,10'd370};
ram[1147] = {-9'd27,10'd373};
ram[1148] = {-9'd24,10'd376};
ram[1149] = {-9'd21,10'd380};
ram[1150] = {-9'd18,10'd383};
ram[1151] = {-9'd15,10'd386};
ram[1152] = {-9'd15,10'd386};
ram[1153] = {-9'd11,10'd389};
ram[1154] = {-9'd8,10'd392};
ram[1155] = {-9'd5,10'd395};
ram[1156] = {-9'd2,10'd398};
ram[1157] = {9'd1,-10'd399};
ram[1158] = {9'd4,-10'd396};
ram[1159] = {9'd7,-10'd393};
ram[1160] = {9'd10,-10'd390};
ram[1161] = {9'd14,-10'd387};
ram[1162] = {9'd17,-10'd384};
ram[1163] = {9'd20,-10'd381};
ram[1164] = {9'd23,-10'd377};
ram[1165] = {9'd26,-10'd374};
ram[1166] = {9'd29,-10'd371};
ram[1167] = {9'd32,-10'd368};
ram[1168] = {9'd36,-10'd365};
ram[1169] = {9'd39,-10'd362};
ram[1170] = {9'd42,-10'd359};
ram[1171] = {9'd45,-10'd355};
ram[1172] = {9'd48,-10'd352};
ram[1173] = {9'd51,-10'd349};
ram[1174] = {9'd54,-10'd346};
ram[1175] = {9'd58,-10'd343};
ram[1176] = {9'd61,-10'd340};
ram[1177] = {9'd64,-10'd337};
ram[1178] = {9'd67,-10'd334};
ram[1179] = {9'd70,-10'd330};
ram[1180] = {9'd73,-10'd327};
ram[1181] = {9'd76,-10'd324};
ram[1182] = {9'd80,-10'd321};
ram[1183] = {9'd83,-10'd318};
ram[1184] = {9'd86,-10'd315};
ram[1185] = {9'd89,-10'd312};
ram[1186] = {9'd92,-10'd308};
ram[1187] = {9'd95,-10'd305};
ram[1188] = {9'd98,-10'd302};
ram[1189] = {-9'd99,-10'd299};
ram[1190] = {-9'd96,-10'd296};
ram[1191] = {-9'd92,-10'd293};
ram[1192] = {-9'd89,-10'd290};
ram[1193] = {-9'd86,-10'd286};
ram[1194] = {-9'd83,-10'd283};
ram[1195] = {-9'd80,-10'd280};
ram[1196] = {-9'd77,-10'd277};
ram[1197] = {-9'd74,-10'd274};
ram[1198] = {-9'd70,-10'd271};
ram[1199] = {-9'd67,-10'd268};
ram[1200] = {-9'd64,-10'd264};
ram[1201] = {-9'd61,-10'd261};
ram[1202] = {-9'd58,-10'd258};
ram[1203] = {-9'd55,-10'd255};
ram[1204] = {-9'd52,-10'd252};
ram[1205] = {-9'd48,-10'd249};
ram[1206] = {-9'd45,-10'd246};
ram[1207] = {-9'd42,-10'd242};
ram[1208] = {-9'd39,-10'd239};
ram[1209] = {-9'd36,-10'd236};
ram[1210] = {-9'd33,-10'd233};
ram[1211] = {-9'd30,-10'd230};
ram[1212] = {-9'd26,-10'd227};
ram[1213] = {-9'd23,-10'd224};
ram[1214] = {-9'd20,-10'd220};
ram[1215] = {-9'd17,-10'd217};
ram[1216] = {-9'd14,-10'd214};
ram[1217] = {-9'd11,-10'd211};
ram[1218] = {-9'd8,-10'd208};
ram[1219] = {-9'd4,-10'd205};
ram[1220] = {-9'd1,-10'd202};
ram[1221] = {9'd2,-10'd198};
ram[1222] = {9'd5,-10'd195};
ram[1223] = {9'd8,-10'd192};
ram[1224] = {9'd11,-10'd189};
ram[1225] = {9'd14,-10'd186};
ram[1226] = {9'd18,-10'd183};
ram[1227] = {9'd21,-10'd180};
ram[1228] = {9'd24,-10'd176};
ram[1229] = {9'd27,-10'd173};
ram[1230] = {9'd30,-10'd170};
ram[1231] = {9'd33,-10'd167};
ram[1232] = {9'd36,-10'd164};
ram[1233] = {9'd40,-10'd161};
ram[1234] = {9'd43,-10'd158};
ram[1235] = {9'd46,-10'd154};
ram[1236] = {9'd49,-10'd151};
ram[1237] = {9'd52,-10'd148};
ram[1238] = {9'd55,-10'd145};
ram[1239] = {9'd58,-10'd142};
ram[1240] = {9'd62,-10'd139};
ram[1241] = {9'd65,-10'd136};
ram[1242] = {9'd68,-10'd132};
ram[1243] = {9'd71,-10'd129};
ram[1244] = {9'd74,-10'd126};
ram[1245] = {9'd77,-10'd123};
ram[1246] = {9'd80,-10'd120};
ram[1247] = {9'd84,-10'd117};
ram[1248] = {9'd87,-10'd114};
ram[1249] = {9'd90,-10'd110};
ram[1250] = {9'd93,-10'd107};
ram[1251] = {9'd96,-10'd104};
ram[1252] = {9'd99,-10'd101};
ram[1253] = {-9'd98,-10'd98};
ram[1254] = {-9'd95,-10'd95};
ram[1255] = {-9'd92,-10'd92};
ram[1256] = {-9'd88,-10'd88};
ram[1257] = {-9'd85,-10'd85};
ram[1258] = {-9'd82,-10'd82};
ram[1259] = {-9'd79,-10'd79};
ram[1260] = {-9'd76,-10'd76};
ram[1261] = {-9'd73,-10'd73};
ram[1262] = {-9'd70,-10'd70};
ram[1263] = {-9'd66,-10'd66};
ram[1264] = {-9'd63,-10'd63};
ram[1265] = {-9'd60,-10'd60};
ram[1266] = {-9'd57,-10'd57};
ram[1267] = {-9'd54,-10'd54};
ram[1268] = {-9'd51,-10'd51};
ram[1269] = {-9'd48,-10'd48};
ram[1270] = {-9'd44,-10'd44};
ram[1271] = {-9'd41,-10'd41};
ram[1272] = {-9'd38,-10'd38};
ram[1273] = {-9'd35,-10'd35};
ram[1274] = {-9'd32,-10'd32};
ram[1275] = {-9'd29,-10'd29};
ram[1276] = {-9'd26,-10'd26};
ram[1277] = {-9'd22,-10'd22};
ram[1278] = {-9'd19,-10'd19};
ram[1279] = {-9'd16,-10'd16};
ram[1280] = {-9'd16,-10'd16};
ram[1281] = {-9'd13,-10'd13};
ram[1282] = {-9'd10,-10'd10};
ram[1283] = {-9'd7,-10'd7};
ram[1284] = {-9'd4,-10'd4};
ram[1285] = {9'd0,10'd0};
ram[1286] = {9'd3,10'd3};
ram[1287] = {9'd6,10'd6};
ram[1288] = {9'd9,10'd9};
ram[1289] = {9'd12,10'd12};
ram[1290] = {9'd15,10'd15};
ram[1291] = {9'd18,10'd18};
ram[1292] = {9'd21,10'd21};
ram[1293] = {9'd25,10'd25};
ram[1294] = {9'd28,10'd28};
ram[1295] = {9'd31,10'd31};
ram[1296] = {9'd34,10'd34};
ram[1297] = {9'd37,10'd37};
ram[1298] = {9'd40,10'd40};
ram[1299] = {9'd43,10'd43};
ram[1300] = {9'd47,10'd47};
ram[1301] = {9'd50,10'd50};
ram[1302] = {9'd53,10'd53};
ram[1303] = {9'd56,10'd56};
ram[1304] = {9'd59,10'd59};
ram[1305] = {9'd62,10'd62};
ram[1306] = {9'd65,10'd65};
ram[1307] = {9'd69,10'd69};
ram[1308] = {9'd72,10'd72};
ram[1309] = {9'd75,10'd75};
ram[1310] = {9'd78,10'd78};
ram[1311] = {9'd81,10'd81};
ram[1312] = {9'd84,10'd84};
ram[1313] = {9'd87,10'd87};
ram[1314] = {9'd91,10'd91};
ram[1315] = {9'd94,10'd94};
ram[1316] = {9'd97,10'd97};
ram[1317] = {-9'd100,10'd100};
ram[1318] = {-9'd97,10'd103};
ram[1319] = {-9'd94,10'd106};
ram[1320] = {-9'd91,10'd109};
ram[1321] = {-9'd88,10'd113};
ram[1322] = {-9'd85,10'd116};
ram[1323] = {-9'd81,10'd119};
ram[1324] = {-9'd78,10'd122};
ram[1325] = {-9'd75,10'd125};
ram[1326] = {-9'd72,10'd128};
ram[1327] = {-9'd69,10'd131};
ram[1328] = {-9'd66,10'd135};
ram[1329] = {-9'd63,10'd138};
ram[1330] = {-9'd59,10'd141};
ram[1331] = {-9'd56,10'd144};
ram[1332] = {-9'd53,10'd147};
ram[1333] = {-9'd50,10'd150};
ram[1334] = {-9'd47,10'd153};
ram[1335] = {-9'd44,10'd157};
ram[1336] = {-9'd41,10'd160};
ram[1337] = {-9'd37,10'd163};
ram[1338] = {-9'd34,10'd166};
ram[1339] = {-9'd31,10'd169};
ram[1340] = {-9'd28,10'd172};
ram[1341] = {-9'd25,10'd175};
ram[1342] = {-9'd22,10'd179};
ram[1343] = {-9'd19,10'd182};
ram[1344] = {-9'd15,10'd185};
ram[1345] = {-9'd12,10'd188};
ram[1346] = {-9'd9,10'd191};
ram[1347] = {-9'd6,10'd194};
ram[1348] = {-9'd3,10'd197};
ram[1349] = {9'd0,10'd201};
ram[1350] = {9'd3,10'd204};
ram[1351] = {9'd7,10'd207};
ram[1352] = {9'd10,10'd210};
ram[1353] = {9'd13,10'd213};
ram[1354] = {9'd16,10'd216};
ram[1355] = {9'd19,10'd219};
ram[1356] = {9'd22,10'd223};
ram[1357] = {9'd25,10'd226};
ram[1358] = {9'd29,10'd229};
ram[1359] = {9'd32,10'd232};
ram[1360] = {9'd35,10'd235};
ram[1361] = {9'd38,10'd238};
ram[1362] = {9'd41,10'd241};
ram[1363] = {9'd44,10'd245};
ram[1364] = {9'd47,10'd248};
ram[1365] = {9'd51,10'd251};
ram[1366] = {9'd54,10'd254};
ram[1367] = {9'd57,10'd257};
ram[1368] = {9'd60,10'd260};
ram[1369] = {9'd63,10'd263};
ram[1370] = {9'd66,10'd267};
ram[1371] = {9'd69,10'd270};
ram[1372] = {9'd73,10'd273};
ram[1373] = {9'd76,10'd276};
ram[1374] = {9'd79,10'd279};
ram[1375] = {9'd82,10'd282};
ram[1376] = {9'd85,10'd285};
ram[1377] = {9'd88,10'd289};
ram[1378] = {9'd91,10'd292};
ram[1379] = {9'd95,10'd295};
ram[1380] = {9'd98,10'd298};
ram[1381] = {-9'd99,10'd301};
ram[1382] = {-9'd96,10'd304};
ram[1383] = {-9'd93,10'd307};
ram[1384] = {-9'd90,10'd311};
ram[1385] = {-9'd87,10'd314};
ram[1386] = {-9'd84,10'd317};
ram[1387] = {-9'd81,10'd320};
ram[1388] = {-9'd77,10'd323};
ram[1389] = {-9'd74,10'd326};
ram[1390] = {-9'd71,10'd329};
ram[1391] = {-9'd68,10'd333};
ram[1392] = {-9'd65,10'd336};
ram[1393] = {-9'd62,10'd339};
ram[1394] = {-9'd59,10'd342};
ram[1395] = {-9'd55,10'd345};
ram[1396] = {-9'd52,10'd348};
ram[1397] = {-9'd49,10'd351};
ram[1398] = {-9'd46,10'd354};
ram[1399] = {-9'd43,10'd358};
ram[1400] = {-9'd40,10'd361};
ram[1401] = {-9'd37,10'd364};
ram[1402] = {-9'd33,10'd367};
ram[1403] = {-9'd30,10'd370};
ram[1404] = {-9'd27,10'd373};
ram[1405] = {-9'd24,10'd376};
ram[1406] = {-9'd21,10'd380};
ram[1407] = {-9'd18,10'd383};
ram[1408] = {-9'd18,10'd383};
ram[1409] = {-9'd15,10'd386};
ram[1410] = {-9'd11,10'd389};
ram[1411] = {-9'd8,10'd392};
ram[1412] = {-9'd5,10'd395};
ram[1413] = {-9'd2,10'd398};
ram[1414] = {9'd1,-10'd399};
ram[1415] = {9'd4,-10'd396};
ram[1416] = {9'd7,-10'd393};
ram[1417] = {9'd10,-10'd390};
ram[1418] = {9'd14,-10'd387};
ram[1419] = {9'd17,-10'd384};
ram[1420] = {9'd20,-10'd381};
ram[1421] = {9'd23,-10'd377};
ram[1422] = {9'd26,-10'd374};
ram[1423] = {9'd29,-10'd371};
ram[1424] = {9'd32,-10'd368};
ram[1425] = {9'd36,-10'd365};
ram[1426] = {9'd39,-10'd362};
ram[1427] = {9'd42,-10'd359};
ram[1428] = {9'd45,-10'd355};
ram[1429] = {9'd48,-10'd352};
ram[1430] = {9'd51,-10'd349};
ram[1431] = {9'd54,-10'd346};
ram[1432] = {9'd58,-10'd343};
ram[1433] = {9'd61,-10'd340};
ram[1434] = {9'd64,-10'd337};
ram[1435] = {9'd67,-10'd334};
ram[1436] = {9'd70,-10'd330};
ram[1437] = {9'd73,-10'd327};
ram[1438] = {9'd76,-10'd324};
ram[1439] = {9'd80,-10'd321};
ram[1440] = {9'd83,-10'd318};
ram[1441] = {9'd86,-10'd315};
ram[1442] = {9'd89,-10'd312};
ram[1443] = {9'd92,-10'd308};
ram[1444] = {9'd95,-10'd305};
ram[1445] = {9'd98,-10'd302};
ram[1446] = {-9'd99,-10'd299};
ram[1447] = {-9'd96,-10'd296};
ram[1448] = {-9'd92,-10'd293};
ram[1449] = {-9'd89,-10'd290};
ram[1450] = {-9'd86,-10'd286};
ram[1451] = {-9'd83,-10'd283};
ram[1452] = {-9'd80,-10'd280};
ram[1453] = {-9'd77,-10'd277};
ram[1454] = {-9'd74,-10'd274};
ram[1455] = {-9'd70,-10'd271};
ram[1456] = {-9'd67,-10'd268};
ram[1457] = {-9'd64,-10'd264};
ram[1458] = {-9'd61,-10'd261};
ram[1459] = {-9'd58,-10'd258};
ram[1460] = {-9'd55,-10'd255};
ram[1461] = {-9'd52,-10'd252};
ram[1462] = {-9'd48,-10'd249};
ram[1463] = {-9'd45,-10'd246};
ram[1464] = {-9'd42,-10'd242};
ram[1465] = {-9'd39,-10'd239};
ram[1466] = {-9'd36,-10'd236};
ram[1467] = {-9'd33,-10'd233};
ram[1468] = {-9'd30,-10'd230};
ram[1469] = {-9'd26,-10'd227};
ram[1470] = {-9'd23,-10'd224};
ram[1471] = {-9'd20,-10'd220};
ram[1472] = {-9'd17,-10'd217};
ram[1473] = {-9'd14,-10'd214};
ram[1474] = {-9'd11,-10'd211};
ram[1475] = {-9'd8,-10'd208};
ram[1476] = {-9'd4,-10'd205};
ram[1477] = {-9'd1,-10'd202};
ram[1478] = {9'd2,-10'd198};
ram[1479] = {9'd5,-10'd195};
ram[1480] = {9'd8,-10'd192};
ram[1481] = {9'd11,-10'd189};
ram[1482] = {9'd14,-10'd186};
ram[1483] = {9'd18,-10'd183};
ram[1484] = {9'd21,-10'd180};
ram[1485] = {9'd24,-10'd176};
ram[1486] = {9'd27,-10'd173};
ram[1487] = {9'd30,-10'd170};
ram[1488] = {9'd33,-10'd167};
ram[1489] = {9'd36,-10'd164};
ram[1490] = {9'd40,-10'd161};
ram[1491] = {9'd43,-10'd158};
ram[1492] = {9'd46,-10'd154};
ram[1493] = {9'd49,-10'd151};
ram[1494] = {9'd52,-10'd148};
ram[1495] = {9'd55,-10'd145};
ram[1496] = {9'd58,-10'd142};
ram[1497] = {9'd62,-10'd139};
ram[1498] = {9'd65,-10'd136};
ram[1499] = {9'd68,-10'd132};
ram[1500] = {9'd71,-10'd129};
ram[1501] = {9'd74,-10'd126};
ram[1502] = {9'd77,-10'd123};
ram[1503] = {9'd80,-10'd120};
ram[1504] = {9'd84,-10'd117};
ram[1505] = {9'd87,-10'd114};
ram[1506] = {9'd90,-10'd110};
ram[1507] = {9'd93,-10'd107};
ram[1508] = {9'd96,-10'd104};
ram[1509] = {9'd99,-10'd101};
ram[1510] = {-9'd98,-10'd98};
ram[1511] = {-9'd95,-10'd95};
ram[1512] = {-9'd92,-10'd92};
ram[1513] = {-9'd88,-10'd88};
ram[1514] = {-9'd85,-10'd85};
ram[1515] = {-9'd82,-10'd82};
ram[1516] = {-9'd79,-10'd79};
ram[1517] = {-9'd76,-10'd76};
ram[1518] = {-9'd73,-10'd73};
ram[1519] = {-9'd70,-10'd70};
ram[1520] = {-9'd66,-10'd66};
ram[1521] = {-9'd63,-10'd63};
ram[1522] = {-9'd60,-10'd60};
ram[1523] = {-9'd57,-10'd57};
ram[1524] = {-9'd54,-10'd54};
ram[1525] = {-9'd51,-10'd51};
ram[1526] = {-9'd48,-10'd48};
ram[1527] = {-9'd44,-10'd44};
ram[1528] = {-9'd41,-10'd41};
ram[1529] = {-9'd38,-10'd38};
ram[1530] = {-9'd35,-10'd35};
ram[1531] = {-9'd32,-10'd32};
ram[1532] = {-9'd29,-10'd29};
ram[1533] = {-9'd26,-10'd26};
ram[1534] = {-9'd22,-10'd22};
ram[1535] = {-9'd19,-10'd19};
ram[1536] = {-9'd19,-10'd19};
ram[1537] = {-9'd16,-10'd16};
ram[1538] = {-9'd13,-10'd13};
ram[1539] = {-9'd10,-10'd10};
ram[1540] = {-9'd7,-10'd7};
ram[1541] = {-9'd4,-10'd4};
ram[1542] = {9'd0,10'd0};
ram[1543] = {9'd3,10'd3};
ram[1544] = {9'd6,10'd6};
ram[1545] = {9'd9,10'd9};
ram[1546] = {9'd12,10'd12};
ram[1547] = {9'd15,10'd15};
ram[1548] = {9'd18,10'd18};
ram[1549] = {9'd21,10'd21};
ram[1550] = {9'd25,10'd25};
ram[1551] = {9'd28,10'd28};
ram[1552] = {9'd31,10'd31};
ram[1553] = {9'd34,10'd34};
ram[1554] = {9'd37,10'd37};
ram[1555] = {9'd40,10'd40};
ram[1556] = {9'd43,10'd43};
ram[1557] = {9'd47,10'd47};
ram[1558] = {9'd50,10'd50};
ram[1559] = {9'd53,10'd53};
ram[1560] = {9'd56,10'd56};
ram[1561] = {9'd59,10'd59};
ram[1562] = {9'd62,10'd62};
ram[1563] = {9'd65,10'd65};
ram[1564] = {9'd69,10'd69};
ram[1565] = {9'd72,10'd72};
ram[1566] = {9'd75,10'd75};
ram[1567] = {9'd78,10'd78};
ram[1568] = {9'd81,10'd81};
ram[1569] = {9'd84,10'd84};
ram[1570] = {9'd87,10'd87};
ram[1571] = {9'd91,10'd91};
ram[1572] = {9'd94,10'd94};
ram[1573] = {9'd97,10'd97};
ram[1574] = {-9'd100,10'd100};
ram[1575] = {-9'd97,10'd103};
ram[1576] = {-9'd94,10'd106};
ram[1577] = {-9'd91,10'd109};
ram[1578] = {-9'd88,10'd113};
ram[1579] = {-9'd85,10'd116};
ram[1580] = {-9'd81,10'd119};
ram[1581] = {-9'd78,10'd122};
ram[1582] = {-9'd75,10'd125};
ram[1583] = {-9'd72,10'd128};
ram[1584] = {-9'd69,10'd131};
ram[1585] = {-9'd66,10'd135};
ram[1586] = {-9'd63,10'd138};
ram[1587] = {-9'd59,10'd141};
ram[1588] = {-9'd56,10'd144};
ram[1589] = {-9'd53,10'd147};
ram[1590] = {-9'd50,10'd150};
ram[1591] = {-9'd47,10'd153};
ram[1592] = {-9'd44,10'd157};
ram[1593] = {-9'd41,10'd160};
ram[1594] = {-9'd37,10'd163};
ram[1595] = {-9'd34,10'd166};
ram[1596] = {-9'd31,10'd169};
ram[1597] = {-9'd28,10'd172};
ram[1598] = {-9'd25,10'd175};
ram[1599] = {-9'd22,10'd179};
ram[1600] = {-9'd19,10'd182};
ram[1601] = {-9'd15,10'd185};
ram[1602] = {-9'd12,10'd188};
ram[1603] = {-9'd9,10'd191};
ram[1604] = {-9'd6,10'd194};
ram[1605] = {-9'd3,10'd197};
ram[1606] = {9'd0,10'd201};
ram[1607] = {9'd3,10'd204};
ram[1608] = {9'd7,10'd207};
ram[1609] = {9'd10,10'd210};
ram[1610] = {9'd13,10'd213};
ram[1611] = {9'd16,10'd216};
ram[1612] = {9'd19,10'd219};
ram[1613] = {9'd22,10'd223};
ram[1614] = {9'd25,10'd226};
ram[1615] = {9'd29,10'd229};
ram[1616] = {9'd32,10'd232};
ram[1617] = {9'd35,10'd235};
ram[1618] = {9'd38,10'd238};
ram[1619] = {9'd41,10'd241};
ram[1620] = {9'd44,10'd245};
ram[1621] = {9'd47,10'd248};
ram[1622] = {9'd51,10'd251};
ram[1623] = {9'd54,10'd254};
ram[1624] = {9'd57,10'd257};
ram[1625] = {9'd60,10'd260};
ram[1626] = {9'd63,10'd263};
ram[1627] = {9'd66,10'd267};
ram[1628] = {9'd69,10'd270};
ram[1629] = {9'd73,10'd273};
ram[1630] = {9'd76,10'd276};
ram[1631] = {9'd79,10'd279};
ram[1632] = {9'd82,10'd282};
ram[1633] = {9'd85,10'd285};
ram[1634] = {9'd88,10'd289};
ram[1635] = {9'd91,10'd292};
ram[1636] = {9'd95,10'd295};
ram[1637] = {9'd98,10'd298};
ram[1638] = {-9'd99,10'd301};
ram[1639] = {-9'd96,10'd304};
ram[1640] = {-9'd93,10'd307};
ram[1641] = {-9'd90,10'd311};
ram[1642] = {-9'd87,10'd314};
ram[1643] = {-9'd84,10'd317};
ram[1644] = {-9'd81,10'd320};
ram[1645] = {-9'd77,10'd323};
ram[1646] = {-9'd74,10'd326};
ram[1647] = {-9'd71,10'd329};
ram[1648] = {-9'd68,10'd333};
ram[1649] = {-9'd65,10'd336};
ram[1650] = {-9'd62,10'd339};
ram[1651] = {-9'd59,10'd342};
ram[1652] = {-9'd55,10'd345};
ram[1653] = {-9'd52,10'd348};
ram[1654] = {-9'd49,10'd351};
ram[1655] = {-9'd46,10'd354};
ram[1656] = {-9'd43,10'd358};
ram[1657] = {-9'd40,10'd361};
ram[1658] = {-9'd37,10'd364};
ram[1659] = {-9'd33,10'd367};
ram[1660] = {-9'd30,10'd370};
ram[1661] = {-9'd27,10'd373};
ram[1662] = {-9'd24,10'd376};
ram[1663] = {-9'd21,10'd380};
ram[1664] = {-9'd21,10'd380};
ram[1665] = {-9'd18,10'd383};
ram[1666] = {-9'd15,10'd386};
ram[1667] = {-9'd11,10'd389};
ram[1668] = {-9'd8,10'd392};
ram[1669] = {-9'd5,10'd395};
ram[1670] = {-9'd2,10'd398};
ram[1671] = {9'd1,-10'd399};
ram[1672] = {9'd4,-10'd396};
ram[1673] = {9'd7,-10'd393};
ram[1674] = {9'd10,-10'd390};
ram[1675] = {9'd14,-10'd387};
ram[1676] = {9'd17,-10'd384};
ram[1677] = {9'd20,-10'd381};
ram[1678] = {9'd23,-10'd377};
ram[1679] = {9'd26,-10'd374};
ram[1680] = {9'd29,-10'd371};
ram[1681] = {9'd32,-10'd368};
ram[1682] = {9'd36,-10'd365};
ram[1683] = {9'd39,-10'd362};
ram[1684] = {9'd42,-10'd359};
ram[1685] = {9'd45,-10'd355};
ram[1686] = {9'd48,-10'd352};
ram[1687] = {9'd51,-10'd349};
ram[1688] = {9'd54,-10'd346};
ram[1689] = {9'd58,-10'd343};
ram[1690] = {9'd61,-10'd340};
ram[1691] = {9'd64,-10'd337};
ram[1692] = {9'd67,-10'd334};
ram[1693] = {9'd70,-10'd330};
ram[1694] = {9'd73,-10'd327};
ram[1695] = {9'd76,-10'd324};
ram[1696] = {9'd80,-10'd321};
ram[1697] = {9'd83,-10'd318};
ram[1698] = {9'd86,-10'd315};
ram[1699] = {9'd89,-10'd312};
ram[1700] = {9'd92,-10'd308};
ram[1701] = {9'd95,-10'd305};
ram[1702] = {9'd98,-10'd302};
ram[1703] = {-9'd99,-10'd299};
ram[1704] = {-9'd96,-10'd296};
ram[1705] = {-9'd92,-10'd293};
ram[1706] = {-9'd89,-10'd290};
ram[1707] = {-9'd86,-10'd286};
ram[1708] = {-9'd83,-10'd283};
ram[1709] = {-9'd80,-10'd280};
ram[1710] = {-9'd77,-10'd277};
ram[1711] = {-9'd74,-10'd274};
ram[1712] = {-9'd70,-10'd271};
ram[1713] = {-9'd67,-10'd268};
ram[1714] = {-9'd64,-10'd264};
ram[1715] = {-9'd61,-10'd261};
ram[1716] = {-9'd58,-10'd258};
ram[1717] = {-9'd55,-10'd255};
ram[1718] = {-9'd52,-10'd252};
ram[1719] = {-9'd48,-10'd249};
ram[1720] = {-9'd45,-10'd246};
ram[1721] = {-9'd42,-10'd242};
ram[1722] = {-9'd39,-10'd239};
ram[1723] = {-9'd36,-10'd236};
ram[1724] = {-9'd33,-10'd233};
ram[1725] = {-9'd30,-10'd230};
ram[1726] = {-9'd26,-10'd227};
ram[1727] = {-9'd23,-10'd224};
ram[1728] = {-9'd20,-10'd220};
ram[1729] = {-9'd17,-10'd217};
ram[1730] = {-9'd14,-10'd214};
ram[1731] = {-9'd11,-10'd211};
ram[1732] = {-9'd8,-10'd208};
ram[1733] = {-9'd4,-10'd205};
ram[1734] = {-9'd1,-10'd202};
ram[1735] = {9'd2,-10'd198};
ram[1736] = {9'd5,-10'd195};
ram[1737] = {9'd8,-10'd192};
ram[1738] = {9'd11,-10'd189};
ram[1739] = {9'd14,-10'd186};
ram[1740] = {9'd18,-10'd183};
ram[1741] = {9'd21,-10'd180};
ram[1742] = {9'd24,-10'd176};
ram[1743] = {9'd27,-10'd173};
ram[1744] = {9'd30,-10'd170};
ram[1745] = {9'd33,-10'd167};
ram[1746] = {9'd36,-10'd164};
ram[1747] = {9'd40,-10'd161};
ram[1748] = {9'd43,-10'd158};
ram[1749] = {9'd46,-10'd154};
ram[1750] = {9'd49,-10'd151};
ram[1751] = {9'd52,-10'd148};
ram[1752] = {9'd55,-10'd145};
ram[1753] = {9'd58,-10'd142};
ram[1754] = {9'd62,-10'd139};
ram[1755] = {9'd65,-10'd136};
ram[1756] = {9'd68,-10'd132};
ram[1757] = {9'd71,-10'd129};
ram[1758] = {9'd74,-10'd126};
ram[1759] = {9'd77,-10'd123};
ram[1760] = {9'd80,-10'd120};
ram[1761] = {9'd84,-10'd117};
ram[1762] = {9'd87,-10'd114};
ram[1763] = {9'd90,-10'd110};
ram[1764] = {9'd93,-10'd107};
ram[1765] = {9'd96,-10'd104};
ram[1766] = {9'd99,-10'd101};
ram[1767] = {-9'd98,-10'd98};
ram[1768] = {-9'd95,-10'd95};
ram[1769] = {-9'd92,-10'd92};
ram[1770] = {-9'd88,-10'd88};
ram[1771] = {-9'd85,-10'd85};
ram[1772] = {-9'd82,-10'd82};
ram[1773] = {-9'd79,-10'd79};
ram[1774] = {-9'd76,-10'd76};
ram[1775] = {-9'd73,-10'd73};
ram[1776] = {-9'd70,-10'd70};
ram[1777] = {-9'd66,-10'd66};
ram[1778] = {-9'd63,-10'd63};
ram[1779] = {-9'd60,-10'd60};
ram[1780] = {-9'd57,-10'd57};
ram[1781] = {-9'd54,-10'd54};
ram[1782] = {-9'd51,-10'd51};
ram[1783] = {-9'd48,-10'd48};
ram[1784] = {-9'd44,-10'd44};
ram[1785] = {-9'd41,-10'd41};
ram[1786] = {-9'd38,-10'd38};
ram[1787] = {-9'd35,-10'd35};
ram[1788] = {-9'd32,-10'd32};
ram[1789] = {-9'd29,-10'd29};
ram[1790] = {-9'd26,-10'd26};
ram[1791] = {-9'd22,-10'd22};
ram[1792] = {-9'd22,-10'd22};
ram[1793] = {-9'd19,-10'd19};
ram[1794] = {-9'd16,-10'd16};
ram[1795] = {-9'd13,-10'd13};
ram[1796] = {-9'd10,-10'd10};
ram[1797] = {-9'd7,-10'd7};
ram[1798] = {-9'd4,-10'd4};
ram[1799] = {9'd0,10'd0};
ram[1800] = {9'd3,10'd3};
ram[1801] = {9'd6,10'd6};
ram[1802] = {9'd9,10'd9};
ram[1803] = {9'd12,10'd12};
ram[1804] = {9'd15,10'd15};
ram[1805] = {9'd18,10'd18};
ram[1806] = {9'd21,10'd21};
ram[1807] = {9'd25,10'd25};
ram[1808] = {9'd28,10'd28};
ram[1809] = {9'd31,10'd31};
ram[1810] = {9'd34,10'd34};
ram[1811] = {9'd37,10'd37};
ram[1812] = {9'd40,10'd40};
ram[1813] = {9'd43,10'd43};
ram[1814] = {9'd47,10'd47};
ram[1815] = {9'd50,10'd50};
ram[1816] = {9'd53,10'd53};
ram[1817] = {9'd56,10'd56};
ram[1818] = {9'd59,10'd59};
ram[1819] = {9'd62,10'd62};
ram[1820] = {9'd65,10'd65};
ram[1821] = {9'd69,10'd69};
ram[1822] = {9'd72,10'd72};
ram[1823] = {9'd75,10'd75};
ram[1824] = {9'd78,10'd78};
ram[1825] = {9'd81,10'd81};
ram[1826] = {9'd84,10'd84};
ram[1827] = {9'd87,10'd87};
ram[1828] = {9'd91,10'd91};
ram[1829] = {9'd94,10'd94};
ram[1830] = {9'd97,10'd97};
ram[1831] = {-9'd100,10'd100};
ram[1832] = {-9'd97,10'd103};
ram[1833] = {-9'd94,10'd106};
ram[1834] = {-9'd91,10'd109};
ram[1835] = {-9'd88,10'd113};
ram[1836] = {-9'd85,10'd116};
ram[1837] = {-9'd81,10'd119};
ram[1838] = {-9'd78,10'd122};
ram[1839] = {-9'd75,10'd125};
ram[1840] = {-9'd72,10'd128};
ram[1841] = {-9'd69,10'd131};
ram[1842] = {-9'd66,10'd135};
ram[1843] = {-9'd63,10'd138};
ram[1844] = {-9'd59,10'd141};
ram[1845] = {-9'd56,10'd144};
ram[1846] = {-9'd53,10'd147};
ram[1847] = {-9'd50,10'd150};
ram[1848] = {-9'd47,10'd153};
ram[1849] = {-9'd44,10'd157};
ram[1850] = {-9'd41,10'd160};
ram[1851] = {-9'd37,10'd163};
ram[1852] = {-9'd34,10'd166};
ram[1853] = {-9'd31,10'd169};
ram[1854] = {-9'd28,10'd172};
ram[1855] = {-9'd25,10'd175};
ram[1856] = {-9'd22,10'd179};
ram[1857] = {-9'd19,10'd182};
ram[1858] = {-9'd15,10'd185};
ram[1859] = {-9'd12,10'd188};
ram[1860] = {-9'd9,10'd191};
ram[1861] = {-9'd6,10'd194};
ram[1862] = {-9'd3,10'd197};
ram[1863] = {9'd0,10'd201};
ram[1864] = {9'd3,10'd204};
ram[1865] = {9'd7,10'd207};
ram[1866] = {9'd10,10'd210};
ram[1867] = {9'd13,10'd213};
ram[1868] = {9'd16,10'd216};
ram[1869] = {9'd19,10'd219};
ram[1870] = {9'd22,10'd223};
ram[1871] = {9'd25,10'd226};
ram[1872] = {9'd29,10'd229};
ram[1873] = {9'd32,10'd232};
ram[1874] = {9'd35,10'd235};
ram[1875] = {9'd38,10'd238};
ram[1876] = {9'd41,10'd241};
ram[1877] = {9'd44,10'd245};
ram[1878] = {9'd47,10'd248};
ram[1879] = {9'd51,10'd251};
ram[1880] = {9'd54,10'd254};
ram[1881] = {9'd57,10'd257};
ram[1882] = {9'd60,10'd260};
ram[1883] = {9'd63,10'd263};
ram[1884] = {9'd66,10'd267};
ram[1885] = {9'd69,10'd270};
ram[1886] = {9'd73,10'd273};
ram[1887] = {9'd76,10'd276};
ram[1888] = {9'd79,10'd279};
ram[1889] = {9'd82,10'd282};
ram[1890] = {9'd85,10'd285};
ram[1891] = {9'd88,10'd289};
ram[1892] = {9'd91,10'd292};
ram[1893] = {9'd95,10'd295};
ram[1894] = {9'd98,10'd298};
ram[1895] = {-9'd99,10'd301};
ram[1896] = {-9'd96,10'd304};
ram[1897] = {-9'd93,10'd307};
ram[1898] = {-9'd90,10'd311};
ram[1899] = {-9'd87,10'd314};
ram[1900] = {-9'd84,10'd317};
ram[1901] = {-9'd81,10'd320};
ram[1902] = {-9'd77,10'd323};
ram[1903] = {-9'd74,10'd326};
ram[1904] = {-9'd71,10'd329};
ram[1905] = {-9'd68,10'd333};
ram[1906] = {-9'd65,10'd336};
ram[1907] = {-9'd62,10'd339};
ram[1908] = {-9'd59,10'd342};
ram[1909] = {-9'd55,10'd345};
ram[1910] = {-9'd52,10'd348};
ram[1911] = {-9'd49,10'd351};
ram[1912] = {-9'd46,10'd354};
ram[1913] = {-9'd43,10'd358};
ram[1914] = {-9'd40,10'd361};
ram[1915] = {-9'd37,10'd364};
ram[1916] = {-9'd33,10'd367};
ram[1917] = {-9'd30,10'd370};
ram[1918] = {-9'd27,10'd373};
ram[1919] = {-9'd24,10'd376};
ram[1920] = {-9'd24,10'd376};
ram[1921] = {-9'd21,10'd380};
ram[1922] = {-9'd18,10'd383};
ram[1923] = {-9'd15,10'd386};
ram[1924] = {-9'd11,10'd389};
ram[1925] = {-9'd8,10'd392};
ram[1926] = {-9'd5,10'd395};
ram[1927] = {-9'd2,10'd398};
ram[1928] = {9'd1,-10'd399};
ram[1929] = {9'd4,-10'd396};
ram[1930] = {9'd7,-10'd393};
ram[1931] = {9'd10,-10'd390};
ram[1932] = {9'd14,-10'd387};
ram[1933] = {9'd17,-10'd384};
ram[1934] = {9'd20,-10'd381};
ram[1935] = {9'd23,-10'd377};
ram[1936] = {9'd26,-10'd374};
ram[1937] = {9'd29,-10'd371};
ram[1938] = {9'd32,-10'd368};
ram[1939] = {9'd36,-10'd365};
ram[1940] = {9'd39,-10'd362};
ram[1941] = {9'd42,-10'd359};
ram[1942] = {9'd45,-10'd355};
ram[1943] = {9'd48,-10'd352};
ram[1944] = {9'd51,-10'd349};
ram[1945] = {9'd54,-10'd346};
ram[1946] = {9'd58,-10'd343};
ram[1947] = {9'd61,-10'd340};
ram[1948] = {9'd64,-10'd337};
ram[1949] = {9'd67,-10'd334};
ram[1950] = {9'd70,-10'd330};
ram[1951] = {9'd73,-10'd327};
ram[1952] = {9'd76,-10'd324};
ram[1953] = {9'd80,-10'd321};
ram[1954] = {9'd83,-10'd318};
ram[1955] = {9'd86,-10'd315};
ram[1956] = {9'd89,-10'd312};
ram[1957] = {9'd92,-10'd308};
ram[1958] = {9'd95,-10'd305};
ram[1959] = {9'd98,-10'd302};
ram[1960] = {-9'd99,-10'd299};
ram[1961] = {-9'd96,-10'd296};
ram[1962] = {-9'd92,-10'd293};
ram[1963] = {-9'd89,-10'd290};
ram[1964] = {-9'd86,-10'd286};
ram[1965] = {-9'd83,-10'd283};
ram[1966] = {-9'd80,-10'd280};
ram[1967] = {-9'd77,-10'd277};
ram[1968] = {-9'd74,-10'd274};
ram[1969] = {-9'd70,-10'd271};
ram[1970] = {-9'd67,-10'd268};
ram[1971] = {-9'd64,-10'd264};
ram[1972] = {-9'd61,-10'd261};
ram[1973] = {-9'd58,-10'd258};
ram[1974] = {-9'd55,-10'd255};
ram[1975] = {-9'd52,-10'd252};
ram[1976] = {-9'd48,-10'd249};
ram[1977] = {-9'd45,-10'd246};
ram[1978] = {-9'd42,-10'd242};
ram[1979] = {-9'd39,-10'd239};
ram[1980] = {-9'd36,-10'd236};
ram[1981] = {-9'd33,-10'd233};
ram[1982] = {-9'd30,-10'd230};
ram[1983] = {-9'd26,-10'd227};
ram[1984] = {-9'd23,-10'd224};
ram[1985] = {-9'd20,-10'd220};
ram[1986] = {-9'd17,-10'd217};
ram[1987] = {-9'd14,-10'd214};
ram[1988] = {-9'd11,-10'd211};
ram[1989] = {-9'd8,-10'd208};
ram[1990] = {-9'd4,-10'd205};
ram[1991] = {-9'd1,-10'd202};
ram[1992] = {9'd2,-10'd198};
ram[1993] = {9'd5,-10'd195};
ram[1994] = {9'd8,-10'd192};
ram[1995] = {9'd11,-10'd189};
ram[1996] = {9'd14,-10'd186};
ram[1997] = {9'd18,-10'd183};
ram[1998] = {9'd21,-10'd180};
ram[1999] = {9'd24,-10'd176};
ram[2000] = {9'd27,-10'd173};
ram[2001] = {9'd30,-10'd170};
ram[2002] = {9'd33,-10'd167};
ram[2003] = {9'd36,-10'd164};
ram[2004] = {9'd40,-10'd161};
ram[2005] = {9'd43,-10'd158};
ram[2006] = {9'd46,-10'd154};
ram[2007] = {9'd49,-10'd151};
ram[2008] = {9'd52,-10'd148};
ram[2009] = {9'd55,-10'd145};
ram[2010] = {9'd58,-10'd142};
ram[2011] = {9'd62,-10'd139};
ram[2012] = {9'd65,-10'd136};
ram[2013] = {9'd68,-10'd132};
ram[2014] = {9'd71,-10'd129};
ram[2015] = {9'd74,-10'd126};
ram[2016] = {9'd77,-10'd123};
ram[2017] = {9'd80,-10'd120};
ram[2018] = {9'd84,-10'd117};
ram[2019] = {9'd87,-10'd114};
ram[2020] = {9'd90,-10'd110};
ram[2021] = {9'd93,-10'd107};
ram[2022] = {9'd96,-10'd104};
ram[2023] = {9'd99,-10'd101};
ram[2024] = {-9'd98,-10'd98};
ram[2025] = {-9'd95,-10'd95};
ram[2026] = {-9'd92,-10'd92};
ram[2027] = {-9'd88,-10'd88};
ram[2028] = {-9'd85,-10'd85};
ram[2029] = {-9'd82,-10'd82};
ram[2030] = {-9'd79,-10'd79};
ram[2031] = {-9'd76,-10'd76};
ram[2032] = {-9'd73,-10'd73};
ram[2033] = {-9'd70,-10'd70};
ram[2034] = {-9'd66,-10'd66};
ram[2035] = {-9'd63,-10'd63};
ram[2036] = {-9'd60,-10'd60};
ram[2037] = {-9'd57,-10'd57};
ram[2038] = {-9'd54,-10'd54};
ram[2039] = {-9'd51,-10'd51};
ram[2040] = {-9'd48,-10'd48};
ram[2041] = {-9'd44,-10'd44};
ram[2042] = {-9'd41,-10'd41};
ram[2043] = {-9'd38,-10'd38};
ram[2044] = {-9'd35,-10'd35};
ram[2045] = {-9'd32,-10'd32};
ram[2046] = {-9'd29,-10'd29};
ram[2047] = {-9'd26,-10'd26};
ram[2048] = {-9'd26,-10'd26};
ram[2049] = {-9'd22,-10'd22};
ram[2050] = {-9'd19,-10'd19};
ram[2051] = {-9'd16,-10'd16};
ram[2052] = {-9'd13,-10'd13};
ram[2053] = {-9'd10,-10'd10};
ram[2054] = {-9'd7,-10'd7};
ram[2055] = {-9'd4,-10'd4};
ram[2056] = {9'd0,10'd0};
ram[2057] = {9'd3,10'd3};
ram[2058] = {9'd6,10'd6};
ram[2059] = {9'd9,10'd9};
ram[2060] = {9'd12,10'd12};
ram[2061] = {9'd15,10'd15};
ram[2062] = {9'd18,10'd18};
ram[2063] = {9'd21,10'd21};
ram[2064] = {9'd25,10'd25};
ram[2065] = {9'd28,10'd28};
ram[2066] = {9'd31,10'd31};
ram[2067] = {9'd34,10'd34};
ram[2068] = {9'd37,10'd37};
ram[2069] = {9'd40,10'd40};
ram[2070] = {9'd43,10'd43};
ram[2071] = {9'd47,10'd47};
ram[2072] = {9'd50,10'd50};
ram[2073] = {9'd53,10'd53};
ram[2074] = {9'd56,10'd56};
ram[2075] = {9'd59,10'd59};
ram[2076] = {9'd62,10'd62};
ram[2077] = {9'd65,10'd65};
ram[2078] = {9'd69,10'd69};
ram[2079] = {9'd72,10'd72};
ram[2080] = {9'd75,10'd75};
ram[2081] = {9'd78,10'd78};
ram[2082] = {9'd81,10'd81};
ram[2083] = {9'd84,10'd84};
ram[2084] = {9'd87,10'd87};
ram[2085] = {9'd91,10'd91};
ram[2086] = {9'd94,10'd94};
ram[2087] = {9'd97,10'd97};
ram[2088] = {-9'd100,10'd100};
ram[2089] = {-9'd97,10'd103};
ram[2090] = {-9'd94,10'd106};
ram[2091] = {-9'd91,10'd109};
ram[2092] = {-9'd88,10'd113};
ram[2093] = {-9'd85,10'd116};
ram[2094] = {-9'd81,10'd119};
ram[2095] = {-9'd78,10'd122};
ram[2096] = {-9'd75,10'd125};
ram[2097] = {-9'd72,10'd128};
ram[2098] = {-9'd69,10'd131};
ram[2099] = {-9'd66,10'd135};
ram[2100] = {-9'd63,10'd138};
ram[2101] = {-9'd59,10'd141};
ram[2102] = {-9'd56,10'd144};
ram[2103] = {-9'd53,10'd147};
ram[2104] = {-9'd50,10'd150};
ram[2105] = {-9'd47,10'd153};
ram[2106] = {-9'd44,10'd157};
ram[2107] = {-9'd41,10'd160};
ram[2108] = {-9'd37,10'd163};
ram[2109] = {-9'd34,10'd166};
ram[2110] = {-9'd31,10'd169};
ram[2111] = {-9'd28,10'd172};
ram[2112] = {-9'd25,10'd175};
ram[2113] = {-9'd22,10'd179};
ram[2114] = {-9'd19,10'd182};
ram[2115] = {-9'd15,10'd185};
ram[2116] = {-9'd12,10'd188};
ram[2117] = {-9'd9,10'd191};
ram[2118] = {-9'd6,10'd194};
ram[2119] = {-9'd3,10'd197};
ram[2120] = {9'd0,10'd201};
ram[2121] = {9'd3,10'd204};
ram[2122] = {9'd7,10'd207};
ram[2123] = {9'd10,10'd210};
ram[2124] = {9'd13,10'd213};
ram[2125] = {9'd16,10'd216};
ram[2126] = {9'd19,10'd219};
ram[2127] = {9'd22,10'd223};
ram[2128] = {9'd25,10'd226};
ram[2129] = {9'd29,10'd229};
ram[2130] = {9'd32,10'd232};
ram[2131] = {9'd35,10'd235};
ram[2132] = {9'd38,10'd238};
ram[2133] = {9'd41,10'd241};
ram[2134] = {9'd44,10'd245};
ram[2135] = {9'd47,10'd248};
ram[2136] = {9'd51,10'd251};
ram[2137] = {9'd54,10'd254};
ram[2138] = {9'd57,10'd257};
ram[2139] = {9'd60,10'd260};
ram[2140] = {9'd63,10'd263};
ram[2141] = {9'd66,10'd267};
ram[2142] = {9'd69,10'd270};
ram[2143] = {9'd73,10'd273};
ram[2144] = {9'd76,10'd276};
ram[2145] = {9'd79,10'd279};
ram[2146] = {9'd82,10'd282};
ram[2147] = {9'd85,10'd285};
ram[2148] = {9'd88,10'd289};
ram[2149] = {9'd91,10'd292};
ram[2150] = {9'd95,10'd295};
ram[2151] = {9'd98,10'd298};
ram[2152] = {-9'd99,10'd301};
ram[2153] = {-9'd96,10'd304};
ram[2154] = {-9'd93,10'd307};
ram[2155] = {-9'd90,10'd311};
ram[2156] = {-9'd87,10'd314};
ram[2157] = {-9'd84,10'd317};
ram[2158] = {-9'd81,10'd320};
ram[2159] = {-9'd77,10'd323};
ram[2160] = {-9'd74,10'd326};
ram[2161] = {-9'd71,10'd329};
ram[2162] = {-9'd68,10'd333};
ram[2163] = {-9'd65,10'd336};
ram[2164] = {-9'd62,10'd339};
ram[2165] = {-9'd59,10'd342};
ram[2166] = {-9'd55,10'd345};
ram[2167] = {-9'd52,10'd348};
ram[2168] = {-9'd49,10'd351};
ram[2169] = {-9'd46,10'd354};
ram[2170] = {-9'd43,10'd358};
ram[2171] = {-9'd40,10'd361};
ram[2172] = {-9'd37,10'd364};
ram[2173] = {-9'd33,10'd367};
ram[2174] = {-9'd30,10'd370};
ram[2175] = {-9'd27,10'd373};
ram[2176] = {-9'd27,10'd373};
ram[2177] = {-9'd24,10'd376};
ram[2178] = {-9'd21,10'd380};
ram[2179] = {-9'd18,10'd383};
ram[2180] = {-9'd15,10'd386};
ram[2181] = {-9'd11,10'd389};
ram[2182] = {-9'd8,10'd392};
ram[2183] = {-9'd5,10'd395};
ram[2184] = {-9'd2,10'd398};
ram[2185] = {9'd1,-10'd399};
ram[2186] = {9'd4,-10'd396};
ram[2187] = {9'd7,-10'd393};
ram[2188] = {9'd10,-10'd390};
ram[2189] = {9'd14,-10'd387};
ram[2190] = {9'd17,-10'd384};
ram[2191] = {9'd20,-10'd381};
ram[2192] = {9'd23,-10'd377};
ram[2193] = {9'd26,-10'd374};
ram[2194] = {9'd29,-10'd371};
ram[2195] = {9'd32,-10'd368};
ram[2196] = {9'd36,-10'd365};
ram[2197] = {9'd39,-10'd362};
ram[2198] = {9'd42,-10'd359};
ram[2199] = {9'd45,-10'd355};
ram[2200] = {9'd48,-10'd352};
ram[2201] = {9'd51,-10'd349};
ram[2202] = {9'd54,-10'd346};
ram[2203] = {9'd58,-10'd343};
ram[2204] = {9'd61,-10'd340};
ram[2205] = {9'd64,-10'd337};
ram[2206] = {9'd67,-10'd334};
ram[2207] = {9'd70,-10'd330};
ram[2208] = {9'd73,-10'd327};
ram[2209] = {9'd76,-10'd324};
ram[2210] = {9'd80,-10'd321};
ram[2211] = {9'd83,-10'd318};
ram[2212] = {9'd86,-10'd315};
ram[2213] = {9'd89,-10'd312};
ram[2214] = {9'd92,-10'd308};
ram[2215] = {9'd95,-10'd305};
ram[2216] = {9'd98,-10'd302};
ram[2217] = {-9'd99,-10'd299};
ram[2218] = {-9'd96,-10'd296};
ram[2219] = {-9'd92,-10'd293};
ram[2220] = {-9'd89,-10'd290};
ram[2221] = {-9'd86,-10'd286};
ram[2222] = {-9'd83,-10'd283};
ram[2223] = {-9'd80,-10'd280};
ram[2224] = {-9'd77,-10'd277};
ram[2225] = {-9'd74,-10'd274};
ram[2226] = {-9'd70,-10'd271};
ram[2227] = {-9'd67,-10'd268};
ram[2228] = {-9'd64,-10'd264};
ram[2229] = {-9'd61,-10'd261};
ram[2230] = {-9'd58,-10'd258};
ram[2231] = {-9'd55,-10'd255};
ram[2232] = {-9'd52,-10'd252};
ram[2233] = {-9'd48,-10'd249};
ram[2234] = {-9'd45,-10'd246};
ram[2235] = {-9'd42,-10'd242};
ram[2236] = {-9'd39,-10'd239};
ram[2237] = {-9'd36,-10'd236};
ram[2238] = {-9'd33,-10'd233};
ram[2239] = {-9'd30,-10'd230};
ram[2240] = {-9'd26,-10'd227};
ram[2241] = {-9'd23,-10'd224};
ram[2242] = {-9'd20,-10'd220};
ram[2243] = {-9'd17,-10'd217};
ram[2244] = {-9'd14,-10'd214};
ram[2245] = {-9'd11,-10'd211};
ram[2246] = {-9'd8,-10'd208};
ram[2247] = {-9'd4,-10'd205};
ram[2248] = {-9'd1,-10'd202};
ram[2249] = {9'd2,-10'd198};
ram[2250] = {9'd5,-10'd195};
ram[2251] = {9'd8,-10'd192};
ram[2252] = {9'd11,-10'd189};
ram[2253] = {9'd14,-10'd186};
ram[2254] = {9'd18,-10'd183};
ram[2255] = {9'd21,-10'd180};
ram[2256] = {9'd24,-10'd176};
ram[2257] = {9'd27,-10'd173};
ram[2258] = {9'd30,-10'd170};
ram[2259] = {9'd33,-10'd167};
ram[2260] = {9'd36,-10'd164};
ram[2261] = {9'd40,-10'd161};
ram[2262] = {9'd43,-10'd158};
ram[2263] = {9'd46,-10'd154};
ram[2264] = {9'd49,-10'd151};
ram[2265] = {9'd52,-10'd148};
ram[2266] = {9'd55,-10'd145};
ram[2267] = {9'd58,-10'd142};
ram[2268] = {9'd62,-10'd139};
ram[2269] = {9'd65,-10'd136};
ram[2270] = {9'd68,-10'd132};
ram[2271] = {9'd71,-10'd129};
ram[2272] = {9'd74,-10'd126};
ram[2273] = {9'd77,-10'd123};
ram[2274] = {9'd80,-10'd120};
ram[2275] = {9'd84,-10'd117};
ram[2276] = {9'd87,-10'd114};
ram[2277] = {9'd90,-10'd110};
ram[2278] = {9'd93,-10'd107};
ram[2279] = {9'd96,-10'd104};
ram[2280] = {9'd99,-10'd101};
ram[2281] = {-9'd98,-10'd98};
ram[2282] = {-9'd95,-10'd95};
ram[2283] = {-9'd92,-10'd92};
ram[2284] = {-9'd88,-10'd88};
ram[2285] = {-9'd85,-10'd85};
ram[2286] = {-9'd82,-10'd82};
ram[2287] = {-9'd79,-10'd79};
ram[2288] = {-9'd76,-10'd76};
ram[2289] = {-9'd73,-10'd73};
ram[2290] = {-9'd70,-10'd70};
ram[2291] = {-9'd66,-10'd66};
ram[2292] = {-9'd63,-10'd63};
ram[2293] = {-9'd60,-10'd60};
ram[2294] = {-9'd57,-10'd57};
ram[2295] = {-9'd54,-10'd54};
ram[2296] = {-9'd51,-10'd51};
ram[2297] = {-9'd48,-10'd48};
ram[2298] = {-9'd44,-10'd44};
ram[2299] = {-9'd41,-10'd41};
ram[2300] = {-9'd38,-10'd38};
ram[2301] = {-9'd35,-10'd35};
ram[2302] = {-9'd32,-10'd32};
ram[2303] = {-9'd29,-10'd29};
ram[2304] = {-9'd29,-10'd29};
ram[2305] = {-9'd26,-10'd26};
ram[2306] = {-9'd22,-10'd22};
ram[2307] = {-9'd19,-10'd19};
ram[2308] = {-9'd16,-10'd16};
ram[2309] = {-9'd13,-10'd13};
ram[2310] = {-9'd10,-10'd10};
ram[2311] = {-9'd7,-10'd7};
ram[2312] = {-9'd4,-10'd4};
ram[2313] = {9'd0,10'd0};
ram[2314] = {9'd3,10'd3};
ram[2315] = {9'd6,10'd6};
ram[2316] = {9'd9,10'd9};
ram[2317] = {9'd12,10'd12};
ram[2318] = {9'd15,10'd15};
ram[2319] = {9'd18,10'd18};
ram[2320] = {9'd21,10'd21};
ram[2321] = {9'd25,10'd25};
ram[2322] = {9'd28,10'd28};
ram[2323] = {9'd31,10'd31};
ram[2324] = {9'd34,10'd34};
ram[2325] = {9'd37,10'd37};
ram[2326] = {9'd40,10'd40};
ram[2327] = {9'd43,10'd43};
ram[2328] = {9'd47,10'd47};
ram[2329] = {9'd50,10'd50};
ram[2330] = {9'd53,10'd53};
ram[2331] = {9'd56,10'd56};
ram[2332] = {9'd59,10'd59};
ram[2333] = {9'd62,10'd62};
ram[2334] = {9'd65,10'd65};
ram[2335] = {9'd69,10'd69};
ram[2336] = {9'd72,10'd72};
ram[2337] = {9'd75,10'd75};
ram[2338] = {9'd78,10'd78};
ram[2339] = {9'd81,10'd81};
ram[2340] = {9'd84,10'd84};
ram[2341] = {9'd87,10'd87};
ram[2342] = {9'd91,10'd91};
ram[2343] = {9'd94,10'd94};
ram[2344] = {9'd97,10'd97};
ram[2345] = {-9'd100,10'd100};
ram[2346] = {-9'd97,10'd103};
ram[2347] = {-9'd94,10'd106};
ram[2348] = {-9'd91,10'd109};
ram[2349] = {-9'd88,10'd113};
ram[2350] = {-9'd85,10'd116};
ram[2351] = {-9'd81,10'd119};
ram[2352] = {-9'd78,10'd122};
ram[2353] = {-9'd75,10'd125};
ram[2354] = {-9'd72,10'd128};
ram[2355] = {-9'd69,10'd131};
ram[2356] = {-9'd66,10'd135};
ram[2357] = {-9'd63,10'd138};
ram[2358] = {-9'd59,10'd141};
ram[2359] = {-9'd56,10'd144};
ram[2360] = {-9'd53,10'd147};
ram[2361] = {-9'd50,10'd150};
ram[2362] = {-9'd47,10'd153};
ram[2363] = {-9'd44,10'd157};
ram[2364] = {-9'd41,10'd160};
ram[2365] = {-9'd37,10'd163};
ram[2366] = {-9'd34,10'd166};
ram[2367] = {-9'd31,10'd169};
ram[2368] = {-9'd28,10'd172};
ram[2369] = {-9'd25,10'd175};
ram[2370] = {-9'd22,10'd179};
ram[2371] = {-9'd19,10'd182};
ram[2372] = {-9'd15,10'd185};
ram[2373] = {-9'd12,10'd188};
ram[2374] = {-9'd9,10'd191};
ram[2375] = {-9'd6,10'd194};
ram[2376] = {-9'd3,10'd197};
ram[2377] = {9'd0,10'd201};
ram[2378] = {9'd3,10'd204};
ram[2379] = {9'd7,10'd207};
ram[2380] = {9'd10,10'd210};
ram[2381] = {9'd13,10'd213};
ram[2382] = {9'd16,10'd216};
ram[2383] = {9'd19,10'd219};
ram[2384] = {9'd22,10'd223};
ram[2385] = {9'd25,10'd226};
ram[2386] = {9'd29,10'd229};
ram[2387] = {9'd32,10'd232};
ram[2388] = {9'd35,10'd235};
ram[2389] = {9'd38,10'd238};
ram[2390] = {9'd41,10'd241};
ram[2391] = {9'd44,10'd245};
ram[2392] = {9'd47,10'd248};
ram[2393] = {9'd51,10'd251};
ram[2394] = {9'd54,10'd254};
ram[2395] = {9'd57,10'd257};
ram[2396] = {9'd60,10'd260};
ram[2397] = {9'd63,10'd263};
ram[2398] = {9'd66,10'd267};
ram[2399] = {9'd69,10'd270};
ram[2400] = {9'd73,10'd273};
ram[2401] = {9'd76,10'd276};
ram[2402] = {9'd79,10'd279};
ram[2403] = {9'd82,10'd282};
ram[2404] = {9'd85,10'd285};
ram[2405] = {9'd88,10'd289};
ram[2406] = {9'd91,10'd292};
ram[2407] = {9'd95,10'd295};
ram[2408] = {9'd98,10'd298};
ram[2409] = {-9'd99,10'd301};
ram[2410] = {-9'd96,10'd304};
ram[2411] = {-9'd93,10'd307};
ram[2412] = {-9'd90,10'd311};
ram[2413] = {-9'd87,10'd314};
ram[2414] = {-9'd84,10'd317};
ram[2415] = {-9'd81,10'd320};
ram[2416] = {-9'd77,10'd323};
ram[2417] = {-9'd74,10'd326};
ram[2418] = {-9'd71,10'd329};
ram[2419] = {-9'd68,10'd333};
ram[2420] = {-9'd65,10'd336};
ram[2421] = {-9'd62,10'd339};
ram[2422] = {-9'd59,10'd342};
ram[2423] = {-9'd55,10'd345};
ram[2424] = {-9'd52,10'd348};
ram[2425] = {-9'd49,10'd351};
ram[2426] = {-9'd46,10'd354};
ram[2427] = {-9'd43,10'd358};
ram[2428] = {-9'd40,10'd361};
ram[2429] = {-9'd37,10'd364};
ram[2430] = {-9'd33,10'd367};
ram[2431] = {-9'd30,10'd370};
ram[2432] = {-9'd30,10'd370};
ram[2433] = {-9'd27,10'd373};
ram[2434] = {-9'd24,10'd376};
ram[2435] = {-9'd21,10'd380};
ram[2436] = {-9'd18,10'd383};
ram[2437] = {-9'd15,10'd386};
ram[2438] = {-9'd11,10'd389};
ram[2439] = {-9'd8,10'd392};
ram[2440] = {-9'd5,10'd395};
ram[2441] = {-9'd2,10'd398};
ram[2442] = {9'd1,-10'd399};
ram[2443] = {9'd4,-10'd396};
ram[2444] = {9'd7,-10'd393};
ram[2445] = {9'd10,-10'd390};
ram[2446] = {9'd14,-10'd387};
ram[2447] = {9'd17,-10'd384};
ram[2448] = {9'd20,-10'd381};
ram[2449] = {9'd23,-10'd377};
ram[2450] = {9'd26,-10'd374};
ram[2451] = {9'd29,-10'd371};
ram[2452] = {9'd32,-10'd368};
ram[2453] = {9'd36,-10'd365};
ram[2454] = {9'd39,-10'd362};
ram[2455] = {9'd42,-10'd359};
ram[2456] = {9'd45,-10'd355};
ram[2457] = {9'd48,-10'd352};
ram[2458] = {9'd51,-10'd349};
ram[2459] = {9'd54,-10'd346};
ram[2460] = {9'd58,-10'd343};
ram[2461] = {9'd61,-10'd340};
ram[2462] = {9'd64,-10'd337};
ram[2463] = {9'd67,-10'd334};
ram[2464] = {9'd70,-10'd330};
ram[2465] = {9'd73,-10'd327};
ram[2466] = {9'd76,-10'd324};
ram[2467] = {9'd80,-10'd321};
ram[2468] = {9'd83,-10'd318};
ram[2469] = {9'd86,-10'd315};
ram[2470] = {9'd89,-10'd312};
ram[2471] = {9'd92,-10'd308};
ram[2472] = {9'd95,-10'd305};
ram[2473] = {9'd98,-10'd302};
ram[2474] = {-9'd99,-10'd299};
ram[2475] = {-9'd96,-10'd296};
ram[2476] = {-9'd92,-10'd293};
ram[2477] = {-9'd89,-10'd290};
ram[2478] = {-9'd86,-10'd286};
ram[2479] = {-9'd83,-10'd283};
ram[2480] = {-9'd80,-10'd280};
ram[2481] = {-9'd77,-10'd277};
ram[2482] = {-9'd74,-10'd274};
ram[2483] = {-9'd70,-10'd271};
ram[2484] = {-9'd67,-10'd268};
ram[2485] = {-9'd64,-10'd264};
ram[2486] = {-9'd61,-10'd261};
ram[2487] = {-9'd58,-10'd258};
ram[2488] = {-9'd55,-10'd255};
ram[2489] = {-9'd52,-10'd252};
ram[2490] = {-9'd48,-10'd249};
ram[2491] = {-9'd45,-10'd246};
ram[2492] = {-9'd42,-10'd242};
ram[2493] = {-9'd39,-10'd239};
ram[2494] = {-9'd36,-10'd236};
ram[2495] = {-9'd33,-10'd233};
ram[2496] = {-9'd30,-10'd230};
ram[2497] = {-9'd26,-10'd227};
ram[2498] = {-9'd23,-10'd224};
ram[2499] = {-9'd20,-10'd220};
ram[2500] = {-9'd17,-10'd217};
ram[2501] = {-9'd14,-10'd214};
ram[2502] = {-9'd11,-10'd211};
ram[2503] = {-9'd8,-10'd208};
ram[2504] = {-9'd4,-10'd205};
ram[2505] = {-9'd1,-10'd202};
ram[2506] = {9'd2,-10'd198};
ram[2507] = {9'd5,-10'd195};
ram[2508] = {9'd8,-10'd192};
ram[2509] = {9'd11,-10'd189};
ram[2510] = {9'd14,-10'd186};
ram[2511] = {9'd18,-10'd183};
ram[2512] = {9'd21,-10'd180};
ram[2513] = {9'd24,-10'd176};
ram[2514] = {9'd27,-10'd173};
ram[2515] = {9'd30,-10'd170};
ram[2516] = {9'd33,-10'd167};
ram[2517] = {9'd36,-10'd164};
ram[2518] = {9'd40,-10'd161};
ram[2519] = {9'd43,-10'd158};
ram[2520] = {9'd46,-10'd154};
ram[2521] = {9'd49,-10'd151};
ram[2522] = {9'd52,-10'd148};
ram[2523] = {9'd55,-10'd145};
ram[2524] = {9'd58,-10'd142};
ram[2525] = {9'd62,-10'd139};
ram[2526] = {9'd65,-10'd136};
ram[2527] = {9'd68,-10'd132};
ram[2528] = {9'd71,-10'd129};
ram[2529] = {9'd74,-10'd126};
ram[2530] = {9'd77,-10'd123};
ram[2531] = {9'd80,-10'd120};
ram[2532] = {9'd84,-10'd117};
ram[2533] = {9'd87,-10'd114};
ram[2534] = {9'd90,-10'd110};
ram[2535] = {9'd93,-10'd107};
ram[2536] = {9'd96,-10'd104};
ram[2537] = {9'd99,-10'd101};
ram[2538] = {-9'd98,-10'd98};
ram[2539] = {-9'd95,-10'd95};
ram[2540] = {-9'd92,-10'd92};
ram[2541] = {-9'd88,-10'd88};
ram[2542] = {-9'd85,-10'd85};
ram[2543] = {-9'd82,-10'd82};
ram[2544] = {-9'd79,-10'd79};
ram[2545] = {-9'd76,-10'd76};
ram[2546] = {-9'd73,-10'd73};
ram[2547] = {-9'd70,-10'd70};
ram[2548] = {-9'd66,-10'd66};
ram[2549] = {-9'd63,-10'd63};
ram[2550] = {-9'd60,-10'd60};
ram[2551] = {-9'd57,-10'd57};
ram[2552] = {-9'd54,-10'd54};
ram[2553] = {-9'd51,-10'd51};
ram[2554] = {-9'd48,-10'd48};
ram[2555] = {-9'd44,-10'd44};
ram[2556] = {-9'd41,-10'd41};
ram[2557] = {-9'd38,-10'd38};
ram[2558] = {-9'd35,-10'd35};
ram[2559] = {-9'd32,-10'd32};
ram[2560] = {-9'd32,-10'd32};
ram[2561] = {-9'd29,-10'd29};
ram[2562] = {-9'd26,-10'd26};
ram[2563] = {-9'd22,-10'd22};
ram[2564] = {-9'd19,-10'd19};
ram[2565] = {-9'd16,-10'd16};
ram[2566] = {-9'd13,-10'd13};
ram[2567] = {-9'd10,-10'd10};
ram[2568] = {-9'd7,-10'd7};
ram[2569] = {-9'd4,-10'd4};
ram[2570] = {9'd0,10'd0};
ram[2571] = {9'd3,10'd3};
ram[2572] = {9'd6,10'd6};
ram[2573] = {9'd9,10'd9};
ram[2574] = {9'd12,10'd12};
ram[2575] = {9'd15,10'd15};
ram[2576] = {9'd18,10'd18};
ram[2577] = {9'd21,10'd21};
ram[2578] = {9'd25,10'd25};
ram[2579] = {9'd28,10'd28};
ram[2580] = {9'd31,10'd31};
ram[2581] = {9'd34,10'd34};
ram[2582] = {9'd37,10'd37};
ram[2583] = {9'd40,10'd40};
ram[2584] = {9'd43,10'd43};
ram[2585] = {9'd47,10'd47};
ram[2586] = {9'd50,10'd50};
ram[2587] = {9'd53,10'd53};
ram[2588] = {9'd56,10'd56};
ram[2589] = {9'd59,10'd59};
ram[2590] = {9'd62,10'd62};
ram[2591] = {9'd65,10'd65};
ram[2592] = {9'd69,10'd69};
ram[2593] = {9'd72,10'd72};
ram[2594] = {9'd75,10'd75};
ram[2595] = {9'd78,10'd78};
ram[2596] = {9'd81,10'd81};
ram[2597] = {9'd84,10'd84};
ram[2598] = {9'd87,10'd87};
ram[2599] = {9'd91,10'd91};
ram[2600] = {9'd94,10'd94};
ram[2601] = {9'd97,10'd97};
ram[2602] = {-9'd100,10'd100};
ram[2603] = {-9'd97,10'd103};
ram[2604] = {-9'd94,10'd106};
ram[2605] = {-9'd91,10'd109};
ram[2606] = {-9'd88,10'd113};
ram[2607] = {-9'd85,10'd116};
ram[2608] = {-9'd81,10'd119};
ram[2609] = {-9'd78,10'd122};
ram[2610] = {-9'd75,10'd125};
ram[2611] = {-9'd72,10'd128};
ram[2612] = {-9'd69,10'd131};
ram[2613] = {-9'd66,10'd135};
ram[2614] = {-9'd63,10'd138};
ram[2615] = {-9'd59,10'd141};
ram[2616] = {-9'd56,10'd144};
ram[2617] = {-9'd53,10'd147};
ram[2618] = {-9'd50,10'd150};
ram[2619] = {-9'd47,10'd153};
ram[2620] = {-9'd44,10'd157};
ram[2621] = {-9'd41,10'd160};
ram[2622] = {-9'd37,10'd163};
ram[2623] = {-9'd34,10'd166};
ram[2624] = {-9'd31,10'd169};
ram[2625] = {-9'd28,10'd172};
ram[2626] = {-9'd25,10'd175};
ram[2627] = {-9'd22,10'd179};
ram[2628] = {-9'd19,10'd182};
ram[2629] = {-9'd15,10'd185};
ram[2630] = {-9'd12,10'd188};
ram[2631] = {-9'd9,10'd191};
ram[2632] = {-9'd6,10'd194};
ram[2633] = {-9'd3,10'd197};
ram[2634] = {9'd0,10'd201};
ram[2635] = {9'd3,10'd204};
ram[2636] = {9'd7,10'd207};
ram[2637] = {9'd10,10'd210};
ram[2638] = {9'd13,10'd213};
ram[2639] = {9'd16,10'd216};
ram[2640] = {9'd19,10'd219};
ram[2641] = {9'd22,10'd223};
ram[2642] = {9'd25,10'd226};
ram[2643] = {9'd29,10'd229};
ram[2644] = {9'd32,10'd232};
ram[2645] = {9'd35,10'd235};
ram[2646] = {9'd38,10'd238};
ram[2647] = {9'd41,10'd241};
ram[2648] = {9'd44,10'd245};
ram[2649] = {9'd47,10'd248};
ram[2650] = {9'd51,10'd251};
ram[2651] = {9'd54,10'd254};
ram[2652] = {9'd57,10'd257};
ram[2653] = {9'd60,10'd260};
ram[2654] = {9'd63,10'd263};
ram[2655] = {9'd66,10'd267};
ram[2656] = {9'd69,10'd270};
ram[2657] = {9'd73,10'd273};
ram[2658] = {9'd76,10'd276};
ram[2659] = {9'd79,10'd279};
ram[2660] = {9'd82,10'd282};
ram[2661] = {9'd85,10'd285};
ram[2662] = {9'd88,10'd289};
ram[2663] = {9'd91,10'd292};
ram[2664] = {9'd95,10'd295};
ram[2665] = {9'd98,10'd298};
ram[2666] = {-9'd99,10'd301};
ram[2667] = {-9'd96,10'd304};
ram[2668] = {-9'd93,10'd307};
ram[2669] = {-9'd90,10'd311};
ram[2670] = {-9'd87,10'd314};
ram[2671] = {-9'd84,10'd317};
ram[2672] = {-9'd81,10'd320};
ram[2673] = {-9'd77,10'd323};
ram[2674] = {-9'd74,10'd326};
ram[2675] = {-9'd71,10'd329};
ram[2676] = {-9'd68,10'd333};
ram[2677] = {-9'd65,10'd336};
ram[2678] = {-9'd62,10'd339};
ram[2679] = {-9'd59,10'd342};
ram[2680] = {-9'd55,10'd345};
ram[2681] = {-9'd52,10'd348};
ram[2682] = {-9'd49,10'd351};
ram[2683] = {-9'd46,10'd354};
ram[2684] = {-9'd43,10'd358};
ram[2685] = {-9'd40,10'd361};
ram[2686] = {-9'd37,10'd364};
ram[2687] = {-9'd33,10'd367};
ram[2688] = {-9'd33,10'd367};
ram[2689] = {-9'd30,10'd370};
ram[2690] = {-9'd27,10'd373};
ram[2691] = {-9'd24,10'd376};
ram[2692] = {-9'd21,10'd380};
ram[2693] = {-9'd18,10'd383};
ram[2694] = {-9'd15,10'd386};
ram[2695] = {-9'd11,10'd389};
ram[2696] = {-9'd8,10'd392};
ram[2697] = {-9'd5,10'd395};
ram[2698] = {-9'd2,10'd398};
ram[2699] = {9'd1,-10'd399};
ram[2700] = {9'd4,-10'd396};
ram[2701] = {9'd7,-10'd393};
ram[2702] = {9'd10,-10'd390};
ram[2703] = {9'd14,-10'd387};
ram[2704] = {9'd17,-10'd384};
ram[2705] = {9'd20,-10'd381};
ram[2706] = {9'd23,-10'd377};
ram[2707] = {9'd26,-10'd374};
ram[2708] = {9'd29,-10'd371};
ram[2709] = {9'd32,-10'd368};
ram[2710] = {9'd36,-10'd365};
ram[2711] = {9'd39,-10'd362};
ram[2712] = {9'd42,-10'd359};
ram[2713] = {9'd45,-10'd355};
ram[2714] = {9'd48,-10'd352};
ram[2715] = {9'd51,-10'd349};
ram[2716] = {9'd54,-10'd346};
ram[2717] = {9'd58,-10'd343};
ram[2718] = {9'd61,-10'd340};
ram[2719] = {9'd64,-10'd337};
ram[2720] = {9'd67,-10'd334};
ram[2721] = {9'd70,-10'd330};
ram[2722] = {9'd73,-10'd327};
ram[2723] = {9'd76,-10'd324};
ram[2724] = {9'd80,-10'd321};
ram[2725] = {9'd83,-10'd318};
ram[2726] = {9'd86,-10'd315};
ram[2727] = {9'd89,-10'd312};
ram[2728] = {9'd92,-10'd308};
ram[2729] = {9'd95,-10'd305};
ram[2730] = {9'd98,-10'd302};
ram[2731] = {-9'd99,-10'd299};
ram[2732] = {-9'd96,-10'd296};
ram[2733] = {-9'd92,-10'd293};
ram[2734] = {-9'd89,-10'd290};
ram[2735] = {-9'd86,-10'd286};
ram[2736] = {-9'd83,-10'd283};
ram[2737] = {-9'd80,-10'd280};
ram[2738] = {-9'd77,-10'd277};
ram[2739] = {-9'd74,-10'd274};
ram[2740] = {-9'd70,-10'd271};
ram[2741] = {-9'd67,-10'd268};
ram[2742] = {-9'd64,-10'd264};
ram[2743] = {-9'd61,-10'd261};
ram[2744] = {-9'd58,-10'd258};
ram[2745] = {-9'd55,-10'd255};
ram[2746] = {-9'd52,-10'd252};
ram[2747] = {-9'd48,-10'd249};
ram[2748] = {-9'd45,-10'd246};
ram[2749] = {-9'd42,-10'd242};
ram[2750] = {-9'd39,-10'd239};
ram[2751] = {-9'd36,-10'd236};
ram[2752] = {-9'd33,-10'd233};
ram[2753] = {-9'd30,-10'd230};
ram[2754] = {-9'd26,-10'd227};
ram[2755] = {-9'd23,-10'd224};
ram[2756] = {-9'd20,-10'd220};
ram[2757] = {-9'd17,-10'd217};
ram[2758] = {-9'd14,-10'd214};
ram[2759] = {-9'd11,-10'd211};
ram[2760] = {-9'd8,-10'd208};
ram[2761] = {-9'd4,-10'd205};
ram[2762] = {-9'd1,-10'd202};
ram[2763] = {9'd2,-10'd198};
ram[2764] = {9'd5,-10'd195};
ram[2765] = {9'd8,-10'd192};
ram[2766] = {9'd11,-10'd189};
ram[2767] = {9'd14,-10'd186};
ram[2768] = {9'd18,-10'd183};
ram[2769] = {9'd21,-10'd180};
ram[2770] = {9'd24,-10'd176};
ram[2771] = {9'd27,-10'd173};
ram[2772] = {9'd30,-10'd170};
ram[2773] = {9'd33,-10'd167};
ram[2774] = {9'd36,-10'd164};
ram[2775] = {9'd40,-10'd161};
ram[2776] = {9'd43,-10'd158};
ram[2777] = {9'd46,-10'd154};
ram[2778] = {9'd49,-10'd151};
ram[2779] = {9'd52,-10'd148};
ram[2780] = {9'd55,-10'd145};
ram[2781] = {9'd58,-10'd142};
ram[2782] = {9'd62,-10'd139};
ram[2783] = {9'd65,-10'd136};
ram[2784] = {9'd68,-10'd132};
ram[2785] = {9'd71,-10'd129};
ram[2786] = {9'd74,-10'd126};
ram[2787] = {9'd77,-10'd123};
ram[2788] = {9'd80,-10'd120};
ram[2789] = {9'd84,-10'd117};
ram[2790] = {9'd87,-10'd114};
ram[2791] = {9'd90,-10'd110};
ram[2792] = {9'd93,-10'd107};
ram[2793] = {9'd96,-10'd104};
ram[2794] = {9'd99,-10'd101};
ram[2795] = {-9'd98,-10'd98};
ram[2796] = {-9'd95,-10'd95};
ram[2797] = {-9'd92,-10'd92};
ram[2798] = {-9'd88,-10'd88};
ram[2799] = {-9'd85,-10'd85};
ram[2800] = {-9'd82,-10'd82};
ram[2801] = {-9'd79,-10'd79};
ram[2802] = {-9'd76,-10'd76};
ram[2803] = {-9'd73,-10'd73};
ram[2804] = {-9'd70,-10'd70};
ram[2805] = {-9'd66,-10'd66};
ram[2806] = {-9'd63,-10'd63};
ram[2807] = {-9'd60,-10'd60};
ram[2808] = {-9'd57,-10'd57};
ram[2809] = {-9'd54,-10'd54};
ram[2810] = {-9'd51,-10'd51};
ram[2811] = {-9'd48,-10'd48};
ram[2812] = {-9'd44,-10'd44};
ram[2813] = {-9'd41,-10'd41};
ram[2814] = {-9'd38,-10'd38};
ram[2815] = {-9'd35,-10'd35};
ram[2816] = {-9'd35,-10'd35};
ram[2817] = {-9'd32,-10'd32};
ram[2818] = {-9'd29,-10'd29};
ram[2819] = {-9'd26,-10'd26};
ram[2820] = {-9'd22,-10'd22};
ram[2821] = {-9'd19,-10'd19};
ram[2822] = {-9'd16,-10'd16};
ram[2823] = {-9'd13,-10'd13};
ram[2824] = {-9'd10,-10'd10};
ram[2825] = {-9'd7,-10'd7};
ram[2826] = {-9'd4,-10'd4};
ram[2827] = {9'd0,10'd0};
ram[2828] = {9'd3,10'd3};
ram[2829] = {9'd6,10'd6};
ram[2830] = {9'd9,10'd9};
ram[2831] = {9'd12,10'd12};
ram[2832] = {9'd15,10'd15};
ram[2833] = {9'd18,10'd18};
ram[2834] = {9'd21,10'd21};
ram[2835] = {9'd25,10'd25};
ram[2836] = {9'd28,10'd28};
ram[2837] = {9'd31,10'd31};
ram[2838] = {9'd34,10'd34};
ram[2839] = {9'd37,10'd37};
ram[2840] = {9'd40,10'd40};
ram[2841] = {9'd43,10'd43};
ram[2842] = {9'd47,10'd47};
ram[2843] = {9'd50,10'd50};
ram[2844] = {9'd53,10'd53};
ram[2845] = {9'd56,10'd56};
ram[2846] = {9'd59,10'd59};
ram[2847] = {9'd62,10'd62};
ram[2848] = {9'd65,10'd65};
ram[2849] = {9'd69,10'd69};
ram[2850] = {9'd72,10'd72};
ram[2851] = {9'd75,10'd75};
ram[2852] = {9'd78,10'd78};
ram[2853] = {9'd81,10'd81};
ram[2854] = {9'd84,10'd84};
ram[2855] = {9'd87,10'd87};
ram[2856] = {9'd91,10'd91};
ram[2857] = {9'd94,10'd94};
ram[2858] = {9'd97,10'd97};
ram[2859] = {-9'd100,10'd100};
ram[2860] = {-9'd97,10'd103};
ram[2861] = {-9'd94,10'd106};
ram[2862] = {-9'd91,10'd109};
ram[2863] = {-9'd88,10'd113};
ram[2864] = {-9'd85,10'd116};
ram[2865] = {-9'd81,10'd119};
ram[2866] = {-9'd78,10'd122};
ram[2867] = {-9'd75,10'd125};
ram[2868] = {-9'd72,10'd128};
ram[2869] = {-9'd69,10'd131};
ram[2870] = {-9'd66,10'd135};
ram[2871] = {-9'd63,10'd138};
ram[2872] = {-9'd59,10'd141};
ram[2873] = {-9'd56,10'd144};
ram[2874] = {-9'd53,10'd147};
ram[2875] = {-9'd50,10'd150};
ram[2876] = {-9'd47,10'd153};
ram[2877] = {-9'd44,10'd157};
ram[2878] = {-9'd41,10'd160};
ram[2879] = {-9'd37,10'd163};
ram[2880] = {-9'd34,10'd166};
ram[2881] = {-9'd31,10'd169};
ram[2882] = {-9'd28,10'd172};
ram[2883] = {-9'd25,10'd175};
ram[2884] = {-9'd22,10'd179};
ram[2885] = {-9'd19,10'd182};
ram[2886] = {-9'd15,10'd185};
ram[2887] = {-9'd12,10'd188};
ram[2888] = {-9'd9,10'd191};
ram[2889] = {-9'd6,10'd194};
ram[2890] = {-9'd3,10'd197};
ram[2891] = {9'd0,10'd201};
ram[2892] = {9'd3,10'd204};
ram[2893] = {9'd7,10'd207};
ram[2894] = {9'd10,10'd210};
ram[2895] = {9'd13,10'd213};
ram[2896] = {9'd16,10'd216};
ram[2897] = {9'd19,10'd219};
ram[2898] = {9'd22,10'd223};
ram[2899] = {9'd25,10'd226};
ram[2900] = {9'd29,10'd229};
ram[2901] = {9'd32,10'd232};
ram[2902] = {9'd35,10'd235};
ram[2903] = {9'd38,10'd238};
ram[2904] = {9'd41,10'd241};
ram[2905] = {9'd44,10'd245};
ram[2906] = {9'd47,10'd248};
ram[2907] = {9'd51,10'd251};
ram[2908] = {9'd54,10'd254};
ram[2909] = {9'd57,10'd257};
ram[2910] = {9'd60,10'd260};
ram[2911] = {9'd63,10'd263};
ram[2912] = {9'd66,10'd267};
ram[2913] = {9'd69,10'd270};
ram[2914] = {9'd73,10'd273};
ram[2915] = {9'd76,10'd276};
ram[2916] = {9'd79,10'd279};
ram[2917] = {9'd82,10'd282};
ram[2918] = {9'd85,10'd285};
ram[2919] = {9'd88,10'd289};
ram[2920] = {9'd91,10'd292};
ram[2921] = {9'd95,10'd295};
ram[2922] = {9'd98,10'd298};
ram[2923] = {-9'd99,10'd301};
ram[2924] = {-9'd96,10'd304};
ram[2925] = {-9'd93,10'd307};
ram[2926] = {-9'd90,10'd311};
ram[2927] = {-9'd87,10'd314};
ram[2928] = {-9'd84,10'd317};
ram[2929] = {-9'd81,10'd320};
ram[2930] = {-9'd77,10'd323};
ram[2931] = {-9'd74,10'd326};
ram[2932] = {-9'd71,10'd329};
ram[2933] = {-9'd68,10'd333};
ram[2934] = {-9'd65,10'd336};
ram[2935] = {-9'd62,10'd339};
ram[2936] = {-9'd59,10'd342};
ram[2937] = {-9'd55,10'd345};
ram[2938] = {-9'd52,10'd348};
ram[2939] = {-9'd49,10'd351};
ram[2940] = {-9'd46,10'd354};
ram[2941] = {-9'd43,10'd358};
ram[2942] = {-9'd40,10'd361};
ram[2943] = {-9'd37,10'd364};
ram[2944] = {-9'd37,10'd364};
ram[2945] = {-9'd33,10'd367};
ram[2946] = {-9'd30,10'd370};
ram[2947] = {-9'd27,10'd373};
ram[2948] = {-9'd24,10'd376};
ram[2949] = {-9'd21,10'd380};
ram[2950] = {-9'd18,10'd383};
ram[2951] = {-9'd15,10'd386};
ram[2952] = {-9'd11,10'd389};
ram[2953] = {-9'd8,10'd392};
ram[2954] = {-9'd5,10'd395};
ram[2955] = {-9'd2,10'd398};
ram[2956] = {9'd1,-10'd399};
ram[2957] = {9'd4,-10'd396};
ram[2958] = {9'd7,-10'd393};
ram[2959] = {9'd10,-10'd390};
ram[2960] = {9'd14,-10'd387};
ram[2961] = {9'd17,-10'd384};
ram[2962] = {9'd20,-10'd381};
ram[2963] = {9'd23,-10'd377};
ram[2964] = {9'd26,-10'd374};
ram[2965] = {9'd29,-10'd371};
ram[2966] = {9'd32,-10'd368};
ram[2967] = {9'd36,-10'd365};
ram[2968] = {9'd39,-10'd362};
ram[2969] = {9'd42,-10'd359};
ram[2970] = {9'd45,-10'd355};
ram[2971] = {9'd48,-10'd352};
ram[2972] = {9'd51,-10'd349};
ram[2973] = {9'd54,-10'd346};
ram[2974] = {9'd58,-10'd343};
ram[2975] = {9'd61,-10'd340};
ram[2976] = {9'd64,-10'd337};
ram[2977] = {9'd67,-10'd334};
ram[2978] = {9'd70,-10'd330};
ram[2979] = {9'd73,-10'd327};
ram[2980] = {9'd76,-10'd324};
ram[2981] = {9'd80,-10'd321};
ram[2982] = {9'd83,-10'd318};
ram[2983] = {9'd86,-10'd315};
ram[2984] = {9'd89,-10'd312};
ram[2985] = {9'd92,-10'd308};
ram[2986] = {9'd95,-10'd305};
ram[2987] = {9'd98,-10'd302};
ram[2988] = {-9'd99,-10'd299};
ram[2989] = {-9'd96,-10'd296};
ram[2990] = {-9'd92,-10'd293};
ram[2991] = {-9'd89,-10'd290};
ram[2992] = {-9'd86,-10'd286};
ram[2993] = {-9'd83,-10'd283};
ram[2994] = {-9'd80,-10'd280};
ram[2995] = {-9'd77,-10'd277};
ram[2996] = {-9'd74,-10'd274};
ram[2997] = {-9'd70,-10'd271};
ram[2998] = {-9'd67,-10'd268};
ram[2999] = {-9'd64,-10'd264};
ram[3000] = {-9'd61,-10'd261};
ram[3001] = {-9'd58,-10'd258};
ram[3002] = {-9'd55,-10'd255};
ram[3003] = {-9'd52,-10'd252};
ram[3004] = {-9'd48,-10'd249};
ram[3005] = {-9'd45,-10'd246};
ram[3006] = {-9'd42,-10'd242};
ram[3007] = {-9'd39,-10'd239};
ram[3008] = {-9'd36,-10'd236};
ram[3009] = {-9'd33,-10'd233};
ram[3010] = {-9'd30,-10'd230};
ram[3011] = {-9'd26,-10'd227};
ram[3012] = {-9'd23,-10'd224};
ram[3013] = {-9'd20,-10'd220};
ram[3014] = {-9'd17,-10'd217};
ram[3015] = {-9'd14,-10'd214};
ram[3016] = {-9'd11,-10'd211};
ram[3017] = {-9'd8,-10'd208};
ram[3018] = {-9'd4,-10'd205};
ram[3019] = {-9'd1,-10'd202};
ram[3020] = {9'd2,-10'd198};
ram[3021] = {9'd5,-10'd195};
ram[3022] = {9'd8,-10'd192};
ram[3023] = {9'd11,-10'd189};
ram[3024] = {9'd14,-10'd186};
ram[3025] = {9'd18,-10'd183};
ram[3026] = {9'd21,-10'd180};
ram[3027] = {9'd24,-10'd176};
ram[3028] = {9'd27,-10'd173};
ram[3029] = {9'd30,-10'd170};
ram[3030] = {9'd33,-10'd167};
ram[3031] = {9'd36,-10'd164};
ram[3032] = {9'd40,-10'd161};
ram[3033] = {9'd43,-10'd158};
ram[3034] = {9'd46,-10'd154};
ram[3035] = {9'd49,-10'd151};
ram[3036] = {9'd52,-10'd148};
ram[3037] = {9'd55,-10'd145};
ram[3038] = {9'd58,-10'd142};
ram[3039] = {9'd62,-10'd139};
ram[3040] = {9'd65,-10'd136};
ram[3041] = {9'd68,-10'd132};
ram[3042] = {9'd71,-10'd129};
ram[3043] = {9'd74,-10'd126};
ram[3044] = {9'd77,-10'd123};
ram[3045] = {9'd80,-10'd120};
ram[3046] = {9'd84,-10'd117};
ram[3047] = {9'd87,-10'd114};
ram[3048] = {9'd90,-10'd110};
ram[3049] = {9'd93,-10'd107};
ram[3050] = {9'd96,-10'd104};
ram[3051] = {9'd99,-10'd101};
ram[3052] = {-9'd98,-10'd98};
ram[3053] = {-9'd95,-10'd95};
ram[3054] = {-9'd92,-10'd92};
ram[3055] = {-9'd88,-10'd88};
ram[3056] = {-9'd85,-10'd85};
ram[3057] = {-9'd82,-10'd82};
ram[3058] = {-9'd79,-10'd79};
ram[3059] = {-9'd76,-10'd76};
ram[3060] = {-9'd73,-10'd73};
ram[3061] = {-9'd70,-10'd70};
ram[3062] = {-9'd66,-10'd66};
ram[3063] = {-9'd63,-10'd63};
ram[3064] = {-9'd60,-10'd60};
ram[3065] = {-9'd57,-10'd57};
ram[3066] = {-9'd54,-10'd54};
ram[3067] = {-9'd51,-10'd51};
ram[3068] = {-9'd48,-10'd48};
ram[3069] = {-9'd44,-10'd44};
ram[3070] = {-9'd41,-10'd41};
ram[3071] = {-9'd38,-10'd38};
ram[3072] = {-9'd38,-10'd38};
ram[3073] = {-9'd35,-10'd35};
ram[3074] = {-9'd32,-10'd32};
ram[3075] = {-9'd29,-10'd29};
ram[3076] = {-9'd26,-10'd26};
ram[3077] = {-9'd22,-10'd22};
ram[3078] = {-9'd19,-10'd19};
ram[3079] = {-9'd16,-10'd16};
ram[3080] = {-9'd13,-10'd13};
ram[3081] = {-9'd10,-10'd10};
ram[3082] = {-9'd7,-10'd7};
ram[3083] = {-9'd4,-10'd4};
ram[3084] = {9'd0,10'd0};
ram[3085] = {9'd3,10'd3};
ram[3086] = {9'd6,10'd6};
ram[3087] = {9'd9,10'd9};
ram[3088] = {9'd12,10'd12};
ram[3089] = {9'd15,10'd15};
ram[3090] = {9'd18,10'd18};
ram[3091] = {9'd21,10'd21};
ram[3092] = {9'd25,10'd25};
ram[3093] = {9'd28,10'd28};
ram[3094] = {9'd31,10'd31};
ram[3095] = {9'd34,10'd34};
ram[3096] = {9'd37,10'd37};
ram[3097] = {9'd40,10'd40};
ram[3098] = {9'd43,10'd43};
ram[3099] = {9'd47,10'd47};
ram[3100] = {9'd50,10'd50};
ram[3101] = {9'd53,10'd53};
ram[3102] = {9'd56,10'd56};
ram[3103] = {9'd59,10'd59};
ram[3104] = {9'd62,10'd62};
ram[3105] = {9'd65,10'd65};
ram[3106] = {9'd69,10'd69};
ram[3107] = {9'd72,10'd72};
ram[3108] = {9'd75,10'd75};
ram[3109] = {9'd78,10'd78};
ram[3110] = {9'd81,10'd81};
ram[3111] = {9'd84,10'd84};
ram[3112] = {9'd87,10'd87};
ram[3113] = {9'd91,10'd91};
ram[3114] = {9'd94,10'd94};
ram[3115] = {9'd97,10'd97};
ram[3116] = {-9'd100,10'd100};
ram[3117] = {-9'd97,10'd103};
ram[3118] = {-9'd94,10'd106};
ram[3119] = {-9'd91,10'd109};
ram[3120] = {-9'd88,10'd113};
ram[3121] = {-9'd85,10'd116};
ram[3122] = {-9'd81,10'd119};
ram[3123] = {-9'd78,10'd122};
ram[3124] = {-9'd75,10'd125};
ram[3125] = {-9'd72,10'd128};
ram[3126] = {-9'd69,10'd131};
ram[3127] = {-9'd66,10'd135};
ram[3128] = {-9'd63,10'd138};
ram[3129] = {-9'd59,10'd141};
ram[3130] = {-9'd56,10'd144};
ram[3131] = {-9'd53,10'd147};
ram[3132] = {-9'd50,10'd150};
ram[3133] = {-9'd47,10'd153};
ram[3134] = {-9'd44,10'd157};
ram[3135] = {-9'd41,10'd160};
ram[3136] = {-9'd37,10'd163};
ram[3137] = {-9'd34,10'd166};
ram[3138] = {-9'd31,10'd169};
ram[3139] = {-9'd28,10'd172};
ram[3140] = {-9'd25,10'd175};
ram[3141] = {-9'd22,10'd179};
ram[3142] = {-9'd19,10'd182};
ram[3143] = {-9'd15,10'd185};
ram[3144] = {-9'd12,10'd188};
ram[3145] = {-9'd9,10'd191};
ram[3146] = {-9'd6,10'd194};
ram[3147] = {-9'd3,10'd197};
ram[3148] = {9'd0,10'd201};
ram[3149] = {9'd3,10'd204};
ram[3150] = {9'd7,10'd207};
ram[3151] = {9'd10,10'd210};
ram[3152] = {9'd13,10'd213};
ram[3153] = {9'd16,10'd216};
ram[3154] = {9'd19,10'd219};
ram[3155] = {9'd22,10'd223};
ram[3156] = {9'd25,10'd226};
ram[3157] = {9'd29,10'd229};
ram[3158] = {9'd32,10'd232};
ram[3159] = {9'd35,10'd235};
ram[3160] = {9'd38,10'd238};
ram[3161] = {9'd41,10'd241};
ram[3162] = {9'd44,10'd245};
ram[3163] = {9'd47,10'd248};
ram[3164] = {9'd51,10'd251};
ram[3165] = {9'd54,10'd254};
ram[3166] = {9'd57,10'd257};
ram[3167] = {9'd60,10'd260};
ram[3168] = {9'd63,10'd263};
ram[3169] = {9'd66,10'd267};
ram[3170] = {9'd69,10'd270};
ram[3171] = {9'd73,10'd273};
ram[3172] = {9'd76,10'd276};
ram[3173] = {9'd79,10'd279};
ram[3174] = {9'd82,10'd282};
ram[3175] = {9'd85,10'd285};
ram[3176] = {9'd88,10'd289};
ram[3177] = {9'd91,10'd292};
ram[3178] = {9'd95,10'd295};
ram[3179] = {9'd98,10'd298};
ram[3180] = {-9'd99,10'd301};
ram[3181] = {-9'd96,10'd304};
ram[3182] = {-9'd93,10'd307};
ram[3183] = {-9'd90,10'd311};
ram[3184] = {-9'd87,10'd314};
ram[3185] = {-9'd84,10'd317};
ram[3186] = {-9'd81,10'd320};
ram[3187] = {-9'd77,10'd323};
ram[3188] = {-9'd74,10'd326};
ram[3189] = {-9'd71,10'd329};
ram[3190] = {-9'd68,10'd333};
ram[3191] = {-9'd65,10'd336};
ram[3192] = {-9'd62,10'd339};
ram[3193] = {-9'd59,10'd342};
ram[3194] = {-9'd55,10'd345};
ram[3195] = {-9'd52,10'd348};
ram[3196] = {-9'd49,10'd351};
ram[3197] = {-9'd46,10'd354};
ram[3198] = {-9'd43,10'd358};
ram[3199] = {-9'd40,10'd361};
ram[3200] = {-9'd40,10'd361};
ram[3201] = {-9'd37,10'd364};
ram[3202] = {-9'd33,10'd367};
ram[3203] = {-9'd30,10'd370};
ram[3204] = {-9'd27,10'd373};
ram[3205] = {-9'd24,10'd376};
ram[3206] = {-9'd21,10'd380};
ram[3207] = {-9'd18,10'd383};
ram[3208] = {-9'd15,10'd386};
ram[3209] = {-9'd11,10'd389};
ram[3210] = {-9'd8,10'd392};
ram[3211] = {-9'd5,10'd395};
ram[3212] = {-9'd2,10'd398};
ram[3213] = {9'd1,-10'd399};
ram[3214] = {9'd4,-10'd396};
ram[3215] = {9'd7,-10'd393};
ram[3216] = {9'd10,-10'd390};
ram[3217] = {9'd14,-10'd387};
ram[3218] = {9'd17,-10'd384};
ram[3219] = {9'd20,-10'd381};
ram[3220] = {9'd23,-10'd377};
ram[3221] = {9'd26,-10'd374};
ram[3222] = {9'd29,-10'd371};
ram[3223] = {9'd32,-10'd368};
ram[3224] = {9'd36,-10'd365};
ram[3225] = {9'd39,-10'd362};
ram[3226] = {9'd42,-10'd359};
ram[3227] = {9'd45,-10'd355};
ram[3228] = {9'd48,-10'd352};
ram[3229] = {9'd51,-10'd349};
ram[3230] = {9'd54,-10'd346};
ram[3231] = {9'd58,-10'd343};
ram[3232] = {9'd61,-10'd340};
ram[3233] = {9'd64,-10'd337};
ram[3234] = {9'd67,-10'd334};
ram[3235] = {9'd70,-10'd330};
ram[3236] = {9'd73,-10'd327};
ram[3237] = {9'd76,-10'd324};
ram[3238] = {9'd80,-10'd321};
ram[3239] = {9'd83,-10'd318};
ram[3240] = {9'd86,-10'd315};
ram[3241] = {9'd89,-10'd312};
ram[3242] = {9'd92,-10'd308};
ram[3243] = {9'd95,-10'd305};
ram[3244] = {9'd98,-10'd302};
ram[3245] = {-9'd99,-10'd299};
ram[3246] = {-9'd96,-10'd296};
ram[3247] = {-9'd92,-10'd293};
ram[3248] = {-9'd89,-10'd290};
ram[3249] = {-9'd86,-10'd286};
ram[3250] = {-9'd83,-10'd283};
ram[3251] = {-9'd80,-10'd280};
ram[3252] = {-9'd77,-10'd277};
ram[3253] = {-9'd74,-10'd274};
ram[3254] = {-9'd70,-10'd271};
ram[3255] = {-9'd67,-10'd268};
ram[3256] = {-9'd64,-10'd264};
ram[3257] = {-9'd61,-10'd261};
ram[3258] = {-9'd58,-10'd258};
ram[3259] = {-9'd55,-10'd255};
ram[3260] = {-9'd52,-10'd252};
ram[3261] = {-9'd48,-10'd249};
ram[3262] = {-9'd45,-10'd246};
ram[3263] = {-9'd42,-10'd242};
ram[3264] = {-9'd39,-10'd239};
ram[3265] = {-9'd36,-10'd236};
ram[3266] = {-9'd33,-10'd233};
ram[3267] = {-9'd30,-10'd230};
ram[3268] = {-9'd26,-10'd227};
ram[3269] = {-9'd23,-10'd224};
ram[3270] = {-9'd20,-10'd220};
ram[3271] = {-9'd17,-10'd217};
ram[3272] = {-9'd14,-10'd214};
ram[3273] = {-9'd11,-10'd211};
ram[3274] = {-9'd8,-10'd208};
ram[3275] = {-9'd4,-10'd205};
ram[3276] = {-9'd1,-10'd202};
ram[3277] = {9'd2,-10'd198};
ram[3278] = {9'd5,-10'd195};
ram[3279] = {9'd8,-10'd192};
ram[3280] = {9'd11,-10'd189};
ram[3281] = {9'd14,-10'd186};
ram[3282] = {9'd18,-10'd183};
ram[3283] = {9'd21,-10'd180};
ram[3284] = {9'd24,-10'd176};
ram[3285] = {9'd27,-10'd173};
ram[3286] = {9'd30,-10'd170};
ram[3287] = {9'd33,-10'd167};
ram[3288] = {9'd36,-10'd164};
ram[3289] = {9'd40,-10'd161};
ram[3290] = {9'd43,-10'd158};
ram[3291] = {9'd46,-10'd154};
ram[3292] = {9'd49,-10'd151};
ram[3293] = {9'd52,-10'd148};
ram[3294] = {9'd55,-10'd145};
ram[3295] = {9'd58,-10'd142};
ram[3296] = {9'd62,-10'd139};
ram[3297] = {9'd65,-10'd136};
ram[3298] = {9'd68,-10'd132};
ram[3299] = {9'd71,-10'd129};
ram[3300] = {9'd74,-10'd126};
ram[3301] = {9'd77,-10'd123};
ram[3302] = {9'd80,-10'd120};
ram[3303] = {9'd84,-10'd117};
ram[3304] = {9'd87,-10'd114};
ram[3305] = {9'd90,-10'd110};
ram[3306] = {9'd93,-10'd107};
ram[3307] = {9'd96,-10'd104};
ram[3308] = {9'd99,-10'd101};
ram[3309] = {-9'd98,-10'd98};
ram[3310] = {-9'd95,-10'd95};
ram[3311] = {-9'd92,-10'd92};
ram[3312] = {-9'd88,-10'd88};
ram[3313] = {-9'd85,-10'd85};
ram[3314] = {-9'd82,-10'd82};
ram[3315] = {-9'd79,-10'd79};
ram[3316] = {-9'd76,-10'd76};
ram[3317] = {-9'd73,-10'd73};
ram[3318] = {-9'd70,-10'd70};
ram[3319] = {-9'd66,-10'd66};
ram[3320] = {-9'd63,-10'd63};
ram[3321] = {-9'd60,-10'd60};
ram[3322] = {-9'd57,-10'd57};
ram[3323] = {-9'd54,-10'd54};
ram[3324] = {-9'd51,-10'd51};
ram[3325] = {-9'd48,-10'd48};
ram[3326] = {-9'd44,-10'd44};
ram[3327] = {-9'd41,-10'd41};
ram[3328] = {-9'd41,-10'd41};
ram[3329] = {-9'd38,-10'd38};
ram[3330] = {-9'd35,-10'd35};
ram[3331] = {-9'd32,-10'd32};
ram[3332] = {-9'd29,-10'd29};
ram[3333] = {-9'd26,-10'd26};
ram[3334] = {-9'd22,-10'd22};
ram[3335] = {-9'd19,-10'd19};
ram[3336] = {-9'd16,-10'd16};
ram[3337] = {-9'd13,-10'd13};
ram[3338] = {-9'd10,-10'd10};
ram[3339] = {-9'd7,-10'd7};
ram[3340] = {-9'd4,-10'd4};
ram[3341] = {9'd0,10'd0};
ram[3342] = {9'd3,10'd3};
ram[3343] = {9'd6,10'd6};
ram[3344] = {9'd9,10'd9};
ram[3345] = {9'd12,10'd12};
ram[3346] = {9'd15,10'd15};
ram[3347] = {9'd18,10'd18};
ram[3348] = {9'd21,10'd21};
ram[3349] = {9'd25,10'd25};
ram[3350] = {9'd28,10'd28};
ram[3351] = {9'd31,10'd31};
ram[3352] = {9'd34,10'd34};
ram[3353] = {9'd37,10'd37};
ram[3354] = {9'd40,10'd40};
ram[3355] = {9'd43,10'd43};
ram[3356] = {9'd47,10'd47};
ram[3357] = {9'd50,10'd50};
ram[3358] = {9'd53,10'd53};
ram[3359] = {9'd56,10'd56};
ram[3360] = {9'd59,10'd59};
ram[3361] = {9'd62,10'd62};
ram[3362] = {9'd65,10'd65};
ram[3363] = {9'd69,10'd69};
ram[3364] = {9'd72,10'd72};
ram[3365] = {9'd75,10'd75};
ram[3366] = {9'd78,10'd78};
ram[3367] = {9'd81,10'd81};
ram[3368] = {9'd84,10'd84};
ram[3369] = {9'd87,10'd87};
ram[3370] = {9'd91,10'd91};
ram[3371] = {9'd94,10'd94};
ram[3372] = {9'd97,10'd97};
ram[3373] = {-9'd100,10'd100};
ram[3374] = {-9'd97,10'd103};
ram[3375] = {-9'd94,10'd106};
ram[3376] = {-9'd91,10'd109};
ram[3377] = {-9'd88,10'd113};
ram[3378] = {-9'd85,10'd116};
ram[3379] = {-9'd81,10'd119};
ram[3380] = {-9'd78,10'd122};
ram[3381] = {-9'd75,10'd125};
ram[3382] = {-9'd72,10'd128};
ram[3383] = {-9'd69,10'd131};
ram[3384] = {-9'd66,10'd135};
ram[3385] = {-9'd63,10'd138};
ram[3386] = {-9'd59,10'd141};
ram[3387] = {-9'd56,10'd144};
ram[3388] = {-9'd53,10'd147};
ram[3389] = {-9'd50,10'd150};
ram[3390] = {-9'd47,10'd153};
ram[3391] = {-9'd44,10'd157};
ram[3392] = {-9'd41,10'd160};
ram[3393] = {-9'd37,10'd163};
ram[3394] = {-9'd34,10'd166};
ram[3395] = {-9'd31,10'd169};
ram[3396] = {-9'd28,10'd172};
ram[3397] = {-9'd25,10'd175};
ram[3398] = {-9'd22,10'd179};
ram[3399] = {-9'd19,10'd182};
ram[3400] = {-9'd15,10'd185};
ram[3401] = {-9'd12,10'd188};
ram[3402] = {-9'd9,10'd191};
ram[3403] = {-9'd6,10'd194};
ram[3404] = {-9'd3,10'd197};
ram[3405] = {9'd0,10'd201};
ram[3406] = {9'd3,10'd204};
ram[3407] = {9'd7,10'd207};
ram[3408] = {9'd10,10'd210};
ram[3409] = {9'd13,10'd213};
ram[3410] = {9'd16,10'd216};
ram[3411] = {9'd19,10'd219};
ram[3412] = {9'd22,10'd223};
ram[3413] = {9'd25,10'd226};
ram[3414] = {9'd29,10'd229};
ram[3415] = {9'd32,10'd232};
ram[3416] = {9'd35,10'd235};
ram[3417] = {9'd38,10'd238};
ram[3418] = {9'd41,10'd241};
ram[3419] = {9'd44,10'd245};
ram[3420] = {9'd47,10'd248};
ram[3421] = {9'd51,10'd251};
ram[3422] = {9'd54,10'd254};
ram[3423] = {9'd57,10'd257};
ram[3424] = {9'd60,10'd260};
ram[3425] = {9'd63,10'd263};
ram[3426] = {9'd66,10'd267};
ram[3427] = {9'd69,10'd270};
ram[3428] = {9'd73,10'd273};
ram[3429] = {9'd76,10'd276};
ram[3430] = {9'd79,10'd279};
ram[3431] = {9'd82,10'd282};
ram[3432] = {9'd85,10'd285};
ram[3433] = {9'd88,10'd289};
ram[3434] = {9'd91,10'd292};
ram[3435] = {9'd95,10'd295};
ram[3436] = {9'd98,10'd298};
ram[3437] = {-9'd99,10'd301};
ram[3438] = {-9'd96,10'd304};
ram[3439] = {-9'd93,10'd307};
ram[3440] = {-9'd90,10'd311};
ram[3441] = {-9'd87,10'd314};
ram[3442] = {-9'd84,10'd317};
ram[3443] = {-9'd81,10'd320};
ram[3444] = {-9'd77,10'd323};
ram[3445] = {-9'd74,10'd326};
ram[3446] = {-9'd71,10'd329};
ram[3447] = {-9'd68,10'd333};
ram[3448] = {-9'd65,10'd336};
ram[3449] = {-9'd62,10'd339};
ram[3450] = {-9'd59,10'd342};
ram[3451] = {-9'd55,10'd345};
ram[3452] = {-9'd52,10'd348};
ram[3453] = {-9'd49,10'd351};
ram[3454] = {-9'd46,10'd354};
ram[3455] = {-9'd43,10'd358};
ram[3456] = {-9'd43,10'd358};
ram[3457] = {-9'd40,10'd361};
ram[3458] = {-9'd37,10'd364};
ram[3459] = {-9'd33,10'd367};
ram[3460] = {-9'd30,10'd370};
ram[3461] = {-9'd27,10'd373};
ram[3462] = {-9'd24,10'd376};
ram[3463] = {-9'd21,10'd380};
ram[3464] = {-9'd18,10'd383};
ram[3465] = {-9'd15,10'd386};
ram[3466] = {-9'd11,10'd389};
ram[3467] = {-9'd8,10'd392};
ram[3468] = {-9'd5,10'd395};
ram[3469] = {-9'd2,10'd398};
ram[3470] = {9'd1,-10'd399};
ram[3471] = {9'd4,-10'd396};
ram[3472] = {9'd7,-10'd393};
ram[3473] = {9'd10,-10'd390};
ram[3474] = {9'd14,-10'd387};
ram[3475] = {9'd17,-10'd384};
ram[3476] = {9'd20,-10'd381};
ram[3477] = {9'd23,-10'd377};
ram[3478] = {9'd26,-10'd374};
ram[3479] = {9'd29,-10'd371};
ram[3480] = {9'd32,-10'd368};
ram[3481] = {9'd36,-10'd365};
ram[3482] = {9'd39,-10'd362};
ram[3483] = {9'd42,-10'd359};
ram[3484] = {9'd45,-10'd355};
ram[3485] = {9'd48,-10'd352};
ram[3486] = {9'd51,-10'd349};
ram[3487] = {9'd54,-10'd346};
ram[3488] = {9'd58,-10'd343};
ram[3489] = {9'd61,-10'd340};
ram[3490] = {9'd64,-10'd337};
ram[3491] = {9'd67,-10'd334};
ram[3492] = {9'd70,-10'd330};
ram[3493] = {9'd73,-10'd327};
ram[3494] = {9'd76,-10'd324};
ram[3495] = {9'd80,-10'd321};
ram[3496] = {9'd83,-10'd318};
ram[3497] = {9'd86,-10'd315};
ram[3498] = {9'd89,-10'd312};
ram[3499] = {9'd92,-10'd308};
ram[3500] = {9'd95,-10'd305};
ram[3501] = {9'd98,-10'd302};
ram[3502] = {-9'd99,-10'd299};
ram[3503] = {-9'd96,-10'd296};
ram[3504] = {-9'd92,-10'd293};
ram[3505] = {-9'd89,-10'd290};
ram[3506] = {-9'd86,-10'd286};
ram[3507] = {-9'd83,-10'd283};
ram[3508] = {-9'd80,-10'd280};
ram[3509] = {-9'd77,-10'd277};
ram[3510] = {-9'd74,-10'd274};
ram[3511] = {-9'd70,-10'd271};
ram[3512] = {-9'd67,-10'd268};
ram[3513] = {-9'd64,-10'd264};
ram[3514] = {-9'd61,-10'd261};
ram[3515] = {-9'd58,-10'd258};
ram[3516] = {-9'd55,-10'd255};
ram[3517] = {-9'd52,-10'd252};
ram[3518] = {-9'd48,-10'd249};
ram[3519] = {-9'd45,-10'd246};
ram[3520] = {-9'd42,-10'd242};
ram[3521] = {-9'd39,-10'd239};
ram[3522] = {-9'd36,-10'd236};
ram[3523] = {-9'd33,-10'd233};
ram[3524] = {-9'd30,-10'd230};
ram[3525] = {-9'd26,-10'd227};
ram[3526] = {-9'd23,-10'd224};
ram[3527] = {-9'd20,-10'd220};
ram[3528] = {-9'd17,-10'd217};
ram[3529] = {-9'd14,-10'd214};
ram[3530] = {-9'd11,-10'd211};
ram[3531] = {-9'd8,-10'd208};
ram[3532] = {-9'd4,-10'd205};
ram[3533] = {-9'd1,-10'd202};
ram[3534] = {9'd2,-10'd198};
ram[3535] = {9'd5,-10'd195};
ram[3536] = {9'd8,-10'd192};
ram[3537] = {9'd11,-10'd189};
ram[3538] = {9'd14,-10'd186};
ram[3539] = {9'd18,-10'd183};
ram[3540] = {9'd21,-10'd180};
ram[3541] = {9'd24,-10'd176};
ram[3542] = {9'd27,-10'd173};
ram[3543] = {9'd30,-10'd170};
ram[3544] = {9'd33,-10'd167};
ram[3545] = {9'd36,-10'd164};
ram[3546] = {9'd40,-10'd161};
ram[3547] = {9'd43,-10'd158};
ram[3548] = {9'd46,-10'd154};
ram[3549] = {9'd49,-10'd151};
ram[3550] = {9'd52,-10'd148};
ram[3551] = {9'd55,-10'd145};
ram[3552] = {9'd58,-10'd142};
ram[3553] = {9'd62,-10'd139};
ram[3554] = {9'd65,-10'd136};
ram[3555] = {9'd68,-10'd132};
ram[3556] = {9'd71,-10'd129};
ram[3557] = {9'd74,-10'd126};
ram[3558] = {9'd77,-10'd123};
ram[3559] = {9'd80,-10'd120};
ram[3560] = {9'd84,-10'd117};
ram[3561] = {9'd87,-10'd114};
ram[3562] = {9'd90,-10'd110};
ram[3563] = {9'd93,-10'd107};
ram[3564] = {9'd96,-10'd104};
ram[3565] = {9'd99,-10'd101};
ram[3566] = {-9'd98,-10'd98};
ram[3567] = {-9'd95,-10'd95};
ram[3568] = {-9'd92,-10'd92};
ram[3569] = {-9'd88,-10'd88};
ram[3570] = {-9'd85,-10'd85};
ram[3571] = {-9'd82,-10'd82};
ram[3572] = {-9'd79,-10'd79};
ram[3573] = {-9'd76,-10'd76};
ram[3574] = {-9'd73,-10'd73};
ram[3575] = {-9'd70,-10'd70};
ram[3576] = {-9'd66,-10'd66};
ram[3577] = {-9'd63,-10'd63};
ram[3578] = {-9'd60,-10'd60};
ram[3579] = {-9'd57,-10'd57};
ram[3580] = {-9'd54,-10'd54};
ram[3581] = {-9'd51,-10'd51};
ram[3582] = {-9'd48,-10'd48};
ram[3583] = {-9'd44,-10'd44};
ram[3584] = {-9'd44,-10'd44};
ram[3585] = {-9'd41,-10'd41};
ram[3586] = {-9'd38,-10'd38};
ram[3587] = {-9'd35,-10'd35};
ram[3588] = {-9'd32,-10'd32};
ram[3589] = {-9'd29,-10'd29};
ram[3590] = {-9'd26,-10'd26};
ram[3591] = {-9'd22,-10'd22};
ram[3592] = {-9'd19,-10'd19};
ram[3593] = {-9'd16,-10'd16};
ram[3594] = {-9'd13,-10'd13};
ram[3595] = {-9'd10,-10'd10};
ram[3596] = {-9'd7,-10'd7};
ram[3597] = {-9'd4,-10'd4};
ram[3598] = {9'd0,10'd0};
ram[3599] = {9'd3,10'd3};
ram[3600] = {9'd6,10'd6};
ram[3601] = {9'd9,10'd9};
ram[3602] = {9'd12,10'd12};
ram[3603] = {9'd15,10'd15};
ram[3604] = {9'd18,10'd18};
ram[3605] = {9'd21,10'd21};
ram[3606] = {9'd25,10'd25};
ram[3607] = {9'd28,10'd28};
ram[3608] = {9'd31,10'd31};
ram[3609] = {9'd34,10'd34};
ram[3610] = {9'd37,10'd37};
ram[3611] = {9'd40,10'd40};
ram[3612] = {9'd43,10'd43};
ram[3613] = {9'd47,10'd47};
ram[3614] = {9'd50,10'd50};
ram[3615] = {9'd53,10'd53};
ram[3616] = {9'd56,10'd56};
ram[3617] = {9'd59,10'd59};
ram[3618] = {9'd62,10'd62};
ram[3619] = {9'd65,10'd65};
ram[3620] = {9'd69,10'd69};
ram[3621] = {9'd72,10'd72};
ram[3622] = {9'd75,10'd75};
ram[3623] = {9'd78,10'd78};
ram[3624] = {9'd81,10'd81};
ram[3625] = {9'd84,10'd84};
ram[3626] = {9'd87,10'd87};
ram[3627] = {9'd91,10'd91};
ram[3628] = {9'd94,10'd94};
ram[3629] = {9'd97,10'd97};
ram[3630] = {-9'd100,10'd100};
ram[3631] = {-9'd97,10'd103};
ram[3632] = {-9'd94,10'd106};
ram[3633] = {-9'd91,10'd109};
ram[3634] = {-9'd88,10'd113};
ram[3635] = {-9'd85,10'd116};
ram[3636] = {-9'd81,10'd119};
ram[3637] = {-9'd78,10'd122};
ram[3638] = {-9'd75,10'd125};
ram[3639] = {-9'd72,10'd128};
ram[3640] = {-9'd69,10'd131};
ram[3641] = {-9'd66,10'd135};
ram[3642] = {-9'd63,10'd138};
ram[3643] = {-9'd59,10'd141};
ram[3644] = {-9'd56,10'd144};
ram[3645] = {-9'd53,10'd147};
ram[3646] = {-9'd50,10'd150};
ram[3647] = {-9'd47,10'd153};
ram[3648] = {-9'd44,10'd157};
ram[3649] = {-9'd41,10'd160};
ram[3650] = {-9'd37,10'd163};
ram[3651] = {-9'd34,10'd166};
ram[3652] = {-9'd31,10'd169};
ram[3653] = {-9'd28,10'd172};
ram[3654] = {-9'd25,10'd175};
ram[3655] = {-9'd22,10'd179};
ram[3656] = {-9'd19,10'd182};
ram[3657] = {-9'd15,10'd185};
ram[3658] = {-9'd12,10'd188};
ram[3659] = {-9'd9,10'd191};
ram[3660] = {-9'd6,10'd194};
ram[3661] = {-9'd3,10'd197};
ram[3662] = {9'd0,10'd201};
ram[3663] = {9'd3,10'd204};
ram[3664] = {9'd7,10'd207};
ram[3665] = {9'd10,10'd210};
ram[3666] = {9'd13,10'd213};
ram[3667] = {9'd16,10'd216};
ram[3668] = {9'd19,10'd219};
ram[3669] = {9'd22,10'd223};
ram[3670] = {9'd25,10'd226};
ram[3671] = {9'd29,10'd229};
ram[3672] = {9'd32,10'd232};
ram[3673] = {9'd35,10'd235};
ram[3674] = {9'd38,10'd238};
ram[3675] = {9'd41,10'd241};
ram[3676] = {9'd44,10'd245};
ram[3677] = {9'd47,10'd248};
ram[3678] = {9'd51,10'd251};
ram[3679] = {9'd54,10'd254};
ram[3680] = {9'd57,10'd257};
ram[3681] = {9'd60,10'd260};
ram[3682] = {9'd63,10'd263};
ram[3683] = {9'd66,10'd267};
ram[3684] = {9'd69,10'd270};
ram[3685] = {9'd73,10'd273};
ram[3686] = {9'd76,10'd276};
ram[3687] = {9'd79,10'd279};
ram[3688] = {9'd82,10'd282};
ram[3689] = {9'd85,10'd285};
ram[3690] = {9'd88,10'd289};
ram[3691] = {9'd91,10'd292};
ram[3692] = {9'd95,10'd295};
ram[3693] = {9'd98,10'd298};
ram[3694] = {-9'd99,10'd301};
ram[3695] = {-9'd96,10'd304};
ram[3696] = {-9'd93,10'd307};
ram[3697] = {-9'd90,10'd311};
ram[3698] = {-9'd87,10'd314};
ram[3699] = {-9'd84,10'd317};
ram[3700] = {-9'd81,10'd320};
ram[3701] = {-9'd77,10'd323};
ram[3702] = {-9'd74,10'd326};
ram[3703] = {-9'd71,10'd329};
ram[3704] = {-9'd68,10'd333};
ram[3705] = {-9'd65,10'd336};
ram[3706] = {-9'd62,10'd339};
ram[3707] = {-9'd59,10'd342};
ram[3708] = {-9'd55,10'd345};
ram[3709] = {-9'd52,10'd348};
ram[3710] = {-9'd49,10'd351};
ram[3711] = {-9'd46,10'd354};
ram[3712] = {-9'd46,10'd354};
ram[3713] = {-9'd43,10'd358};
ram[3714] = {-9'd40,10'd361};
ram[3715] = {-9'd37,10'd364};
ram[3716] = {-9'd33,10'd367};
ram[3717] = {-9'd30,10'd370};
ram[3718] = {-9'd27,10'd373};
ram[3719] = {-9'd24,10'd376};
ram[3720] = {-9'd21,10'd380};
ram[3721] = {-9'd18,10'd383};
ram[3722] = {-9'd15,10'd386};
ram[3723] = {-9'd11,10'd389};
ram[3724] = {-9'd8,10'd392};
ram[3725] = {-9'd5,10'd395};
ram[3726] = {-9'd2,10'd398};
ram[3727] = {9'd1,-10'd399};
ram[3728] = {9'd4,-10'd396};
ram[3729] = {9'd7,-10'd393};
ram[3730] = {9'd10,-10'd390};
ram[3731] = {9'd14,-10'd387};
ram[3732] = {9'd17,-10'd384};
ram[3733] = {9'd20,-10'd381};
ram[3734] = {9'd23,-10'd377};
ram[3735] = {9'd26,-10'd374};
ram[3736] = {9'd29,-10'd371};
ram[3737] = {9'd32,-10'd368};
ram[3738] = {9'd36,-10'd365};
ram[3739] = {9'd39,-10'd362};
ram[3740] = {9'd42,-10'd359};
ram[3741] = {9'd45,-10'd355};
ram[3742] = {9'd48,-10'd352};
ram[3743] = {9'd51,-10'd349};
ram[3744] = {9'd54,-10'd346};
ram[3745] = {9'd58,-10'd343};
ram[3746] = {9'd61,-10'd340};
ram[3747] = {9'd64,-10'd337};
ram[3748] = {9'd67,-10'd334};
ram[3749] = {9'd70,-10'd330};
ram[3750] = {9'd73,-10'd327};
ram[3751] = {9'd76,-10'd324};
ram[3752] = {9'd80,-10'd321};
ram[3753] = {9'd83,-10'd318};
ram[3754] = {9'd86,-10'd315};
ram[3755] = {9'd89,-10'd312};
ram[3756] = {9'd92,-10'd308};
ram[3757] = {9'd95,-10'd305};
ram[3758] = {9'd98,-10'd302};
ram[3759] = {-9'd99,-10'd299};
ram[3760] = {-9'd96,-10'd296};
ram[3761] = {-9'd92,-10'd293};
ram[3762] = {-9'd89,-10'd290};
ram[3763] = {-9'd86,-10'd286};
ram[3764] = {-9'd83,-10'd283};
ram[3765] = {-9'd80,-10'd280};
ram[3766] = {-9'd77,-10'd277};
ram[3767] = {-9'd74,-10'd274};
ram[3768] = {-9'd70,-10'd271};
ram[3769] = {-9'd67,-10'd268};
ram[3770] = {-9'd64,-10'd264};
ram[3771] = {-9'd61,-10'd261};
ram[3772] = {-9'd58,-10'd258};
ram[3773] = {-9'd55,-10'd255};
ram[3774] = {-9'd52,-10'd252};
ram[3775] = {-9'd48,-10'd249};
ram[3776] = {-9'd45,-10'd246};
ram[3777] = {-9'd42,-10'd242};
ram[3778] = {-9'd39,-10'd239};
ram[3779] = {-9'd36,-10'd236};
ram[3780] = {-9'd33,-10'd233};
ram[3781] = {-9'd30,-10'd230};
ram[3782] = {-9'd26,-10'd227};
ram[3783] = {-9'd23,-10'd224};
ram[3784] = {-9'd20,-10'd220};
ram[3785] = {-9'd17,-10'd217};
ram[3786] = {-9'd14,-10'd214};
ram[3787] = {-9'd11,-10'd211};
ram[3788] = {-9'd8,-10'd208};
ram[3789] = {-9'd4,-10'd205};
ram[3790] = {-9'd1,-10'd202};
ram[3791] = {9'd2,-10'd198};
ram[3792] = {9'd5,-10'd195};
ram[3793] = {9'd8,-10'd192};
ram[3794] = {9'd11,-10'd189};
ram[3795] = {9'd14,-10'd186};
ram[3796] = {9'd18,-10'd183};
ram[3797] = {9'd21,-10'd180};
ram[3798] = {9'd24,-10'd176};
ram[3799] = {9'd27,-10'd173};
ram[3800] = {9'd30,-10'd170};
ram[3801] = {9'd33,-10'd167};
ram[3802] = {9'd36,-10'd164};
ram[3803] = {9'd40,-10'd161};
ram[3804] = {9'd43,-10'd158};
ram[3805] = {9'd46,-10'd154};
ram[3806] = {9'd49,-10'd151};
ram[3807] = {9'd52,-10'd148};
ram[3808] = {9'd55,-10'd145};
ram[3809] = {9'd58,-10'd142};
ram[3810] = {9'd62,-10'd139};
ram[3811] = {9'd65,-10'd136};
ram[3812] = {9'd68,-10'd132};
ram[3813] = {9'd71,-10'd129};
ram[3814] = {9'd74,-10'd126};
ram[3815] = {9'd77,-10'd123};
ram[3816] = {9'd80,-10'd120};
ram[3817] = {9'd84,-10'd117};
ram[3818] = {9'd87,-10'd114};
ram[3819] = {9'd90,-10'd110};
ram[3820] = {9'd93,-10'd107};
ram[3821] = {9'd96,-10'd104};
ram[3822] = {9'd99,-10'd101};
ram[3823] = {-9'd98,-10'd98};
ram[3824] = {-9'd95,-10'd95};
ram[3825] = {-9'd92,-10'd92};
ram[3826] = {-9'd88,-10'd88};
ram[3827] = {-9'd85,-10'd85};
ram[3828] = {-9'd82,-10'd82};
ram[3829] = {-9'd79,-10'd79};
ram[3830] = {-9'd76,-10'd76};
ram[3831] = {-9'd73,-10'd73};
ram[3832] = {-9'd70,-10'd70};
ram[3833] = {-9'd66,-10'd66};
ram[3834] = {-9'd63,-10'd63};
ram[3835] = {-9'd60,-10'd60};
ram[3836] = {-9'd57,-10'd57};
ram[3837] = {-9'd54,-10'd54};
ram[3838] = {-9'd51,-10'd51};
ram[3839] = {-9'd48,-10'd48};
ram[3840] = {-9'd48,-10'd48};
ram[3841] = {-9'd44,-10'd44};
ram[3842] = {-9'd41,-10'd41};
ram[3843] = {-9'd38,-10'd38};
ram[3844] = {-9'd35,-10'd35};
ram[3845] = {-9'd32,-10'd32};
ram[3846] = {-9'd29,-10'd29};
ram[3847] = {-9'd26,-10'd26};
ram[3848] = {-9'd22,-10'd22};
ram[3849] = {-9'd19,-10'd19};
ram[3850] = {-9'd16,-10'd16};
ram[3851] = {-9'd13,-10'd13};
ram[3852] = {-9'd10,-10'd10};
ram[3853] = {-9'd7,-10'd7};
ram[3854] = {-9'd4,-10'd4};
ram[3855] = {9'd0,10'd0};
ram[3856] = {9'd3,10'd3};
ram[3857] = {9'd6,10'd6};
ram[3858] = {9'd9,10'd9};
ram[3859] = {9'd12,10'd12};
ram[3860] = {9'd15,10'd15};
ram[3861] = {9'd18,10'd18};
ram[3862] = {9'd21,10'd21};
ram[3863] = {9'd25,10'd25};
ram[3864] = {9'd28,10'd28};
ram[3865] = {9'd31,10'd31};
ram[3866] = {9'd34,10'd34};
ram[3867] = {9'd37,10'd37};
ram[3868] = {9'd40,10'd40};
ram[3869] = {9'd43,10'd43};
ram[3870] = {9'd47,10'd47};
ram[3871] = {9'd50,10'd50};
ram[3872] = {9'd53,10'd53};
ram[3873] = {9'd56,10'd56};
ram[3874] = {9'd59,10'd59};
ram[3875] = {9'd62,10'd62};
ram[3876] = {9'd65,10'd65};
ram[3877] = {9'd69,10'd69};
ram[3878] = {9'd72,10'd72};
ram[3879] = {9'd75,10'd75};
ram[3880] = {9'd78,10'd78};
ram[3881] = {9'd81,10'd81};
ram[3882] = {9'd84,10'd84};
ram[3883] = {9'd87,10'd87};
ram[3884] = {9'd91,10'd91};
ram[3885] = {9'd94,10'd94};
ram[3886] = {9'd97,10'd97};
ram[3887] = {-9'd100,10'd100};
ram[3888] = {-9'd97,10'd103};
ram[3889] = {-9'd94,10'd106};
ram[3890] = {-9'd91,10'd109};
ram[3891] = {-9'd88,10'd113};
ram[3892] = {-9'd85,10'd116};
ram[3893] = {-9'd81,10'd119};
ram[3894] = {-9'd78,10'd122};
ram[3895] = {-9'd75,10'd125};
ram[3896] = {-9'd72,10'd128};
ram[3897] = {-9'd69,10'd131};
ram[3898] = {-9'd66,10'd135};
ram[3899] = {-9'd63,10'd138};
ram[3900] = {-9'd59,10'd141};
ram[3901] = {-9'd56,10'd144};
ram[3902] = {-9'd53,10'd147};
ram[3903] = {-9'd50,10'd150};
ram[3904] = {-9'd47,10'd153};
ram[3905] = {-9'd44,10'd157};
ram[3906] = {-9'd41,10'd160};
ram[3907] = {-9'd37,10'd163};
ram[3908] = {-9'd34,10'd166};
ram[3909] = {-9'd31,10'd169};
ram[3910] = {-9'd28,10'd172};
ram[3911] = {-9'd25,10'd175};
ram[3912] = {-9'd22,10'd179};
ram[3913] = {-9'd19,10'd182};
ram[3914] = {-9'd15,10'd185};
ram[3915] = {-9'd12,10'd188};
ram[3916] = {-9'd9,10'd191};
ram[3917] = {-9'd6,10'd194};
ram[3918] = {-9'd3,10'd197};
ram[3919] = {9'd0,10'd201};
ram[3920] = {9'd3,10'd204};
ram[3921] = {9'd7,10'd207};
ram[3922] = {9'd10,10'd210};
ram[3923] = {9'd13,10'd213};
ram[3924] = {9'd16,10'd216};
ram[3925] = {9'd19,10'd219};
ram[3926] = {9'd22,10'd223};
ram[3927] = {9'd25,10'd226};
ram[3928] = {9'd29,10'd229};
ram[3929] = {9'd32,10'd232};
ram[3930] = {9'd35,10'd235};
ram[3931] = {9'd38,10'd238};
ram[3932] = {9'd41,10'd241};
ram[3933] = {9'd44,10'd245};
ram[3934] = {9'd47,10'd248};
ram[3935] = {9'd51,10'd251};
ram[3936] = {9'd54,10'd254};
ram[3937] = {9'd57,10'd257};
ram[3938] = {9'd60,10'd260};
ram[3939] = {9'd63,10'd263};
ram[3940] = {9'd66,10'd267};
ram[3941] = {9'd69,10'd270};
ram[3942] = {9'd73,10'd273};
ram[3943] = {9'd76,10'd276};
ram[3944] = {9'd79,10'd279};
ram[3945] = {9'd82,10'd282};
ram[3946] = {9'd85,10'd285};
ram[3947] = {9'd88,10'd289};
ram[3948] = {9'd91,10'd292};
ram[3949] = {9'd95,10'd295};
ram[3950] = {9'd98,10'd298};
ram[3951] = {-9'd99,10'd301};
ram[3952] = {-9'd96,10'd304};
ram[3953] = {-9'd93,10'd307};
ram[3954] = {-9'd90,10'd311};
ram[3955] = {-9'd87,10'd314};
ram[3956] = {-9'd84,10'd317};
ram[3957] = {-9'd81,10'd320};
ram[3958] = {-9'd77,10'd323};
ram[3959] = {-9'd74,10'd326};
ram[3960] = {-9'd71,10'd329};
ram[3961] = {-9'd68,10'd333};
ram[3962] = {-9'd65,10'd336};
ram[3963] = {-9'd62,10'd339};
ram[3964] = {-9'd59,10'd342};
ram[3965] = {-9'd55,10'd345};
ram[3966] = {-9'd52,10'd348};
ram[3967] = {-9'd49,10'd351};
ram[3968] = {-9'd49,10'd351};
ram[3969] = {-9'd46,10'd354};
ram[3970] = {-9'd43,10'd358};
ram[3971] = {-9'd40,10'd361};
ram[3972] = {-9'd37,10'd364};
ram[3973] = {-9'd33,10'd367};
ram[3974] = {-9'd30,10'd370};
ram[3975] = {-9'd27,10'd373};
ram[3976] = {-9'd24,10'd376};
ram[3977] = {-9'd21,10'd380};
ram[3978] = {-9'd18,10'd383};
ram[3979] = {-9'd15,10'd386};
ram[3980] = {-9'd11,10'd389};
ram[3981] = {-9'd8,10'd392};
ram[3982] = {-9'd5,10'd395};
ram[3983] = {-9'd2,10'd398};
ram[3984] = {9'd1,-10'd399};
ram[3985] = {9'd4,-10'd396};
ram[3986] = {9'd7,-10'd393};
ram[3987] = {9'd10,-10'd390};
ram[3988] = {9'd14,-10'd387};
ram[3989] = {9'd17,-10'd384};
ram[3990] = {9'd20,-10'd381};
ram[3991] = {9'd23,-10'd377};
ram[3992] = {9'd26,-10'd374};
ram[3993] = {9'd29,-10'd371};
ram[3994] = {9'd32,-10'd368};
ram[3995] = {9'd36,-10'd365};
ram[3996] = {9'd39,-10'd362};
ram[3997] = {9'd42,-10'd359};
ram[3998] = {9'd45,-10'd355};
ram[3999] = {9'd48,-10'd352};
ram[4000] = {9'd51,-10'd349};
ram[4001] = {9'd54,-10'd346};
ram[4002] = {9'd58,-10'd343};
ram[4003] = {9'd61,-10'd340};
ram[4004] = {9'd64,-10'd337};
ram[4005] = {9'd67,-10'd334};
ram[4006] = {9'd70,-10'd330};
ram[4007] = {9'd73,-10'd327};
ram[4008] = {9'd76,-10'd324};
ram[4009] = {9'd80,-10'd321};
ram[4010] = {9'd83,-10'd318};
ram[4011] = {9'd86,-10'd315};
ram[4012] = {9'd89,-10'd312};
ram[4013] = {9'd92,-10'd308};
ram[4014] = {9'd95,-10'd305};
ram[4015] = {9'd98,-10'd302};
ram[4016] = {-9'd99,-10'd299};
ram[4017] = {-9'd96,-10'd296};
ram[4018] = {-9'd92,-10'd293};
ram[4019] = {-9'd89,-10'd290};
ram[4020] = {-9'd86,-10'd286};
ram[4021] = {-9'd83,-10'd283};
ram[4022] = {-9'd80,-10'd280};
ram[4023] = {-9'd77,-10'd277};
ram[4024] = {-9'd74,-10'd274};
ram[4025] = {-9'd70,-10'd271};
ram[4026] = {-9'd67,-10'd268};
ram[4027] = {-9'd64,-10'd264};
ram[4028] = {-9'd61,-10'd261};
ram[4029] = {-9'd58,-10'd258};
ram[4030] = {-9'd55,-10'd255};
ram[4031] = {-9'd52,-10'd252};
ram[4032] = {-9'd48,-10'd249};
ram[4033] = {-9'd45,-10'd246};
ram[4034] = {-9'd42,-10'd242};
ram[4035] = {-9'd39,-10'd239};
ram[4036] = {-9'd36,-10'd236};
ram[4037] = {-9'd33,-10'd233};
ram[4038] = {-9'd30,-10'd230};
ram[4039] = {-9'd26,-10'd227};
ram[4040] = {-9'd23,-10'd224};
ram[4041] = {-9'd20,-10'd220};
ram[4042] = {-9'd17,-10'd217};
ram[4043] = {-9'd14,-10'd214};
ram[4044] = {-9'd11,-10'd211};
ram[4045] = {-9'd8,-10'd208};
ram[4046] = {-9'd4,-10'd205};
ram[4047] = {-9'd1,-10'd202};
ram[4048] = {9'd2,-10'd198};
ram[4049] = {9'd5,-10'd195};
ram[4050] = {9'd8,-10'd192};
ram[4051] = {9'd11,-10'd189};
ram[4052] = {9'd14,-10'd186};
ram[4053] = {9'd18,-10'd183};
ram[4054] = {9'd21,-10'd180};
ram[4055] = {9'd24,-10'd176};
ram[4056] = {9'd27,-10'd173};
ram[4057] = {9'd30,-10'd170};
ram[4058] = {9'd33,-10'd167};
ram[4059] = {9'd36,-10'd164};
ram[4060] = {9'd40,-10'd161};
ram[4061] = {9'd43,-10'd158};
ram[4062] = {9'd46,-10'd154};
ram[4063] = {9'd49,-10'd151};
ram[4064] = {9'd52,-10'd148};
ram[4065] = {9'd55,-10'd145};
ram[4066] = {9'd58,-10'd142};
ram[4067] = {9'd62,-10'd139};
ram[4068] = {9'd65,-10'd136};
ram[4069] = {9'd68,-10'd132};
ram[4070] = {9'd71,-10'd129};
ram[4071] = {9'd74,-10'd126};
ram[4072] = {9'd77,-10'd123};
ram[4073] = {9'd80,-10'd120};
ram[4074] = {9'd84,-10'd117};
ram[4075] = {9'd87,-10'd114};
ram[4076] = {9'd90,-10'd110};
ram[4077] = {9'd93,-10'd107};
ram[4078] = {9'd96,-10'd104};
ram[4079] = {9'd99,-10'd101};
ram[4080] = {-9'd98,-10'd98};
ram[4081] = {-9'd95,-10'd95};
ram[4082] = {-9'd92,-10'd92};
ram[4083] = {-9'd88,-10'd88};
ram[4084] = {-9'd85,-10'd85};
ram[4085] = {-9'd82,-10'd82};
ram[4086] = {-9'd79,-10'd79};
ram[4087] = {-9'd76,-10'd76};
ram[4088] = {-9'd73,-10'd73};
ram[4089] = {-9'd70,-10'd70};
ram[4090] = {-9'd66,-10'd66};
ram[4091] = {-9'd63,-10'd63};
ram[4092] = {-9'd60,-10'd60};
ram[4093] = {-9'd57,-10'd57};
ram[4094] = {-9'd54,-10'd54};
ram[4095] = {-9'd51,-10'd51};
ram[4096] = {-9'd51,-10'd51};
ram[4097] = {-9'd48,-10'd48};
ram[4098] = {-9'd44,-10'd44};
ram[4099] = {-9'd41,-10'd41};
ram[4100] = {-9'd38,-10'd38};
ram[4101] = {-9'd35,-10'd35};
ram[4102] = {-9'd32,-10'd32};
ram[4103] = {-9'd29,-10'd29};
ram[4104] = {-9'd26,-10'd26};
ram[4105] = {-9'd22,-10'd22};
ram[4106] = {-9'd19,-10'd19};
ram[4107] = {-9'd16,-10'd16};
ram[4108] = {-9'd13,-10'd13};
ram[4109] = {-9'd10,-10'd10};
ram[4110] = {-9'd7,-10'd7};
ram[4111] = {-9'd4,-10'd4};
ram[4112] = {9'd0,10'd0};
ram[4113] = {9'd3,10'd3};
ram[4114] = {9'd6,10'd6};
ram[4115] = {9'd9,10'd9};
ram[4116] = {9'd12,10'd12};
ram[4117] = {9'd15,10'd15};
ram[4118] = {9'd18,10'd18};
ram[4119] = {9'd21,10'd21};
ram[4120] = {9'd25,10'd25};
ram[4121] = {9'd28,10'd28};
ram[4122] = {9'd31,10'd31};
ram[4123] = {9'd34,10'd34};
ram[4124] = {9'd37,10'd37};
ram[4125] = {9'd40,10'd40};
ram[4126] = {9'd43,10'd43};
ram[4127] = {9'd47,10'd47};
ram[4128] = {9'd50,10'd50};
ram[4129] = {9'd53,10'd53};
ram[4130] = {9'd56,10'd56};
ram[4131] = {9'd59,10'd59};
ram[4132] = {9'd62,10'd62};
ram[4133] = {9'd65,10'd65};
ram[4134] = {9'd69,10'd69};
ram[4135] = {9'd72,10'd72};
ram[4136] = {9'd75,10'd75};
ram[4137] = {9'd78,10'd78};
ram[4138] = {9'd81,10'd81};
ram[4139] = {9'd84,10'd84};
ram[4140] = {9'd87,10'd87};
ram[4141] = {9'd91,10'd91};
ram[4142] = {9'd94,10'd94};
ram[4143] = {9'd97,10'd97};
ram[4144] = {-9'd100,10'd100};
ram[4145] = {-9'd97,10'd103};
ram[4146] = {-9'd94,10'd106};
ram[4147] = {-9'd91,10'd109};
ram[4148] = {-9'd88,10'd113};
ram[4149] = {-9'd85,10'd116};
ram[4150] = {-9'd81,10'd119};
ram[4151] = {-9'd78,10'd122};
ram[4152] = {-9'd75,10'd125};
ram[4153] = {-9'd72,10'd128};
ram[4154] = {-9'd69,10'd131};
ram[4155] = {-9'd66,10'd135};
ram[4156] = {-9'd63,10'd138};
ram[4157] = {-9'd59,10'd141};
ram[4158] = {-9'd56,10'd144};
ram[4159] = {-9'd53,10'd147};
ram[4160] = {-9'd50,10'd150};
ram[4161] = {-9'd47,10'd153};
ram[4162] = {-9'd44,10'd157};
ram[4163] = {-9'd41,10'd160};
ram[4164] = {-9'd37,10'd163};
ram[4165] = {-9'd34,10'd166};
ram[4166] = {-9'd31,10'd169};
ram[4167] = {-9'd28,10'd172};
ram[4168] = {-9'd25,10'd175};
ram[4169] = {-9'd22,10'd179};
ram[4170] = {-9'd19,10'd182};
ram[4171] = {-9'd15,10'd185};
ram[4172] = {-9'd12,10'd188};
ram[4173] = {-9'd9,10'd191};
ram[4174] = {-9'd6,10'd194};
ram[4175] = {-9'd3,10'd197};
ram[4176] = {9'd0,10'd201};
ram[4177] = {9'd3,10'd204};
ram[4178] = {9'd7,10'd207};
ram[4179] = {9'd10,10'd210};
ram[4180] = {9'd13,10'd213};
ram[4181] = {9'd16,10'd216};
ram[4182] = {9'd19,10'd219};
ram[4183] = {9'd22,10'd223};
ram[4184] = {9'd25,10'd226};
ram[4185] = {9'd29,10'd229};
ram[4186] = {9'd32,10'd232};
ram[4187] = {9'd35,10'd235};
ram[4188] = {9'd38,10'd238};
ram[4189] = {9'd41,10'd241};
ram[4190] = {9'd44,10'd245};
ram[4191] = {9'd47,10'd248};
ram[4192] = {9'd51,10'd251};
ram[4193] = {9'd54,10'd254};
ram[4194] = {9'd57,10'd257};
ram[4195] = {9'd60,10'd260};
ram[4196] = {9'd63,10'd263};
ram[4197] = {9'd66,10'd267};
ram[4198] = {9'd69,10'd270};
ram[4199] = {9'd73,10'd273};
ram[4200] = {9'd76,10'd276};
ram[4201] = {9'd79,10'd279};
ram[4202] = {9'd82,10'd282};
ram[4203] = {9'd85,10'd285};
ram[4204] = {9'd88,10'd289};
ram[4205] = {9'd91,10'd292};
ram[4206] = {9'd95,10'd295};
ram[4207] = {9'd98,10'd298};
ram[4208] = {-9'd99,10'd301};
ram[4209] = {-9'd96,10'd304};
ram[4210] = {-9'd93,10'd307};
ram[4211] = {-9'd90,10'd311};
ram[4212] = {-9'd87,10'd314};
ram[4213] = {-9'd84,10'd317};
ram[4214] = {-9'd81,10'd320};
ram[4215] = {-9'd77,10'd323};
ram[4216] = {-9'd74,10'd326};
ram[4217] = {-9'd71,10'd329};
ram[4218] = {-9'd68,10'd333};
ram[4219] = {-9'd65,10'd336};
ram[4220] = {-9'd62,10'd339};
ram[4221] = {-9'd59,10'd342};
ram[4222] = {-9'd55,10'd345};
ram[4223] = {-9'd52,10'd348};
ram[4224] = {-9'd52,10'd348};
ram[4225] = {-9'd49,10'd351};
ram[4226] = {-9'd46,10'd354};
ram[4227] = {-9'd43,10'd358};
ram[4228] = {-9'd40,10'd361};
ram[4229] = {-9'd37,10'd364};
ram[4230] = {-9'd33,10'd367};
ram[4231] = {-9'd30,10'd370};
ram[4232] = {-9'd27,10'd373};
ram[4233] = {-9'd24,10'd376};
ram[4234] = {-9'd21,10'd380};
ram[4235] = {-9'd18,10'd383};
ram[4236] = {-9'd15,10'd386};
ram[4237] = {-9'd11,10'd389};
ram[4238] = {-9'd8,10'd392};
ram[4239] = {-9'd5,10'd395};
ram[4240] = {-9'd2,10'd398};
ram[4241] = {9'd1,-10'd399};
ram[4242] = {9'd4,-10'd396};
ram[4243] = {9'd7,-10'd393};
ram[4244] = {9'd10,-10'd390};
ram[4245] = {9'd14,-10'd387};
ram[4246] = {9'd17,-10'd384};
ram[4247] = {9'd20,-10'd381};
ram[4248] = {9'd23,-10'd377};
ram[4249] = {9'd26,-10'd374};
ram[4250] = {9'd29,-10'd371};
ram[4251] = {9'd32,-10'd368};
ram[4252] = {9'd36,-10'd365};
ram[4253] = {9'd39,-10'd362};
ram[4254] = {9'd42,-10'd359};
ram[4255] = {9'd45,-10'd355};
ram[4256] = {9'd48,-10'd352};
ram[4257] = {9'd51,-10'd349};
ram[4258] = {9'd54,-10'd346};
ram[4259] = {9'd58,-10'd343};
ram[4260] = {9'd61,-10'd340};
ram[4261] = {9'd64,-10'd337};
ram[4262] = {9'd67,-10'd334};
ram[4263] = {9'd70,-10'd330};
ram[4264] = {9'd73,-10'd327};
ram[4265] = {9'd76,-10'd324};
ram[4266] = {9'd80,-10'd321};
ram[4267] = {9'd83,-10'd318};
ram[4268] = {9'd86,-10'd315};
ram[4269] = {9'd89,-10'd312};
ram[4270] = {9'd92,-10'd308};
ram[4271] = {9'd95,-10'd305};
ram[4272] = {9'd98,-10'd302};
ram[4273] = {-9'd99,-10'd299};
ram[4274] = {-9'd96,-10'd296};
ram[4275] = {-9'd92,-10'd293};
ram[4276] = {-9'd89,-10'd290};
ram[4277] = {-9'd86,-10'd286};
ram[4278] = {-9'd83,-10'd283};
ram[4279] = {-9'd80,-10'd280};
ram[4280] = {-9'd77,-10'd277};
ram[4281] = {-9'd74,-10'd274};
ram[4282] = {-9'd70,-10'd271};
ram[4283] = {-9'd67,-10'd268};
ram[4284] = {-9'd64,-10'd264};
ram[4285] = {-9'd61,-10'd261};
ram[4286] = {-9'd58,-10'd258};
ram[4287] = {-9'd55,-10'd255};
ram[4288] = {-9'd52,-10'd252};
ram[4289] = {-9'd48,-10'd249};
ram[4290] = {-9'd45,-10'd246};
ram[4291] = {-9'd42,-10'd242};
ram[4292] = {-9'd39,-10'd239};
ram[4293] = {-9'd36,-10'd236};
ram[4294] = {-9'd33,-10'd233};
ram[4295] = {-9'd30,-10'd230};
ram[4296] = {-9'd26,-10'd227};
ram[4297] = {-9'd23,-10'd224};
ram[4298] = {-9'd20,-10'd220};
ram[4299] = {-9'd17,-10'd217};
ram[4300] = {-9'd14,-10'd214};
ram[4301] = {-9'd11,-10'd211};
ram[4302] = {-9'd8,-10'd208};
ram[4303] = {-9'd4,-10'd205};
ram[4304] = {-9'd1,-10'd202};
ram[4305] = {9'd2,-10'd198};
ram[4306] = {9'd5,-10'd195};
ram[4307] = {9'd8,-10'd192};
ram[4308] = {9'd11,-10'd189};
ram[4309] = {9'd14,-10'd186};
ram[4310] = {9'd18,-10'd183};
ram[4311] = {9'd21,-10'd180};
ram[4312] = {9'd24,-10'd176};
ram[4313] = {9'd27,-10'd173};
ram[4314] = {9'd30,-10'd170};
ram[4315] = {9'd33,-10'd167};
ram[4316] = {9'd36,-10'd164};
ram[4317] = {9'd40,-10'd161};
ram[4318] = {9'd43,-10'd158};
ram[4319] = {9'd46,-10'd154};
ram[4320] = {9'd49,-10'd151};
ram[4321] = {9'd52,-10'd148};
ram[4322] = {9'd55,-10'd145};
ram[4323] = {9'd58,-10'd142};
ram[4324] = {9'd62,-10'd139};
ram[4325] = {9'd65,-10'd136};
ram[4326] = {9'd68,-10'd132};
ram[4327] = {9'd71,-10'd129};
ram[4328] = {9'd74,-10'd126};
ram[4329] = {9'd77,-10'd123};
ram[4330] = {9'd80,-10'd120};
ram[4331] = {9'd84,-10'd117};
ram[4332] = {9'd87,-10'd114};
ram[4333] = {9'd90,-10'd110};
ram[4334] = {9'd93,-10'd107};
ram[4335] = {9'd96,-10'd104};
ram[4336] = {9'd99,-10'd101};
ram[4337] = {-9'd98,-10'd98};
ram[4338] = {-9'd95,-10'd95};
ram[4339] = {-9'd92,-10'd92};
ram[4340] = {-9'd88,-10'd88};
ram[4341] = {-9'd85,-10'd85};
ram[4342] = {-9'd82,-10'd82};
ram[4343] = {-9'd79,-10'd79};
ram[4344] = {-9'd76,-10'd76};
ram[4345] = {-9'd73,-10'd73};
ram[4346] = {-9'd70,-10'd70};
ram[4347] = {-9'd66,-10'd66};
ram[4348] = {-9'd63,-10'd63};
ram[4349] = {-9'd60,-10'd60};
ram[4350] = {-9'd57,-10'd57};
ram[4351] = {-9'd54,-10'd54};
ram[4352] = {-9'd54,-10'd54};
ram[4353] = {-9'd51,-10'd51};
ram[4354] = {-9'd48,-10'd48};
ram[4355] = {-9'd44,-10'd44};
ram[4356] = {-9'd41,-10'd41};
ram[4357] = {-9'd38,-10'd38};
ram[4358] = {-9'd35,-10'd35};
ram[4359] = {-9'd32,-10'd32};
ram[4360] = {-9'd29,-10'd29};
ram[4361] = {-9'd26,-10'd26};
ram[4362] = {-9'd22,-10'd22};
ram[4363] = {-9'd19,-10'd19};
ram[4364] = {-9'd16,-10'd16};
ram[4365] = {-9'd13,-10'd13};
ram[4366] = {-9'd10,-10'd10};
ram[4367] = {-9'd7,-10'd7};
ram[4368] = {-9'd4,-10'd4};
ram[4369] = {9'd0,10'd0};
ram[4370] = {9'd3,10'd3};
ram[4371] = {9'd6,10'd6};
ram[4372] = {9'd9,10'd9};
ram[4373] = {9'd12,10'd12};
ram[4374] = {9'd15,10'd15};
ram[4375] = {9'd18,10'd18};
ram[4376] = {9'd21,10'd21};
ram[4377] = {9'd25,10'd25};
ram[4378] = {9'd28,10'd28};
ram[4379] = {9'd31,10'd31};
ram[4380] = {9'd34,10'd34};
ram[4381] = {9'd37,10'd37};
ram[4382] = {9'd40,10'd40};
ram[4383] = {9'd43,10'd43};
ram[4384] = {9'd47,10'd47};
ram[4385] = {9'd50,10'd50};
ram[4386] = {9'd53,10'd53};
ram[4387] = {9'd56,10'd56};
ram[4388] = {9'd59,10'd59};
ram[4389] = {9'd62,10'd62};
ram[4390] = {9'd65,10'd65};
ram[4391] = {9'd69,10'd69};
ram[4392] = {9'd72,10'd72};
ram[4393] = {9'd75,10'd75};
ram[4394] = {9'd78,10'd78};
ram[4395] = {9'd81,10'd81};
ram[4396] = {9'd84,10'd84};
ram[4397] = {9'd87,10'd87};
ram[4398] = {9'd91,10'd91};
ram[4399] = {9'd94,10'd94};
ram[4400] = {9'd97,10'd97};
ram[4401] = {-9'd100,10'd100};
ram[4402] = {-9'd97,10'd103};
ram[4403] = {-9'd94,10'd106};
ram[4404] = {-9'd91,10'd109};
ram[4405] = {-9'd88,10'd113};
ram[4406] = {-9'd85,10'd116};
ram[4407] = {-9'd81,10'd119};
ram[4408] = {-9'd78,10'd122};
ram[4409] = {-9'd75,10'd125};
ram[4410] = {-9'd72,10'd128};
ram[4411] = {-9'd69,10'd131};
ram[4412] = {-9'd66,10'd135};
ram[4413] = {-9'd63,10'd138};
ram[4414] = {-9'd59,10'd141};
ram[4415] = {-9'd56,10'd144};
ram[4416] = {-9'd53,10'd147};
ram[4417] = {-9'd50,10'd150};
ram[4418] = {-9'd47,10'd153};
ram[4419] = {-9'd44,10'd157};
ram[4420] = {-9'd41,10'd160};
ram[4421] = {-9'd37,10'd163};
ram[4422] = {-9'd34,10'd166};
ram[4423] = {-9'd31,10'd169};
ram[4424] = {-9'd28,10'd172};
ram[4425] = {-9'd25,10'd175};
ram[4426] = {-9'd22,10'd179};
ram[4427] = {-9'd19,10'd182};
ram[4428] = {-9'd15,10'd185};
ram[4429] = {-9'd12,10'd188};
ram[4430] = {-9'd9,10'd191};
ram[4431] = {-9'd6,10'd194};
ram[4432] = {-9'd3,10'd197};
ram[4433] = {9'd0,10'd201};
ram[4434] = {9'd3,10'd204};
ram[4435] = {9'd7,10'd207};
ram[4436] = {9'd10,10'd210};
ram[4437] = {9'd13,10'd213};
ram[4438] = {9'd16,10'd216};
ram[4439] = {9'd19,10'd219};
ram[4440] = {9'd22,10'd223};
ram[4441] = {9'd25,10'd226};
ram[4442] = {9'd29,10'd229};
ram[4443] = {9'd32,10'd232};
ram[4444] = {9'd35,10'd235};
ram[4445] = {9'd38,10'd238};
ram[4446] = {9'd41,10'd241};
ram[4447] = {9'd44,10'd245};
ram[4448] = {9'd47,10'd248};
ram[4449] = {9'd51,10'd251};
ram[4450] = {9'd54,10'd254};
ram[4451] = {9'd57,10'd257};
ram[4452] = {9'd60,10'd260};
ram[4453] = {9'd63,10'd263};
ram[4454] = {9'd66,10'd267};
ram[4455] = {9'd69,10'd270};
ram[4456] = {9'd73,10'd273};
ram[4457] = {9'd76,10'd276};
ram[4458] = {9'd79,10'd279};
ram[4459] = {9'd82,10'd282};
ram[4460] = {9'd85,10'd285};
ram[4461] = {9'd88,10'd289};
ram[4462] = {9'd91,10'd292};
ram[4463] = {9'd95,10'd295};
ram[4464] = {9'd98,10'd298};
ram[4465] = {-9'd99,10'd301};
ram[4466] = {-9'd96,10'd304};
ram[4467] = {-9'd93,10'd307};
ram[4468] = {-9'd90,10'd311};
ram[4469] = {-9'd87,10'd314};
ram[4470] = {-9'd84,10'd317};
ram[4471] = {-9'd81,10'd320};
ram[4472] = {-9'd77,10'd323};
ram[4473] = {-9'd74,10'd326};
ram[4474] = {-9'd71,10'd329};
ram[4475] = {-9'd68,10'd333};
ram[4476] = {-9'd65,10'd336};
ram[4477] = {-9'd62,10'd339};
ram[4478] = {-9'd59,10'd342};
ram[4479] = {-9'd55,10'd345};
ram[4480] = {-9'd55,10'd345};
ram[4481] = {-9'd52,10'd348};
ram[4482] = {-9'd49,10'd351};
ram[4483] = {-9'd46,10'd354};
ram[4484] = {-9'd43,10'd358};
ram[4485] = {-9'd40,10'd361};
ram[4486] = {-9'd37,10'd364};
ram[4487] = {-9'd33,10'd367};
ram[4488] = {-9'd30,10'd370};
ram[4489] = {-9'd27,10'd373};
ram[4490] = {-9'd24,10'd376};
ram[4491] = {-9'd21,10'd380};
ram[4492] = {-9'd18,10'd383};
ram[4493] = {-9'd15,10'd386};
ram[4494] = {-9'd11,10'd389};
ram[4495] = {-9'd8,10'd392};
ram[4496] = {-9'd5,10'd395};
ram[4497] = {-9'd2,10'd398};
ram[4498] = {9'd1,-10'd399};
ram[4499] = {9'd4,-10'd396};
ram[4500] = {9'd7,-10'd393};
ram[4501] = {9'd10,-10'd390};
ram[4502] = {9'd14,-10'd387};
ram[4503] = {9'd17,-10'd384};
ram[4504] = {9'd20,-10'd381};
ram[4505] = {9'd23,-10'd377};
ram[4506] = {9'd26,-10'd374};
ram[4507] = {9'd29,-10'd371};
ram[4508] = {9'd32,-10'd368};
ram[4509] = {9'd36,-10'd365};
ram[4510] = {9'd39,-10'd362};
ram[4511] = {9'd42,-10'd359};
ram[4512] = {9'd45,-10'd355};
ram[4513] = {9'd48,-10'd352};
ram[4514] = {9'd51,-10'd349};
ram[4515] = {9'd54,-10'd346};
ram[4516] = {9'd58,-10'd343};
ram[4517] = {9'd61,-10'd340};
ram[4518] = {9'd64,-10'd337};
ram[4519] = {9'd67,-10'd334};
ram[4520] = {9'd70,-10'd330};
ram[4521] = {9'd73,-10'd327};
ram[4522] = {9'd76,-10'd324};
ram[4523] = {9'd80,-10'd321};
ram[4524] = {9'd83,-10'd318};
ram[4525] = {9'd86,-10'd315};
ram[4526] = {9'd89,-10'd312};
ram[4527] = {9'd92,-10'd308};
ram[4528] = {9'd95,-10'd305};
ram[4529] = {9'd98,-10'd302};
ram[4530] = {-9'd99,-10'd299};
ram[4531] = {-9'd96,-10'd296};
ram[4532] = {-9'd92,-10'd293};
ram[4533] = {-9'd89,-10'd290};
ram[4534] = {-9'd86,-10'd286};
ram[4535] = {-9'd83,-10'd283};
ram[4536] = {-9'd80,-10'd280};
ram[4537] = {-9'd77,-10'd277};
ram[4538] = {-9'd74,-10'd274};
ram[4539] = {-9'd70,-10'd271};
ram[4540] = {-9'd67,-10'd268};
ram[4541] = {-9'd64,-10'd264};
ram[4542] = {-9'd61,-10'd261};
ram[4543] = {-9'd58,-10'd258};
ram[4544] = {-9'd55,-10'd255};
ram[4545] = {-9'd52,-10'd252};
ram[4546] = {-9'd48,-10'd249};
ram[4547] = {-9'd45,-10'd246};
ram[4548] = {-9'd42,-10'd242};
ram[4549] = {-9'd39,-10'd239};
ram[4550] = {-9'd36,-10'd236};
ram[4551] = {-9'd33,-10'd233};
ram[4552] = {-9'd30,-10'd230};
ram[4553] = {-9'd26,-10'd227};
ram[4554] = {-9'd23,-10'd224};
ram[4555] = {-9'd20,-10'd220};
ram[4556] = {-9'd17,-10'd217};
ram[4557] = {-9'd14,-10'd214};
ram[4558] = {-9'd11,-10'd211};
ram[4559] = {-9'd8,-10'd208};
ram[4560] = {-9'd4,-10'd205};
ram[4561] = {-9'd1,-10'd202};
ram[4562] = {9'd2,-10'd198};
ram[4563] = {9'd5,-10'd195};
ram[4564] = {9'd8,-10'd192};
ram[4565] = {9'd11,-10'd189};
ram[4566] = {9'd14,-10'd186};
ram[4567] = {9'd18,-10'd183};
ram[4568] = {9'd21,-10'd180};
ram[4569] = {9'd24,-10'd176};
ram[4570] = {9'd27,-10'd173};
ram[4571] = {9'd30,-10'd170};
ram[4572] = {9'd33,-10'd167};
ram[4573] = {9'd36,-10'd164};
ram[4574] = {9'd40,-10'd161};
ram[4575] = {9'd43,-10'd158};
ram[4576] = {9'd46,-10'd154};
ram[4577] = {9'd49,-10'd151};
ram[4578] = {9'd52,-10'd148};
ram[4579] = {9'd55,-10'd145};
ram[4580] = {9'd58,-10'd142};
ram[4581] = {9'd62,-10'd139};
ram[4582] = {9'd65,-10'd136};
ram[4583] = {9'd68,-10'd132};
ram[4584] = {9'd71,-10'd129};
ram[4585] = {9'd74,-10'd126};
ram[4586] = {9'd77,-10'd123};
ram[4587] = {9'd80,-10'd120};
ram[4588] = {9'd84,-10'd117};
ram[4589] = {9'd87,-10'd114};
ram[4590] = {9'd90,-10'd110};
ram[4591] = {9'd93,-10'd107};
ram[4592] = {9'd96,-10'd104};
ram[4593] = {9'd99,-10'd101};
ram[4594] = {-9'd98,-10'd98};
ram[4595] = {-9'd95,-10'd95};
ram[4596] = {-9'd92,-10'd92};
ram[4597] = {-9'd88,-10'd88};
ram[4598] = {-9'd85,-10'd85};
ram[4599] = {-9'd82,-10'd82};
ram[4600] = {-9'd79,-10'd79};
ram[4601] = {-9'd76,-10'd76};
ram[4602] = {-9'd73,-10'd73};
ram[4603] = {-9'd70,-10'd70};
ram[4604] = {-9'd66,-10'd66};
ram[4605] = {-9'd63,-10'd63};
ram[4606] = {-9'd60,-10'd60};
ram[4607] = {-9'd57,-10'd57};
ram[4608] = {-9'd57,-10'd57};
ram[4609] = {-9'd54,-10'd54};
ram[4610] = {-9'd51,-10'd51};
ram[4611] = {-9'd48,-10'd48};
ram[4612] = {-9'd44,-10'd44};
ram[4613] = {-9'd41,-10'd41};
ram[4614] = {-9'd38,-10'd38};
ram[4615] = {-9'd35,-10'd35};
ram[4616] = {-9'd32,-10'd32};
ram[4617] = {-9'd29,-10'd29};
ram[4618] = {-9'd26,-10'd26};
ram[4619] = {-9'd22,-10'd22};
ram[4620] = {-9'd19,-10'd19};
ram[4621] = {-9'd16,-10'd16};
ram[4622] = {-9'd13,-10'd13};
ram[4623] = {-9'd10,-10'd10};
ram[4624] = {-9'd7,-10'd7};
ram[4625] = {-9'd4,-10'd4};
ram[4626] = {9'd0,10'd0};
ram[4627] = {9'd3,10'd3};
ram[4628] = {9'd6,10'd6};
ram[4629] = {9'd9,10'd9};
ram[4630] = {9'd12,10'd12};
ram[4631] = {9'd15,10'd15};
ram[4632] = {9'd18,10'd18};
ram[4633] = {9'd21,10'd21};
ram[4634] = {9'd25,10'd25};
ram[4635] = {9'd28,10'd28};
ram[4636] = {9'd31,10'd31};
ram[4637] = {9'd34,10'd34};
ram[4638] = {9'd37,10'd37};
ram[4639] = {9'd40,10'd40};
ram[4640] = {9'd43,10'd43};
ram[4641] = {9'd47,10'd47};
ram[4642] = {9'd50,10'd50};
ram[4643] = {9'd53,10'd53};
ram[4644] = {9'd56,10'd56};
ram[4645] = {9'd59,10'd59};
ram[4646] = {9'd62,10'd62};
ram[4647] = {9'd65,10'd65};
ram[4648] = {9'd69,10'd69};
ram[4649] = {9'd72,10'd72};
ram[4650] = {9'd75,10'd75};
ram[4651] = {9'd78,10'd78};
ram[4652] = {9'd81,10'd81};
ram[4653] = {9'd84,10'd84};
ram[4654] = {9'd87,10'd87};
ram[4655] = {9'd91,10'd91};
ram[4656] = {9'd94,10'd94};
ram[4657] = {9'd97,10'd97};
ram[4658] = {-9'd100,10'd100};
ram[4659] = {-9'd97,10'd103};
ram[4660] = {-9'd94,10'd106};
ram[4661] = {-9'd91,10'd109};
ram[4662] = {-9'd88,10'd113};
ram[4663] = {-9'd85,10'd116};
ram[4664] = {-9'd81,10'd119};
ram[4665] = {-9'd78,10'd122};
ram[4666] = {-9'd75,10'd125};
ram[4667] = {-9'd72,10'd128};
ram[4668] = {-9'd69,10'd131};
ram[4669] = {-9'd66,10'd135};
ram[4670] = {-9'd63,10'd138};
ram[4671] = {-9'd59,10'd141};
ram[4672] = {-9'd56,10'd144};
ram[4673] = {-9'd53,10'd147};
ram[4674] = {-9'd50,10'd150};
ram[4675] = {-9'd47,10'd153};
ram[4676] = {-9'd44,10'd157};
ram[4677] = {-9'd41,10'd160};
ram[4678] = {-9'd37,10'd163};
ram[4679] = {-9'd34,10'd166};
ram[4680] = {-9'd31,10'd169};
ram[4681] = {-9'd28,10'd172};
ram[4682] = {-9'd25,10'd175};
ram[4683] = {-9'd22,10'd179};
ram[4684] = {-9'd19,10'd182};
ram[4685] = {-9'd15,10'd185};
ram[4686] = {-9'd12,10'd188};
ram[4687] = {-9'd9,10'd191};
ram[4688] = {-9'd6,10'd194};
ram[4689] = {-9'd3,10'd197};
ram[4690] = {9'd0,10'd201};
ram[4691] = {9'd3,10'd204};
ram[4692] = {9'd7,10'd207};
ram[4693] = {9'd10,10'd210};
ram[4694] = {9'd13,10'd213};
ram[4695] = {9'd16,10'd216};
ram[4696] = {9'd19,10'd219};
ram[4697] = {9'd22,10'd223};
ram[4698] = {9'd25,10'd226};
ram[4699] = {9'd29,10'd229};
ram[4700] = {9'd32,10'd232};
ram[4701] = {9'd35,10'd235};
ram[4702] = {9'd38,10'd238};
ram[4703] = {9'd41,10'd241};
ram[4704] = {9'd44,10'd245};
ram[4705] = {9'd47,10'd248};
ram[4706] = {9'd51,10'd251};
ram[4707] = {9'd54,10'd254};
ram[4708] = {9'd57,10'd257};
ram[4709] = {9'd60,10'd260};
ram[4710] = {9'd63,10'd263};
ram[4711] = {9'd66,10'd267};
ram[4712] = {9'd69,10'd270};
ram[4713] = {9'd73,10'd273};
ram[4714] = {9'd76,10'd276};
ram[4715] = {9'd79,10'd279};
ram[4716] = {9'd82,10'd282};
ram[4717] = {9'd85,10'd285};
ram[4718] = {9'd88,10'd289};
ram[4719] = {9'd91,10'd292};
ram[4720] = {9'd95,10'd295};
ram[4721] = {9'd98,10'd298};
ram[4722] = {-9'd99,10'd301};
ram[4723] = {-9'd96,10'd304};
ram[4724] = {-9'd93,10'd307};
ram[4725] = {-9'd90,10'd311};
ram[4726] = {-9'd87,10'd314};
ram[4727] = {-9'd84,10'd317};
ram[4728] = {-9'd81,10'd320};
ram[4729] = {-9'd77,10'd323};
ram[4730] = {-9'd74,10'd326};
ram[4731] = {-9'd71,10'd329};
ram[4732] = {-9'd68,10'd333};
ram[4733] = {-9'd65,10'd336};
ram[4734] = {-9'd62,10'd339};
ram[4735] = {-9'd59,10'd342};
ram[4736] = {-9'd59,10'd342};
ram[4737] = {-9'd55,10'd345};
ram[4738] = {-9'd52,10'd348};
ram[4739] = {-9'd49,10'd351};
ram[4740] = {-9'd46,10'd354};
ram[4741] = {-9'd43,10'd358};
ram[4742] = {-9'd40,10'd361};
ram[4743] = {-9'd37,10'd364};
ram[4744] = {-9'd33,10'd367};
ram[4745] = {-9'd30,10'd370};
ram[4746] = {-9'd27,10'd373};
ram[4747] = {-9'd24,10'd376};
ram[4748] = {-9'd21,10'd380};
ram[4749] = {-9'd18,10'd383};
ram[4750] = {-9'd15,10'd386};
ram[4751] = {-9'd11,10'd389};
ram[4752] = {-9'd8,10'd392};
ram[4753] = {-9'd5,10'd395};
ram[4754] = {-9'd2,10'd398};
ram[4755] = {9'd1,-10'd399};
ram[4756] = {9'd4,-10'd396};
ram[4757] = {9'd7,-10'd393};
ram[4758] = {9'd10,-10'd390};
ram[4759] = {9'd14,-10'd387};
ram[4760] = {9'd17,-10'd384};
ram[4761] = {9'd20,-10'd381};
ram[4762] = {9'd23,-10'd377};
ram[4763] = {9'd26,-10'd374};
ram[4764] = {9'd29,-10'd371};
ram[4765] = {9'd32,-10'd368};
ram[4766] = {9'd36,-10'd365};
ram[4767] = {9'd39,-10'd362};
ram[4768] = {9'd42,-10'd359};
ram[4769] = {9'd45,-10'd355};
ram[4770] = {9'd48,-10'd352};
ram[4771] = {9'd51,-10'd349};
ram[4772] = {9'd54,-10'd346};
ram[4773] = {9'd58,-10'd343};
ram[4774] = {9'd61,-10'd340};
ram[4775] = {9'd64,-10'd337};
ram[4776] = {9'd67,-10'd334};
ram[4777] = {9'd70,-10'd330};
ram[4778] = {9'd73,-10'd327};
ram[4779] = {9'd76,-10'd324};
ram[4780] = {9'd80,-10'd321};
ram[4781] = {9'd83,-10'd318};
ram[4782] = {9'd86,-10'd315};
ram[4783] = {9'd89,-10'd312};
ram[4784] = {9'd92,-10'd308};
ram[4785] = {9'd95,-10'd305};
ram[4786] = {9'd98,-10'd302};
ram[4787] = {-9'd99,-10'd299};
ram[4788] = {-9'd96,-10'd296};
ram[4789] = {-9'd92,-10'd293};
ram[4790] = {-9'd89,-10'd290};
ram[4791] = {-9'd86,-10'd286};
ram[4792] = {-9'd83,-10'd283};
ram[4793] = {-9'd80,-10'd280};
ram[4794] = {-9'd77,-10'd277};
ram[4795] = {-9'd74,-10'd274};
ram[4796] = {-9'd70,-10'd271};
ram[4797] = {-9'd67,-10'd268};
ram[4798] = {-9'd64,-10'd264};
ram[4799] = {-9'd61,-10'd261};
ram[4800] = {-9'd58,-10'd258};
ram[4801] = {-9'd55,-10'd255};
ram[4802] = {-9'd52,-10'd252};
ram[4803] = {-9'd48,-10'd249};
ram[4804] = {-9'd45,-10'd246};
ram[4805] = {-9'd42,-10'd242};
ram[4806] = {-9'd39,-10'd239};
ram[4807] = {-9'd36,-10'd236};
ram[4808] = {-9'd33,-10'd233};
ram[4809] = {-9'd30,-10'd230};
ram[4810] = {-9'd26,-10'd227};
ram[4811] = {-9'd23,-10'd224};
ram[4812] = {-9'd20,-10'd220};
ram[4813] = {-9'd17,-10'd217};
ram[4814] = {-9'd14,-10'd214};
ram[4815] = {-9'd11,-10'd211};
ram[4816] = {-9'd8,-10'd208};
ram[4817] = {-9'd4,-10'd205};
ram[4818] = {-9'd1,-10'd202};
ram[4819] = {9'd2,-10'd198};
ram[4820] = {9'd5,-10'd195};
ram[4821] = {9'd8,-10'd192};
ram[4822] = {9'd11,-10'd189};
ram[4823] = {9'd14,-10'd186};
ram[4824] = {9'd18,-10'd183};
ram[4825] = {9'd21,-10'd180};
ram[4826] = {9'd24,-10'd176};
ram[4827] = {9'd27,-10'd173};
ram[4828] = {9'd30,-10'd170};
ram[4829] = {9'd33,-10'd167};
ram[4830] = {9'd36,-10'd164};
ram[4831] = {9'd40,-10'd161};
ram[4832] = {9'd43,-10'd158};
ram[4833] = {9'd46,-10'd154};
ram[4834] = {9'd49,-10'd151};
ram[4835] = {9'd52,-10'd148};
ram[4836] = {9'd55,-10'd145};
ram[4837] = {9'd58,-10'd142};
ram[4838] = {9'd62,-10'd139};
ram[4839] = {9'd65,-10'd136};
ram[4840] = {9'd68,-10'd132};
ram[4841] = {9'd71,-10'd129};
ram[4842] = {9'd74,-10'd126};
ram[4843] = {9'd77,-10'd123};
ram[4844] = {9'd80,-10'd120};
ram[4845] = {9'd84,-10'd117};
ram[4846] = {9'd87,-10'd114};
ram[4847] = {9'd90,-10'd110};
ram[4848] = {9'd93,-10'd107};
ram[4849] = {9'd96,-10'd104};
ram[4850] = {9'd99,-10'd101};
ram[4851] = {-9'd98,-10'd98};
ram[4852] = {-9'd95,-10'd95};
ram[4853] = {-9'd92,-10'd92};
ram[4854] = {-9'd88,-10'd88};
ram[4855] = {-9'd85,-10'd85};
ram[4856] = {-9'd82,-10'd82};
ram[4857] = {-9'd79,-10'd79};
ram[4858] = {-9'd76,-10'd76};
ram[4859] = {-9'd73,-10'd73};
ram[4860] = {-9'd70,-10'd70};
ram[4861] = {-9'd66,-10'd66};
ram[4862] = {-9'd63,-10'd63};
ram[4863] = {-9'd60,-10'd60};
ram[4864] = {-9'd60,-10'd60};
ram[4865] = {-9'd57,-10'd57};
ram[4866] = {-9'd54,-10'd54};
ram[4867] = {-9'd51,-10'd51};
ram[4868] = {-9'd48,-10'd48};
ram[4869] = {-9'd44,-10'd44};
ram[4870] = {-9'd41,-10'd41};
ram[4871] = {-9'd38,-10'd38};
ram[4872] = {-9'd35,-10'd35};
ram[4873] = {-9'd32,-10'd32};
ram[4874] = {-9'd29,-10'd29};
ram[4875] = {-9'd26,-10'd26};
ram[4876] = {-9'd22,-10'd22};
ram[4877] = {-9'd19,-10'd19};
ram[4878] = {-9'd16,-10'd16};
ram[4879] = {-9'd13,-10'd13};
ram[4880] = {-9'd10,-10'd10};
ram[4881] = {-9'd7,-10'd7};
ram[4882] = {-9'd4,-10'd4};
ram[4883] = {9'd0,10'd0};
ram[4884] = {9'd3,10'd3};
ram[4885] = {9'd6,10'd6};
ram[4886] = {9'd9,10'd9};
ram[4887] = {9'd12,10'd12};
ram[4888] = {9'd15,10'd15};
ram[4889] = {9'd18,10'd18};
ram[4890] = {9'd21,10'd21};
ram[4891] = {9'd25,10'd25};
ram[4892] = {9'd28,10'd28};
ram[4893] = {9'd31,10'd31};
ram[4894] = {9'd34,10'd34};
ram[4895] = {9'd37,10'd37};
ram[4896] = {9'd40,10'd40};
ram[4897] = {9'd43,10'd43};
ram[4898] = {9'd47,10'd47};
ram[4899] = {9'd50,10'd50};
ram[4900] = {9'd53,10'd53};
ram[4901] = {9'd56,10'd56};
ram[4902] = {9'd59,10'd59};
ram[4903] = {9'd62,10'd62};
ram[4904] = {9'd65,10'd65};
ram[4905] = {9'd69,10'd69};
ram[4906] = {9'd72,10'd72};
ram[4907] = {9'd75,10'd75};
ram[4908] = {9'd78,10'd78};
ram[4909] = {9'd81,10'd81};
ram[4910] = {9'd84,10'd84};
ram[4911] = {9'd87,10'd87};
ram[4912] = {9'd91,10'd91};
ram[4913] = {9'd94,10'd94};
ram[4914] = {9'd97,10'd97};
ram[4915] = {-9'd100,10'd100};
ram[4916] = {-9'd97,10'd103};
ram[4917] = {-9'd94,10'd106};
ram[4918] = {-9'd91,10'd109};
ram[4919] = {-9'd88,10'd113};
ram[4920] = {-9'd85,10'd116};
ram[4921] = {-9'd81,10'd119};
ram[4922] = {-9'd78,10'd122};
ram[4923] = {-9'd75,10'd125};
ram[4924] = {-9'd72,10'd128};
ram[4925] = {-9'd69,10'd131};
ram[4926] = {-9'd66,10'd135};
ram[4927] = {-9'd63,10'd138};
ram[4928] = {-9'd59,10'd141};
ram[4929] = {-9'd56,10'd144};
ram[4930] = {-9'd53,10'd147};
ram[4931] = {-9'd50,10'd150};
ram[4932] = {-9'd47,10'd153};
ram[4933] = {-9'd44,10'd157};
ram[4934] = {-9'd41,10'd160};
ram[4935] = {-9'd37,10'd163};
ram[4936] = {-9'd34,10'd166};
ram[4937] = {-9'd31,10'd169};
ram[4938] = {-9'd28,10'd172};
ram[4939] = {-9'd25,10'd175};
ram[4940] = {-9'd22,10'd179};
ram[4941] = {-9'd19,10'd182};
ram[4942] = {-9'd15,10'd185};
ram[4943] = {-9'd12,10'd188};
ram[4944] = {-9'd9,10'd191};
ram[4945] = {-9'd6,10'd194};
ram[4946] = {-9'd3,10'd197};
ram[4947] = {9'd0,10'd201};
ram[4948] = {9'd3,10'd204};
ram[4949] = {9'd7,10'd207};
ram[4950] = {9'd10,10'd210};
ram[4951] = {9'd13,10'd213};
ram[4952] = {9'd16,10'd216};
ram[4953] = {9'd19,10'd219};
ram[4954] = {9'd22,10'd223};
ram[4955] = {9'd25,10'd226};
ram[4956] = {9'd29,10'd229};
ram[4957] = {9'd32,10'd232};
ram[4958] = {9'd35,10'd235};
ram[4959] = {9'd38,10'd238};
ram[4960] = {9'd41,10'd241};
ram[4961] = {9'd44,10'd245};
ram[4962] = {9'd47,10'd248};
ram[4963] = {9'd51,10'd251};
ram[4964] = {9'd54,10'd254};
ram[4965] = {9'd57,10'd257};
ram[4966] = {9'd60,10'd260};
ram[4967] = {9'd63,10'd263};
ram[4968] = {9'd66,10'd267};
ram[4969] = {9'd69,10'd270};
ram[4970] = {9'd73,10'd273};
ram[4971] = {9'd76,10'd276};
ram[4972] = {9'd79,10'd279};
ram[4973] = {9'd82,10'd282};
ram[4974] = {9'd85,10'd285};
ram[4975] = {9'd88,10'd289};
ram[4976] = {9'd91,10'd292};
ram[4977] = {9'd95,10'd295};
ram[4978] = {9'd98,10'd298};
ram[4979] = {-9'd99,10'd301};
ram[4980] = {-9'd96,10'd304};
ram[4981] = {-9'd93,10'd307};
ram[4982] = {-9'd90,10'd311};
ram[4983] = {-9'd87,10'd314};
ram[4984] = {-9'd84,10'd317};
ram[4985] = {-9'd81,10'd320};
ram[4986] = {-9'd77,10'd323};
ram[4987] = {-9'd74,10'd326};
ram[4988] = {-9'd71,10'd329};
ram[4989] = {-9'd68,10'd333};
ram[4990] = {-9'd65,10'd336};
ram[4991] = {-9'd62,10'd339};
ram[4992] = {-9'd62,10'd339};
ram[4993] = {-9'd59,10'd342};
ram[4994] = {-9'd55,10'd345};
ram[4995] = {-9'd52,10'd348};
ram[4996] = {-9'd49,10'd351};
ram[4997] = {-9'd46,10'd354};
ram[4998] = {-9'd43,10'd358};
ram[4999] = {-9'd40,10'd361};
ram[5000] = {-9'd37,10'd364};
ram[5001] = {-9'd33,10'd367};
ram[5002] = {-9'd30,10'd370};
ram[5003] = {-9'd27,10'd373};
ram[5004] = {-9'd24,10'd376};
ram[5005] = {-9'd21,10'd380};
ram[5006] = {-9'd18,10'd383};
ram[5007] = {-9'd15,10'd386};
ram[5008] = {-9'd11,10'd389};
ram[5009] = {-9'd8,10'd392};
ram[5010] = {-9'd5,10'd395};
ram[5011] = {-9'd2,10'd398};
ram[5012] = {9'd1,-10'd399};
ram[5013] = {9'd4,-10'd396};
ram[5014] = {9'd7,-10'd393};
ram[5015] = {9'd10,-10'd390};
ram[5016] = {9'd14,-10'd387};
ram[5017] = {9'd17,-10'd384};
ram[5018] = {9'd20,-10'd381};
ram[5019] = {9'd23,-10'd377};
ram[5020] = {9'd26,-10'd374};
ram[5021] = {9'd29,-10'd371};
ram[5022] = {9'd32,-10'd368};
ram[5023] = {9'd36,-10'd365};
ram[5024] = {9'd39,-10'd362};
ram[5025] = {9'd42,-10'd359};
ram[5026] = {9'd45,-10'd355};
ram[5027] = {9'd48,-10'd352};
ram[5028] = {9'd51,-10'd349};
ram[5029] = {9'd54,-10'd346};
ram[5030] = {9'd58,-10'd343};
ram[5031] = {9'd61,-10'd340};
ram[5032] = {9'd64,-10'd337};
ram[5033] = {9'd67,-10'd334};
ram[5034] = {9'd70,-10'd330};
ram[5035] = {9'd73,-10'd327};
ram[5036] = {9'd76,-10'd324};
ram[5037] = {9'd80,-10'd321};
ram[5038] = {9'd83,-10'd318};
ram[5039] = {9'd86,-10'd315};
ram[5040] = {9'd89,-10'd312};
ram[5041] = {9'd92,-10'd308};
ram[5042] = {9'd95,-10'd305};
ram[5043] = {9'd98,-10'd302};
ram[5044] = {-9'd99,-10'd299};
ram[5045] = {-9'd96,-10'd296};
ram[5046] = {-9'd92,-10'd293};
ram[5047] = {-9'd89,-10'd290};
ram[5048] = {-9'd86,-10'd286};
ram[5049] = {-9'd83,-10'd283};
ram[5050] = {-9'd80,-10'd280};
ram[5051] = {-9'd77,-10'd277};
ram[5052] = {-9'd74,-10'd274};
ram[5053] = {-9'd70,-10'd271};
ram[5054] = {-9'd67,-10'd268};
ram[5055] = {-9'd64,-10'd264};
ram[5056] = {-9'd61,-10'd261};
ram[5057] = {-9'd58,-10'd258};
ram[5058] = {-9'd55,-10'd255};
ram[5059] = {-9'd52,-10'd252};
ram[5060] = {-9'd48,-10'd249};
ram[5061] = {-9'd45,-10'd246};
ram[5062] = {-9'd42,-10'd242};
ram[5063] = {-9'd39,-10'd239};
ram[5064] = {-9'd36,-10'd236};
ram[5065] = {-9'd33,-10'd233};
ram[5066] = {-9'd30,-10'd230};
ram[5067] = {-9'd26,-10'd227};
ram[5068] = {-9'd23,-10'd224};
ram[5069] = {-9'd20,-10'd220};
ram[5070] = {-9'd17,-10'd217};
ram[5071] = {-9'd14,-10'd214};
ram[5072] = {-9'd11,-10'd211};
ram[5073] = {-9'd8,-10'd208};
ram[5074] = {-9'd4,-10'd205};
ram[5075] = {-9'd1,-10'd202};
ram[5076] = {9'd2,-10'd198};
ram[5077] = {9'd5,-10'd195};
ram[5078] = {9'd8,-10'd192};
ram[5079] = {9'd11,-10'd189};
ram[5080] = {9'd14,-10'd186};
ram[5081] = {9'd18,-10'd183};
ram[5082] = {9'd21,-10'd180};
ram[5083] = {9'd24,-10'd176};
ram[5084] = {9'd27,-10'd173};
ram[5085] = {9'd30,-10'd170};
ram[5086] = {9'd33,-10'd167};
ram[5087] = {9'd36,-10'd164};
ram[5088] = {9'd40,-10'd161};
ram[5089] = {9'd43,-10'd158};
ram[5090] = {9'd46,-10'd154};
ram[5091] = {9'd49,-10'd151};
ram[5092] = {9'd52,-10'd148};
ram[5093] = {9'd55,-10'd145};
ram[5094] = {9'd58,-10'd142};
ram[5095] = {9'd62,-10'd139};
ram[5096] = {9'd65,-10'd136};
ram[5097] = {9'd68,-10'd132};
ram[5098] = {9'd71,-10'd129};
ram[5099] = {9'd74,-10'd126};
ram[5100] = {9'd77,-10'd123};
ram[5101] = {9'd80,-10'd120};
ram[5102] = {9'd84,-10'd117};
ram[5103] = {9'd87,-10'd114};
ram[5104] = {9'd90,-10'd110};
ram[5105] = {9'd93,-10'd107};
ram[5106] = {9'd96,-10'd104};
ram[5107] = {9'd99,-10'd101};
ram[5108] = {-9'd98,-10'd98};
ram[5109] = {-9'd95,-10'd95};
ram[5110] = {-9'd92,-10'd92};
ram[5111] = {-9'd88,-10'd88};
ram[5112] = {-9'd85,-10'd85};
ram[5113] = {-9'd82,-10'd82};
ram[5114] = {-9'd79,-10'd79};
ram[5115] = {-9'd76,-10'd76};
ram[5116] = {-9'd73,-10'd73};
ram[5117] = {-9'd70,-10'd70};
ram[5118] = {-9'd66,-10'd66};
ram[5119] = {-9'd63,-10'd63};
ram[5120] = {-9'd63,-10'd63};
ram[5121] = {-9'd60,-10'd60};
ram[5122] = {-9'd57,-10'd57};
ram[5123] = {-9'd54,-10'd54};
ram[5124] = {-9'd51,-10'd51};
ram[5125] = {-9'd48,-10'd48};
ram[5126] = {-9'd44,-10'd44};
ram[5127] = {-9'd41,-10'd41};
ram[5128] = {-9'd38,-10'd38};
ram[5129] = {-9'd35,-10'd35};
ram[5130] = {-9'd32,-10'd32};
ram[5131] = {-9'd29,-10'd29};
ram[5132] = {-9'd26,-10'd26};
ram[5133] = {-9'd22,-10'd22};
ram[5134] = {-9'd19,-10'd19};
ram[5135] = {-9'd16,-10'd16};
ram[5136] = {-9'd13,-10'd13};
ram[5137] = {-9'd10,-10'd10};
ram[5138] = {-9'd7,-10'd7};
ram[5139] = {-9'd4,-10'd4};
ram[5140] = {9'd0,10'd0};
ram[5141] = {9'd3,10'd3};
ram[5142] = {9'd6,10'd6};
ram[5143] = {9'd9,10'd9};
ram[5144] = {9'd12,10'd12};
ram[5145] = {9'd15,10'd15};
ram[5146] = {9'd18,10'd18};
ram[5147] = {9'd21,10'd21};
ram[5148] = {9'd25,10'd25};
ram[5149] = {9'd28,10'd28};
ram[5150] = {9'd31,10'd31};
ram[5151] = {9'd34,10'd34};
ram[5152] = {9'd37,10'd37};
ram[5153] = {9'd40,10'd40};
ram[5154] = {9'd43,10'd43};
ram[5155] = {9'd47,10'd47};
ram[5156] = {9'd50,10'd50};
ram[5157] = {9'd53,10'd53};
ram[5158] = {9'd56,10'd56};
ram[5159] = {9'd59,10'd59};
ram[5160] = {9'd62,10'd62};
ram[5161] = {9'd65,10'd65};
ram[5162] = {9'd69,10'd69};
ram[5163] = {9'd72,10'd72};
ram[5164] = {9'd75,10'd75};
ram[5165] = {9'd78,10'd78};
ram[5166] = {9'd81,10'd81};
ram[5167] = {9'd84,10'd84};
ram[5168] = {9'd87,10'd87};
ram[5169] = {9'd91,10'd91};
ram[5170] = {9'd94,10'd94};
ram[5171] = {9'd97,10'd97};
ram[5172] = {-9'd100,10'd100};
ram[5173] = {-9'd97,10'd103};
ram[5174] = {-9'd94,10'd106};
ram[5175] = {-9'd91,10'd109};
ram[5176] = {-9'd88,10'd113};
ram[5177] = {-9'd85,10'd116};
ram[5178] = {-9'd81,10'd119};
ram[5179] = {-9'd78,10'd122};
ram[5180] = {-9'd75,10'd125};
ram[5181] = {-9'd72,10'd128};
ram[5182] = {-9'd69,10'd131};
ram[5183] = {-9'd66,10'd135};
ram[5184] = {-9'd63,10'd138};
ram[5185] = {-9'd59,10'd141};
ram[5186] = {-9'd56,10'd144};
ram[5187] = {-9'd53,10'd147};
ram[5188] = {-9'd50,10'd150};
ram[5189] = {-9'd47,10'd153};
ram[5190] = {-9'd44,10'd157};
ram[5191] = {-9'd41,10'd160};
ram[5192] = {-9'd37,10'd163};
ram[5193] = {-9'd34,10'd166};
ram[5194] = {-9'd31,10'd169};
ram[5195] = {-9'd28,10'd172};
ram[5196] = {-9'd25,10'd175};
ram[5197] = {-9'd22,10'd179};
ram[5198] = {-9'd19,10'd182};
ram[5199] = {-9'd15,10'd185};
ram[5200] = {-9'd12,10'd188};
ram[5201] = {-9'd9,10'd191};
ram[5202] = {-9'd6,10'd194};
ram[5203] = {-9'd3,10'd197};
ram[5204] = {9'd0,10'd201};
ram[5205] = {9'd3,10'd204};
ram[5206] = {9'd7,10'd207};
ram[5207] = {9'd10,10'd210};
ram[5208] = {9'd13,10'd213};
ram[5209] = {9'd16,10'd216};
ram[5210] = {9'd19,10'd219};
ram[5211] = {9'd22,10'd223};
ram[5212] = {9'd25,10'd226};
ram[5213] = {9'd29,10'd229};
ram[5214] = {9'd32,10'd232};
ram[5215] = {9'd35,10'd235};
ram[5216] = {9'd38,10'd238};
ram[5217] = {9'd41,10'd241};
ram[5218] = {9'd44,10'd245};
ram[5219] = {9'd47,10'd248};
ram[5220] = {9'd51,10'd251};
ram[5221] = {9'd54,10'd254};
ram[5222] = {9'd57,10'd257};
ram[5223] = {9'd60,10'd260};
ram[5224] = {9'd63,10'd263};
ram[5225] = {9'd66,10'd267};
ram[5226] = {9'd69,10'd270};
ram[5227] = {9'd73,10'd273};
ram[5228] = {9'd76,10'd276};
ram[5229] = {9'd79,10'd279};
ram[5230] = {9'd82,10'd282};
ram[5231] = {9'd85,10'd285};
ram[5232] = {9'd88,10'd289};
ram[5233] = {9'd91,10'd292};
ram[5234] = {9'd95,10'd295};
ram[5235] = {9'd98,10'd298};
ram[5236] = {-9'd99,10'd301};
ram[5237] = {-9'd96,10'd304};
ram[5238] = {-9'd93,10'd307};
ram[5239] = {-9'd90,10'd311};
ram[5240] = {-9'd87,10'd314};
ram[5241] = {-9'd84,10'd317};
ram[5242] = {-9'd81,10'd320};
ram[5243] = {-9'd77,10'd323};
ram[5244] = {-9'd74,10'd326};
ram[5245] = {-9'd71,10'd329};
ram[5246] = {-9'd68,10'd333};
ram[5247] = {-9'd65,10'd336};
ram[5248] = {-9'd65,10'd336};
ram[5249] = {-9'd62,10'd339};
ram[5250] = {-9'd59,10'd342};
ram[5251] = {-9'd55,10'd345};
ram[5252] = {-9'd52,10'd348};
ram[5253] = {-9'd49,10'd351};
ram[5254] = {-9'd46,10'd354};
ram[5255] = {-9'd43,10'd358};
ram[5256] = {-9'd40,10'd361};
ram[5257] = {-9'd37,10'd364};
ram[5258] = {-9'd33,10'd367};
ram[5259] = {-9'd30,10'd370};
ram[5260] = {-9'd27,10'd373};
ram[5261] = {-9'd24,10'd376};
ram[5262] = {-9'd21,10'd380};
ram[5263] = {-9'd18,10'd383};
ram[5264] = {-9'd15,10'd386};
ram[5265] = {-9'd11,10'd389};
ram[5266] = {-9'd8,10'd392};
ram[5267] = {-9'd5,10'd395};
ram[5268] = {-9'd2,10'd398};
ram[5269] = {9'd1,-10'd399};
ram[5270] = {9'd4,-10'd396};
ram[5271] = {9'd7,-10'd393};
ram[5272] = {9'd10,-10'd390};
ram[5273] = {9'd14,-10'd387};
ram[5274] = {9'd17,-10'd384};
ram[5275] = {9'd20,-10'd381};
ram[5276] = {9'd23,-10'd377};
ram[5277] = {9'd26,-10'd374};
ram[5278] = {9'd29,-10'd371};
ram[5279] = {9'd32,-10'd368};
ram[5280] = {9'd36,-10'd365};
ram[5281] = {9'd39,-10'd362};
ram[5282] = {9'd42,-10'd359};
ram[5283] = {9'd45,-10'd355};
ram[5284] = {9'd48,-10'd352};
ram[5285] = {9'd51,-10'd349};
ram[5286] = {9'd54,-10'd346};
ram[5287] = {9'd58,-10'd343};
ram[5288] = {9'd61,-10'd340};
ram[5289] = {9'd64,-10'd337};
ram[5290] = {9'd67,-10'd334};
ram[5291] = {9'd70,-10'd330};
ram[5292] = {9'd73,-10'd327};
ram[5293] = {9'd76,-10'd324};
ram[5294] = {9'd80,-10'd321};
ram[5295] = {9'd83,-10'd318};
ram[5296] = {9'd86,-10'd315};
ram[5297] = {9'd89,-10'd312};
ram[5298] = {9'd92,-10'd308};
ram[5299] = {9'd95,-10'd305};
ram[5300] = {9'd98,-10'd302};
ram[5301] = {-9'd99,-10'd299};
ram[5302] = {-9'd96,-10'd296};
ram[5303] = {-9'd92,-10'd293};
ram[5304] = {-9'd89,-10'd290};
ram[5305] = {-9'd86,-10'd286};
ram[5306] = {-9'd83,-10'd283};
ram[5307] = {-9'd80,-10'd280};
ram[5308] = {-9'd77,-10'd277};
ram[5309] = {-9'd74,-10'd274};
ram[5310] = {-9'd70,-10'd271};
ram[5311] = {-9'd67,-10'd268};
ram[5312] = {-9'd64,-10'd264};
ram[5313] = {-9'd61,-10'd261};
ram[5314] = {-9'd58,-10'd258};
ram[5315] = {-9'd55,-10'd255};
ram[5316] = {-9'd52,-10'd252};
ram[5317] = {-9'd48,-10'd249};
ram[5318] = {-9'd45,-10'd246};
ram[5319] = {-9'd42,-10'd242};
ram[5320] = {-9'd39,-10'd239};
ram[5321] = {-9'd36,-10'd236};
ram[5322] = {-9'd33,-10'd233};
ram[5323] = {-9'd30,-10'd230};
ram[5324] = {-9'd26,-10'd227};
ram[5325] = {-9'd23,-10'd224};
ram[5326] = {-9'd20,-10'd220};
ram[5327] = {-9'd17,-10'd217};
ram[5328] = {-9'd14,-10'd214};
ram[5329] = {-9'd11,-10'd211};
ram[5330] = {-9'd8,-10'd208};
ram[5331] = {-9'd4,-10'd205};
ram[5332] = {-9'd1,-10'd202};
ram[5333] = {9'd2,-10'd198};
ram[5334] = {9'd5,-10'd195};
ram[5335] = {9'd8,-10'd192};
ram[5336] = {9'd11,-10'd189};
ram[5337] = {9'd14,-10'd186};
ram[5338] = {9'd18,-10'd183};
ram[5339] = {9'd21,-10'd180};
ram[5340] = {9'd24,-10'd176};
ram[5341] = {9'd27,-10'd173};
ram[5342] = {9'd30,-10'd170};
ram[5343] = {9'd33,-10'd167};
ram[5344] = {9'd36,-10'd164};
ram[5345] = {9'd40,-10'd161};
ram[5346] = {9'd43,-10'd158};
ram[5347] = {9'd46,-10'd154};
ram[5348] = {9'd49,-10'd151};
ram[5349] = {9'd52,-10'd148};
ram[5350] = {9'd55,-10'd145};
ram[5351] = {9'd58,-10'd142};
ram[5352] = {9'd62,-10'd139};
ram[5353] = {9'd65,-10'd136};
ram[5354] = {9'd68,-10'd132};
ram[5355] = {9'd71,-10'd129};
ram[5356] = {9'd74,-10'd126};
ram[5357] = {9'd77,-10'd123};
ram[5358] = {9'd80,-10'd120};
ram[5359] = {9'd84,-10'd117};
ram[5360] = {9'd87,-10'd114};
ram[5361] = {9'd90,-10'd110};
ram[5362] = {9'd93,-10'd107};
ram[5363] = {9'd96,-10'd104};
ram[5364] = {9'd99,-10'd101};
ram[5365] = {-9'd98,-10'd98};
ram[5366] = {-9'd95,-10'd95};
ram[5367] = {-9'd92,-10'd92};
ram[5368] = {-9'd88,-10'd88};
ram[5369] = {-9'd85,-10'd85};
ram[5370] = {-9'd82,-10'd82};
ram[5371] = {-9'd79,-10'd79};
ram[5372] = {-9'd76,-10'd76};
ram[5373] = {-9'd73,-10'd73};
ram[5374] = {-9'd70,-10'd70};
ram[5375] = {-9'd66,-10'd66};
ram[5376] = {-9'd66,-10'd66};
ram[5377] = {-9'd63,-10'd63};
ram[5378] = {-9'd60,-10'd60};
ram[5379] = {-9'd57,-10'd57};
ram[5380] = {-9'd54,-10'd54};
ram[5381] = {-9'd51,-10'd51};
ram[5382] = {-9'd48,-10'd48};
ram[5383] = {-9'd44,-10'd44};
ram[5384] = {-9'd41,-10'd41};
ram[5385] = {-9'd38,-10'd38};
ram[5386] = {-9'd35,-10'd35};
ram[5387] = {-9'd32,-10'd32};
ram[5388] = {-9'd29,-10'd29};
ram[5389] = {-9'd26,-10'd26};
ram[5390] = {-9'd22,-10'd22};
ram[5391] = {-9'd19,-10'd19};
ram[5392] = {-9'd16,-10'd16};
ram[5393] = {-9'd13,-10'd13};
ram[5394] = {-9'd10,-10'd10};
ram[5395] = {-9'd7,-10'd7};
ram[5396] = {-9'd4,-10'd4};
ram[5397] = {9'd0,10'd0};
ram[5398] = {9'd3,10'd3};
ram[5399] = {9'd6,10'd6};
ram[5400] = {9'd9,10'd9};
ram[5401] = {9'd12,10'd12};
ram[5402] = {9'd15,10'd15};
ram[5403] = {9'd18,10'd18};
ram[5404] = {9'd21,10'd21};
ram[5405] = {9'd25,10'd25};
ram[5406] = {9'd28,10'd28};
ram[5407] = {9'd31,10'd31};
ram[5408] = {9'd34,10'd34};
ram[5409] = {9'd37,10'd37};
ram[5410] = {9'd40,10'd40};
ram[5411] = {9'd43,10'd43};
ram[5412] = {9'd47,10'd47};
ram[5413] = {9'd50,10'd50};
ram[5414] = {9'd53,10'd53};
ram[5415] = {9'd56,10'd56};
ram[5416] = {9'd59,10'd59};
ram[5417] = {9'd62,10'd62};
ram[5418] = {9'd65,10'd65};
ram[5419] = {9'd69,10'd69};
ram[5420] = {9'd72,10'd72};
ram[5421] = {9'd75,10'd75};
ram[5422] = {9'd78,10'd78};
ram[5423] = {9'd81,10'd81};
ram[5424] = {9'd84,10'd84};
ram[5425] = {9'd87,10'd87};
ram[5426] = {9'd91,10'd91};
ram[5427] = {9'd94,10'd94};
ram[5428] = {9'd97,10'd97};
ram[5429] = {-9'd100,10'd100};
ram[5430] = {-9'd97,10'd103};
ram[5431] = {-9'd94,10'd106};
ram[5432] = {-9'd91,10'd109};
ram[5433] = {-9'd88,10'd113};
ram[5434] = {-9'd85,10'd116};
ram[5435] = {-9'd81,10'd119};
ram[5436] = {-9'd78,10'd122};
ram[5437] = {-9'd75,10'd125};
ram[5438] = {-9'd72,10'd128};
ram[5439] = {-9'd69,10'd131};
ram[5440] = {-9'd66,10'd135};
ram[5441] = {-9'd63,10'd138};
ram[5442] = {-9'd59,10'd141};
ram[5443] = {-9'd56,10'd144};
ram[5444] = {-9'd53,10'd147};
ram[5445] = {-9'd50,10'd150};
ram[5446] = {-9'd47,10'd153};
ram[5447] = {-9'd44,10'd157};
ram[5448] = {-9'd41,10'd160};
ram[5449] = {-9'd37,10'd163};
ram[5450] = {-9'd34,10'd166};
ram[5451] = {-9'd31,10'd169};
ram[5452] = {-9'd28,10'd172};
ram[5453] = {-9'd25,10'd175};
ram[5454] = {-9'd22,10'd179};
ram[5455] = {-9'd19,10'd182};
ram[5456] = {-9'd15,10'd185};
ram[5457] = {-9'd12,10'd188};
ram[5458] = {-9'd9,10'd191};
ram[5459] = {-9'd6,10'd194};
ram[5460] = {-9'd3,10'd197};
ram[5461] = {9'd0,10'd201};
ram[5462] = {9'd3,10'd204};
ram[5463] = {9'd7,10'd207};
ram[5464] = {9'd10,10'd210};
ram[5465] = {9'd13,10'd213};
ram[5466] = {9'd16,10'd216};
ram[5467] = {9'd19,10'd219};
ram[5468] = {9'd22,10'd223};
ram[5469] = {9'd25,10'd226};
ram[5470] = {9'd29,10'd229};
ram[5471] = {9'd32,10'd232};
ram[5472] = {9'd35,10'd235};
ram[5473] = {9'd38,10'd238};
ram[5474] = {9'd41,10'd241};
ram[5475] = {9'd44,10'd245};
ram[5476] = {9'd47,10'd248};
ram[5477] = {9'd51,10'd251};
ram[5478] = {9'd54,10'd254};
ram[5479] = {9'd57,10'd257};
ram[5480] = {9'd60,10'd260};
ram[5481] = {9'd63,10'd263};
ram[5482] = {9'd66,10'd267};
ram[5483] = {9'd69,10'd270};
ram[5484] = {9'd73,10'd273};
ram[5485] = {9'd76,10'd276};
ram[5486] = {9'd79,10'd279};
ram[5487] = {9'd82,10'd282};
ram[5488] = {9'd85,10'd285};
ram[5489] = {9'd88,10'd289};
ram[5490] = {9'd91,10'd292};
ram[5491] = {9'd95,10'd295};
ram[5492] = {9'd98,10'd298};
ram[5493] = {-9'd99,10'd301};
ram[5494] = {-9'd96,10'd304};
ram[5495] = {-9'd93,10'd307};
ram[5496] = {-9'd90,10'd311};
ram[5497] = {-9'd87,10'd314};
ram[5498] = {-9'd84,10'd317};
ram[5499] = {-9'd81,10'd320};
ram[5500] = {-9'd77,10'd323};
ram[5501] = {-9'd74,10'd326};
ram[5502] = {-9'd71,10'd329};
ram[5503] = {-9'd68,10'd333};
ram[5504] = {-9'd68,10'd333};
ram[5505] = {-9'd65,10'd336};
ram[5506] = {-9'd62,10'd339};
ram[5507] = {-9'd59,10'd342};
ram[5508] = {-9'd55,10'd345};
ram[5509] = {-9'd52,10'd348};
ram[5510] = {-9'd49,10'd351};
ram[5511] = {-9'd46,10'd354};
ram[5512] = {-9'd43,10'd358};
ram[5513] = {-9'd40,10'd361};
ram[5514] = {-9'd37,10'd364};
ram[5515] = {-9'd33,10'd367};
ram[5516] = {-9'd30,10'd370};
ram[5517] = {-9'd27,10'd373};
ram[5518] = {-9'd24,10'd376};
ram[5519] = {-9'd21,10'd380};
ram[5520] = {-9'd18,10'd383};
ram[5521] = {-9'd15,10'd386};
ram[5522] = {-9'd11,10'd389};
ram[5523] = {-9'd8,10'd392};
ram[5524] = {-9'd5,10'd395};
ram[5525] = {-9'd2,10'd398};
ram[5526] = {9'd1,-10'd399};
ram[5527] = {9'd4,-10'd396};
ram[5528] = {9'd7,-10'd393};
ram[5529] = {9'd10,-10'd390};
ram[5530] = {9'd14,-10'd387};
ram[5531] = {9'd17,-10'd384};
ram[5532] = {9'd20,-10'd381};
ram[5533] = {9'd23,-10'd377};
ram[5534] = {9'd26,-10'd374};
ram[5535] = {9'd29,-10'd371};
ram[5536] = {9'd32,-10'd368};
ram[5537] = {9'd36,-10'd365};
ram[5538] = {9'd39,-10'd362};
ram[5539] = {9'd42,-10'd359};
ram[5540] = {9'd45,-10'd355};
ram[5541] = {9'd48,-10'd352};
ram[5542] = {9'd51,-10'd349};
ram[5543] = {9'd54,-10'd346};
ram[5544] = {9'd58,-10'd343};
ram[5545] = {9'd61,-10'd340};
ram[5546] = {9'd64,-10'd337};
ram[5547] = {9'd67,-10'd334};
ram[5548] = {9'd70,-10'd330};
ram[5549] = {9'd73,-10'd327};
ram[5550] = {9'd76,-10'd324};
ram[5551] = {9'd80,-10'd321};
ram[5552] = {9'd83,-10'd318};
ram[5553] = {9'd86,-10'd315};
ram[5554] = {9'd89,-10'd312};
ram[5555] = {9'd92,-10'd308};
ram[5556] = {9'd95,-10'd305};
ram[5557] = {9'd98,-10'd302};
ram[5558] = {-9'd99,-10'd299};
ram[5559] = {-9'd96,-10'd296};
ram[5560] = {-9'd92,-10'd293};
ram[5561] = {-9'd89,-10'd290};
ram[5562] = {-9'd86,-10'd286};
ram[5563] = {-9'd83,-10'd283};
ram[5564] = {-9'd80,-10'd280};
ram[5565] = {-9'd77,-10'd277};
ram[5566] = {-9'd74,-10'd274};
ram[5567] = {-9'd70,-10'd271};
ram[5568] = {-9'd67,-10'd268};
ram[5569] = {-9'd64,-10'd264};
ram[5570] = {-9'd61,-10'd261};
ram[5571] = {-9'd58,-10'd258};
ram[5572] = {-9'd55,-10'd255};
ram[5573] = {-9'd52,-10'd252};
ram[5574] = {-9'd48,-10'd249};
ram[5575] = {-9'd45,-10'd246};
ram[5576] = {-9'd42,-10'd242};
ram[5577] = {-9'd39,-10'd239};
ram[5578] = {-9'd36,-10'd236};
ram[5579] = {-9'd33,-10'd233};
ram[5580] = {-9'd30,-10'd230};
ram[5581] = {-9'd26,-10'd227};
ram[5582] = {-9'd23,-10'd224};
ram[5583] = {-9'd20,-10'd220};
ram[5584] = {-9'd17,-10'd217};
ram[5585] = {-9'd14,-10'd214};
ram[5586] = {-9'd11,-10'd211};
ram[5587] = {-9'd8,-10'd208};
ram[5588] = {-9'd4,-10'd205};
ram[5589] = {-9'd1,-10'd202};
ram[5590] = {9'd2,-10'd198};
ram[5591] = {9'd5,-10'd195};
ram[5592] = {9'd8,-10'd192};
ram[5593] = {9'd11,-10'd189};
ram[5594] = {9'd14,-10'd186};
ram[5595] = {9'd18,-10'd183};
ram[5596] = {9'd21,-10'd180};
ram[5597] = {9'd24,-10'd176};
ram[5598] = {9'd27,-10'd173};
ram[5599] = {9'd30,-10'd170};
ram[5600] = {9'd33,-10'd167};
ram[5601] = {9'd36,-10'd164};
ram[5602] = {9'd40,-10'd161};
ram[5603] = {9'd43,-10'd158};
ram[5604] = {9'd46,-10'd154};
ram[5605] = {9'd49,-10'd151};
ram[5606] = {9'd52,-10'd148};
ram[5607] = {9'd55,-10'd145};
ram[5608] = {9'd58,-10'd142};
ram[5609] = {9'd62,-10'd139};
ram[5610] = {9'd65,-10'd136};
ram[5611] = {9'd68,-10'd132};
ram[5612] = {9'd71,-10'd129};
ram[5613] = {9'd74,-10'd126};
ram[5614] = {9'd77,-10'd123};
ram[5615] = {9'd80,-10'd120};
ram[5616] = {9'd84,-10'd117};
ram[5617] = {9'd87,-10'd114};
ram[5618] = {9'd90,-10'd110};
ram[5619] = {9'd93,-10'd107};
ram[5620] = {9'd96,-10'd104};
ram[5621] = {9'd99,-10'd101};
ram[5622] = {-9'd98,-10'd98};
ram[5623] = {-9'd95,-10'd95};
ram[5624] = {-9'd92,-10'd92};
ram[5625] = {-9'd88,-10'd88};
ram[5626] = {-9'd85,-10'd85};
ram[5627] = {-9'd82,-10'd82};
ram[5628] = {-9'd79,-10'd79};
ram[5629] = {-9'd76,-10'd76};
ram[5630] = {-9'd73,-10'd73};
ram[5631] = {-9'd70,-10'd70};
ram[5632] = {-9'd70,-10'd70};
ram[5633] = {-9'd66,-10'd66};
ram[5634] = {-9'd63,-10'd63};
ram[5635] = {-9'd60,-10'd60};
ram[5636] = {-9'd57,-10'd57};
ram[5637] = {-9'd54,-10'd54};
ram[5638] = {-9'd51,-10'd51};
ram[5639] = {-9'd48,-10'd48};
ram[5640] = {-9'd44,-10'd44};
ram[5641] = {-9'd41,-10'd41};
ram[5642] = {-9'd38,-10'd38};
ram[5643] = {-9'd35,-10'd35};
ram[5644] = {-9'd32,-10'd32};
ram[5645] = {-9'd29,-10'd29};
ram[5646] = {-9'd26,-10'd26};
ram[5647] = {-9'd22,-10'd22};
ram[5648] = {-9'd19,-10'd19};
ram[5649] = {-9'd16,-10'd16};
ram[5650] = {-9'd13,-10'd13};
ram[5651] = {-9'd10,-10'd10};
ram[5652] = {-9'd7,-10'd7};
ram[5653] = {-9'd4,-10'd4};
ram[5654] = {9'd0,10'd0};
ram[5655] = {9'd3,10'd3};
ram[5656] = {9'd6,10'd6};
ram[5657] = {9'd9,10'd9};
ram[5658] = {9'd12,10'd12};
ram[5659] = {9'd15,10'd15};
ram[5660] = {9'd18,10'd18};
ram[5661] = {9'd21,10'd21};
ram[5662] = {9'd25,10'd25};
ram[5663] = {9'd28,10'd28};
ram[5664] = {9'd31,10'd31};
ram[5665] = {9'd34,10'd34};
ram[5666] = {9'd37,10'd37};
ram[5667] = {9'd40,10'd40};
ram[5668] = {9'd43,10'd43};
ram[5669] = {9'd47,10'd47};
ram[5670] = {9'd50,10'd50};
ram[5671] = {9'd53,10'd53};
ram[5672] = {9'd56,10'd56};
ram[5673] = {9'd59,10'd59};
ram[5674] = {9'd62,10'd62};
ram[5675] = {9'd65,10'd65};
ram[5676] = {9'd69,10'd69};
ram[5677] = {9'd72,10'd72};
ram[5678] = {9'd75,10'd75};
ram[5679] = {9'd78,10'd78};
ram[5680] = {9'd81,10'd81};
ram[5681] = {9'd84,10'd84};
ram[5682] = {9'd87,10'd87};
ram[5683] = {9'd91,10'd91};
ram[5684] = {9'd94,10'd94};
ram[5685] = {9'd97,10'd97};
ram[5686] = {-9'd100,10'd100};
ram[5687] = {-9'd97,10'd103};
ram[5688] = {-9'd94,10'd106};
ram[5689] = {-9'd91,10'd109};
ram[5690] = {-9'd88,10'd113};
ram[5691] = {-9'd85,10'd116};
ram[5692] = {-9'd81,10'd119};
ram[5693] = {-9'd78,10'd122};
ram[5694] = {-9'd75,10'd125};
ram[5695] = {-9'd72,10'd128};
ram[5696] = {-9'd69,10'd131};
ram[5697] = {-9'd66,10'd135};
ram[5698] = {-9'd63,10'd138};
ram[5699] = {-9'd59,10'd141};
ram[5700] = {-9'd56,10'd144};
ram[5701] = {-9'd53,10'd147};
ram[5702] = {-9'd50,10'd150};
ram[5703] = {-9'd47,10'd153};
ram[5704] = {-9'd44,10'd157};
ram[5705] = {-9'd41,10'd160};
ram[5706] = {-9'd37,10'd163};
ram[5707] = {-9'd34,10'd166};
ram[5708] = {-9'd31,10'd169};
ram[5709] = {-9'd28,10'd172};
ram[5710] = {-9'd25,10'd175};
ram[5711] = {-9'd22,10'd179};
ram[5712] = {-9'd19,10'd182};
ram[5713] = {-9'd15,10'd185};
ram[5714] = {-9'd12,10'd188};
ram[5715] = {-9'd9,10'd191};
ram[5716] = {-9'd6,10'd194};
ram[5717] = {-9'd3,10'd197};
ram[5718] = {9'd0,10'd201};
ram[5719] = {9'd3,10'd204};
ram[5720] = {9'd7,10'd207};
ram[5721] = {9'd10,10'd210};
ram[5722] = {9'd13,10'd213};
ram[5723] = {9'd16,10'd216};
ram[5724] = {9'd19,10'd219};
ram[5725] = {9'd22,10'd223};
ram[5726] = {9'd25,10'd226};
ram[5727] = {9'd29,10'd229};
ram[5728] = {9'd32,10'd232};
ram[5729] = {9'd35,10'd235};
ram[5730] = {9'd38,10'd238};
ram[5731] = {9'd41,10'd241};
ram[5732] = {9'd44,10'd245};
ram[5733] = {9'd47,10'd248};
ram[5734] = {9'd51,10'd251};
ram[5735] = {9'd54,10'd254};
ram[5736] = {9'd57,10'd257};
ram[5737] = {9'd60,10'd260};
ram[5738] = {9'd63,10'd263};
ram[5739] = {9'd66,10'd267};
ram[5740] = {9'd69,10'd270};
ram[5741] = {9'd73,10'd273};
ram[5742] = {9'd76,10'd276};
ram[5743] = {9'd79,10'd279};
ram[5744] = {9'd82,10'd282};
ram[5745] = {9'd85,10'd285};
ram[5746] = {9'd88,10'd289};
ram[5747] = {9'd91,10'd292};
ram[5748] = {9'd95,10'd295};
ram[5749] = {9'd98,10'd298};
ram[5750] = {-9'd99,10'd301};
ram[5751] = {-9'd96,10'd304};
ram[5752] = {-9'd93,10'd307};
ram[5753] = {-9'd90,10'd311};
ram[5754] = {-9'd87,10'd314};
ram[5755] = {-9'd84,10'd317};
ram[5756] = {-9'd81,10'd320};
ram[5757] = {-9'd77,10'd323};
ram[5758] = {-9'd74,10'd326};
ram[5759] = {-9'd71,10'd329};
ram[5760] = {-9'd71,10'd329};
ram[5761] = {-9'd68,10'd333};
ram[5762] = {-9'd65,10'd336};
ram[5763] = {-9'd62,10'd339};
ram[5764] = {-9'd59,10'd342};
ram[5765] = {-9'd55,10'd345};
ram[5766] = {-9'd52,10'd348};
ram[5767] = {-9'd49,10'd351};
ram[5768] = {-9'd46,10'd354};
ram[5769] = {-9'd43,10'd358};
ram[5770] = {-9'd40,10'd361};
ram[5771] = {-9'd37,10'd364};
ram[5772] = {-9'd33,10'd367};
ram[5773] = {-9'd30,10'd370};
ram[5774] = {-9'd27,10'd373};
ram[5775] = {-9'd24,10'd376};
ram[5776] = {-9'd21,10'd380};
ram[5777] = {-9'd18,10'd383};
ram[5778] = {-9'd15,10'd386};
ram[5779] = {-9'd11,10'd389};
ram[5780] = {-9'd8,10'd392};
ram[5781] = {-9'd5,10'd395};
ram[5782] = {-9'd2,10'd398};
ram[5783] = {9'd1,-10'd399};
ram[5784] = {9'd4,-10'd396};
ram[5785] = {9'd7,-10'd393};
ram[5786] = {9'd10,-10'd390};
ram[5787] = {9'd14,-10'd387};
ram[5788] = {9'd17,-10'd384};
ram[5789] = {9'd20,-10'd381};
ram[5790] = {9'd23,-10'd377};
ram[5791] = {9'd26,-10'd374};
ram[5792] = {9'd29,-10'd371};
ram[5793] = {9'd32,-10'd368};
ram[5794] = {9'd36,-10'd365};
ram[5795] = {9'd39,-10'd362};
ram[5796] = {9'd42,-10'd359};
ram[5797] = {9'd45,-10'd355};
ram[5798] = {9'd48,-10'd352};
ram[5799] = {9'd51,-10'd349};
ram[5800] = {9'd54,-10'd346};
ram[5801] = {9'd58,-10'd343};
ram[5802] = {9'd61,-10'd340};
ram[5803] = {9'd64,-10'd337};
ram[5804] = {9'd67,-10'd334};
ram[5805] = {9'd70,-10'd330};
ram[5806] = {9'd73,-10'd327};
ram[5807] = {9'd76,-10'd324};
ram[5808] = {9'd80,-10'd321};
ram[5809] = {9'd83,-10'd318};
ram[5810] = {9'd86,-10'd315};
ram[5811] = {9'd89,-10'd312};
ram[5812] = {9'd92,-10'd308};
ram[5813] = {9'd95,-10'd305};
ram[5814] = {9'd98,-10'd302};
ram[5815] = {-9'd99,-10'd299};
ram[5816] = {-9'd96,-10'd296};
ram[5817] = {-9'd92,-10'd293};
ram[5818] = {-9'd89,-10'd290};
ram[5819] = {-9'd86,-10'd286};
ram[5820] = {-9'd83,-10'd283};
ram[5821] = {-9'd80,-10'd280};
ram[5822] = {-9'd77,-10'd277};
ram[5823] = {-9'd74,-10'd274};
ram[5824] = {-9'd70,-10'd271};
ram[5825] = {-9'd67,-10'd268};
ram[5826] = {-9'd64,-10'd264};
ram[5827] = {-9'd61,-10'd261};
ram[5828] = {-9'd58,-10'd258};
ram[5829] = {-9'd55,-10'd255};
ram[5830] = {-9'd52,-10'd252};
ram[5831] = {-9'd48,-10'd249};
ram[5832] = {-9'd45,-10'd246};
ram[5833] = {-9'd42,-10'd242};
ram[5834] = {-9'd39,-10'd239};
ram[5835] = {-9'd36,-10'd236};
ram[5836] = {-9'd33,-10'd233};
ram[5837] = {-9'd30,-10'd230};
ram[5838] = {-9'd26,-10'd227};
ram[5839] = {-9'd23,-10'd224};
ram[5840] = {-9'd20,-10'd220};
ram[5841] = {-9'd17,-10'd217};
ram[5842] = {-9'd14,-10'd214};
ram[5843] = {-9'd11,-10'd211};
ram[5844] = {-9'd8,-10'd208};
ram[5845] = {-9'd4,-10'd205};
ram[5846] = {-9'd1,-10'd202};
ram[5847] = {9'd2,-10'd198};
ram[5848] = {9'd5,-10'd195};
ram[5849] = {9'd8,-10'd192};
ram[5850] = {9'd11,-10'd189};
ram[5851] = {9'd14,-10'd186};
ram[5852] = {9'd18,-10'd183};
ram[5853] = {9'd21,-10'd180};
ram[5854] = {9'd24,-10'd176};
ram[5855] = {9'd27,-10'd173};
ram[5856] = {9'd30,-10'd170};
ram[5857] = {9'd33,-10'd167};
ram[5858] = {9'd36,-10'd164};
ram[5859] = {9'd40,-10'd161};
ram[5860] = {9'd43,-10'd158};
ram[5861] = {9'd46,-10'd154};
ram[5862] = {9'd49,-10'd151};
ram[5863] = {9'd52,-10'd148};
ram[5864] = {9'd55,-10'd145};
ram[5865] = {9'd58,-10'd142};
ram[5866] = {9'd62,-10'd139};
ram[5867] = {9'd65,-10'd136};
ram[5868] = {9'd68,-10'd132};
ram[5869] = {9'd71,-10'd129};
ram[5870] = {9'd74,-10'd126};
ram[5871] = {9'd77,-10'd123};
ram[5872] = {9'd80,-10'd120};
ram[5873] = {9'd84,-10'd117};
ram[5874] = {9'd87,-10'd114};
ram[5875] = {9'd90,-10'd110};
ram[5876] = {9'd93,-10'd107};
ram[5877] = {9'd96,-10'd104};
ram[5878] = {9'd99,-10'd101};
ram[5879] = {-9'd98,-10'd98};
ram[5880] = {-9'd95,-10'd95};
ram[5881] = {-9'd92,-10'd92};
ram[5882] = {-9'd88,-10'd88};
ram[5883] = {-9'd85,-10'd85};
ram[5884] = {-9'd82,-10'd82};
ram[5885] = {-9'd79,-10'd79};
ram[5886] = {-9'd76,-10'd76};
ram[5887] = {-9'd73,-10'd73};
ram[5888] = {-9'd73,-10'd73};
ram[5889] = {-9'd70,-10'd70};
ram[5890] = {-9'd66,-10'd66};
ram[5891] = {-9'd63,-10'd63};
ram[5892] = {-9'd60,-10'd60};
ram[5893] = {-9'd57,-10'd57};
ram[5894] = {-9'd54,-10'd54};
ram[5895] = {-9'd51,-10'd51};
ram[5896] = {-9'd48,-10'd48};
ram[5897] = {-9'd44,-10'd44};
ram[5898] = {-9'd41,-10'd41};
ram[5899] = {-9'd38,-10'd38};
ram[5900] = {-9'd35,-10'd35};
ram[5901] = {-9'd32,-10'd32};
ram[5902] = {-9'd29,-10'd29};
ram[5903] = {-9'd26,-10'd26};
ram[5904] = {-9'd22,-10'd22};
ram[5905] = {-9'd19,-10'd19};
ram[5906] = {-9'd16,-10'd16};
ram[5907] = {-9'd13,-10'd13};
ram[5908] = {-9'd10,-10'd10};
ram[5909] = {-9'd7,-10'd7};
ram[5910] = {-9'd4,-10'd4};
ram[5911] = {9'd0,10'd0};
ram[5912] = {9'd3,10'd3};
ram[5913] = {9'd6,10'd6};
ram[5914] = {9'd9,10'd9};
ram[5915] = {9'd12,10'd12};
ram[5916] = {9'd15,10'd15};
ram[5917] = {9'd18,10'd18};
ram[5918] = {9'd21,10'd21};
ram[5919] = {9'd25,10'd25};
ram[5920] = {9'd28,10'd28};
ram[5921] = {9'd31,10'd31};
ram[5922] = {9'd34,10'd34};
ram[5923] = {9'd37,10'd37};
ram[5924] = {9'd40,10'd40};
ram[5925] = {9'd43,10'd43};
ram[5926] = {9'd47,10'd47};
ram[5927] = {9'd50,10'd50};
ram[5928] = {9'd53,10'd53};
ram[5929] = {9'd56,10'd56};
ram[5930] = {9'd59,10'd59};
ram[5931] = {9'd62,10'd62};
ram[5932] = {9'd65,10'd65};
ram[5933] = {9'd69,10'd69};
ram[5934] = {9'd72,10'd72};
ram[5935] = {9'd75,10'd75};
ram[5936] = {9'd78,10'd78};
ram[5937] = {9'd81,10'd81};
ram[5938] = {9'd84,10'd84};
ram[5939] = {9'd87,10'd87};
ram[5940] = {9'd91,10'd91};
ram[5941] = {9'd94,10'd94};
ram[5942] = {9'd97,10'd97};
ram[5943] = {-9'd100,10'd100};
ram[5944] = {-9'd97,10'd103};
ram[5945] = {-9'd94,10'd106};
ram[5946] = {-9'd91,10'd109};
ram[5947] = {-9'd88,10'd113};
ram[5948] = {-9'd85,10'd116};
ram[5949] = {-9'd81,10'd119};
ram[5950] = {-9'd78,10'd122};
ram[5951] = {-9'd75,10'd125};
ram[5952] = {-9'd72,10'd128};
ram[5953] = {-9'd69,10'd131};
ram[5954] = {-9'd66,10'd135};
ram[5955] = {-9'd63,10'd138};
ram[5956] = {-9'd59,10'd141};
ram[5957] = {-9'd56,10'd144};
ram[5958] = {-9'd53,10'd147};
ram[5959] = {-9'd50,10'd150};
ram[5960] = {-9'd47,10'd153};
ram[5961] = {-9'd44,10'd157};
ram[5962] = {-9'd41,10'd160};
ram[5963] = {-9'd37,10'd163};
ram[5964] = {-9'd34,10'd166};
ram[5965] = {-9'd31,10'd169};
ram[5966] = {-9'd28,10'd172};
ram[5967] = {-9'd25,10'd175};
ram[5968] = {-9'd22,10'd179};
ram[5969] = {-9'd19,10'd182};
ram[5970] = {-9'd15,10'd185};
ram[5971] = {-9'd12,10'd188};
ram[5972] = {-9'd9,10'd191};
ram[5973] = {-9'd6,10'd194};
ram[5974] = {-9'd3,10'd197};
ram[5975] = {9'd0,10'd201};
ram[5976] = {9'd3,10'd204};
ram[5977] = {9'd7,10'd207};
ram[5978] = {9'd10,10'd210};
ram[5979] = {9'd13,10'd213};
ram[5980] = {9'd16,10'd216};
ram[5981] = {9'd19,10'd219};
ram[5982] = {9'd22,10'd223};
ram[5983] = {9'd25,10'd226};
ram[5984] = {9'd29,10'd229};
ram[5985] = {9'd32,10'd232};
ram[5986] = {9'd35,10'd235};
ram[5987] = {9'd38,10'd238};
ram[5988] = {9'd41,10'd241};
ram[5989] = {9'd44,10'd245};
ram[5990] = {9'd47,10'd248};
ram[5991] = {9'd51,10'd251};
ram[5992] = {9'd54,10'd254};
ram[5993] = {9'd57,10'd257};
ram[5994] = {9'd60,10'd260};
ram[5995] = {9'd63,10'd263};
ram[5996] = {9'd66,10'd267};
ram[5997] = {9'd69,10'd270};
ram[5998] = {9'd73,10'd273};
ram[5999] = {9'd76,10'd276};
ram[6000] = {9'd79,10'd279};
ram[6001] = {9'd82,10'd282};
ram[6002] = {9'd85,10'd285};
ram[6003] = {9'd88,10'd289};
ram[6004] = {9'd91,10'd292};
ram[6005] = {9'd95,10'd295};
ram[6006] = {9'd98,10'd298};
ram[6007] = {-9'd99,10'd301};
ram[6008] = {-9'd96,10'd304};
ram[6009] = {-9'd93,10'd307};
ram[6010] = {-9'd90,10'd311};
ram[6011] = {-9'd87,10'd314};
ram[6012] = {-9'd84,10'd317};
ram[6013] = {-9'd81,10'd320};
ram[6014] = {-9'd77,10'd323};
ram[6015] = {-9'd74,10'd326};
ram[6016] = {-9'd74,10'd326};
ram[6017] = {-9'd71,10'd329};
ram[6018] = {-9'd68,10'd333};
ram[6019] = {-9'd65,10'd336};
ram[6020] = {-9'd62,10'd339};
ram[6021] = {-9'd59,10'd342};
ram[6022] = {-9'd55,10'd345};
ram[6023] = {-9'd52,10'd348};
ram[6024] = {-9'd49,10'd351};
ram[6025] = {-9'd46,10'd354};
ram[6026] = {-9'd43,10'd358};
ram[6027] = {-9'd40,10'd361};
ram[6028] = {-9'd37,10'd364};
ram[6029] = {-9'd33,10'd367};
ram[6030] = {-9'd30,10'd370};
ram[6031] = {-9'd27,10'd373};
ram[6032] = {-9'd24,10'd376};
ram[6033] = {-9'd21,10'd380};
ram[6034] = {-9'd18,10'd383};
ram[6035] = {-9'd15,10'd386};
ram[6036] = {-9'd11,10'd389};
ram[6037] = {-9'd8,10'd392};
ram[6038] = {-9'd5,10'd395};
ram[6039] = {-9'd2,10'd398};
ram[6040] = {9'd1,-10'd399};
ram[6041] = {9'd4,-10'd396};
ram[6042] = {9'd7,-10'd393};
ram[6043] = {9'd10,-10'd390};
ram[6044] = {9'd14,-10'd387};
ram[6045] = {9'd17,-10'd384};
ram[6046] = {9'd20,-10'd381};
ram[6047] = {9'd23,-10'd377};
ram[6048] = {9'd26,-10'd374};
ram[6049] = {9'd29,-10'd371};
ram[6050] = {9'd32,-10'd368};
ram[6051] = {9'd36,-10'd365};
ram[6052] = {9'd39,-10'd362};
ram[6053] = {9'd42,-10'd359};
ram[6054] = {9'd45,-10'd355};
ram[6055] = {9'd48,-10'd352};
ram[6056] = {9'd51,-10'd349};
ram[6057] = {9'd54,-10'd346};
ram[6058] = {9'd58,-10'd343};
ram[6059] = {9'd61,-10'd340};
ram[6060] = {9'd64,-10'd337};
ram[6061] = {9'd67,-10'd334};
ram[6062] = {9'd70,-10'd330};
ram[6063] = {9'd73,-10'd327};
ram[6064] = {9'd76,-10'd324};
ram[6065] = {9'd80,-10'd321};
ram[6066] = {9'd83,-10'd318};
ram[6067] = {9'd86,-10'd315};
ram[6068] = {9'd89,-10'd312};
ram[6069] = {9'd92,-10'd308};
ram[6070] = {9'd95,-10'd305};
ram[6071] = {9'd98,-10'd302};
ram[6072] = {-9'd99,-10'd299};
ram[6073] = {-9'd96,-10'd296};
ram[6074] = {-9'd92,-10'd293};
ram[6075] = {-9'd89,-10'd290};
ram[6076] = {-9'd86,-10'd286};
ram[6077] = {-9'd83,-10'd283};
ram[6078] = {-9'd80,-10'd280};
ram[6079] = {-9'd77,-10'd277};
ram[6080] = {-9'd74,-10'd274};
ram[6081] = {-9'd70,-10'd271};
ram[6082] = {-9'd67,-10'd268};
ram[6083] = {-9'd64,-10'd264};
ram[6084] = {-9'd61,-10'd261};
ram[6085] = {-9'd58,-10'd258};
ram[6086] = {-9'd55,-10'd255};
ram[6087] = {-9'd52,-10'd252};
ram[6088] = {-9'd48,-10'd249};
ram[6089] = {-9'd45,-10'd246};
ram[6090] = {-9'd42,-10'd242};
ram[6091] = {-9'd39,-10'd239};
ram[6092] = {-9'd36,-10'd236};
ram[6093] = {-9'd33,-10'd233};
ram[6094] = {-9'd30,-10'd230};
ram[6095] = {-9'd26,-10'd227};
ram[6096] = {-9'd23,-10'd224};
ram[6097] = {-9'd20,-10'd220};
ram[6098] = {-9'd17,-10'd217};
ram[6099] = {-9'd14,-10'd214};
ram[6100] = {-9'd11,-10'd211};
ram[6101] = {-9'd8,-10'd208};
ram[6102] = {-9'd4,-10'd205};
ram[6103] = {-9'd1,-10'd202};
ram[6104] = {9'd2,-10'd198};
ram[6105] = {9'd5,-10'd195};
ram[6106] = {9'd8,-10'd192};
ram[6107] = {9'd11,-10'd189};
ram[6108] = {9'd14,-10'd186};
ram[6109] = {9'd18,-10'd183};
ram[6110] = {9'd21,-10'd180};
ram[6111] = {9'd24,-10'd176};
ram[6112] = {9'd27,-10'd173};
ram[6113] = {9'd30,-10'd170};
ram[6114] = {9'd33,-10'd167};
ram[6115] = {9'd36,-10'd164};
ram[6116] = {9'd40,-10'd161};
ram[6117] = {9'd43,-10'd158};
ram[6118] = {9'd46,-10'd154};
ram[6119] = {9'd49,-10'd151};
ram[6120] = {9'd52,-10'd148};
ram[6121] = {9'd55,-10'd145};
ram[6122] = {9'd58,-10'd142};
ram[6123] = {9'd62,-10'd139};
ram[6124] = {9'd65,-10'd136};
ram[6125] = {9'd68,-10'd132};
ram[6126] = {9'd71,-10'd129};
ram[6127] = {9'd74,-10'd126};
ram[6128] = {9'd77,-10'd123};
ram[6129] = {9'd80,-10'd120};
ram[6130] = {9'd84,-10'd117};
ram[6131] = {9'd87,-10'd114};
ram[6132] = {9'd90,-10'd110};
ram[6133] = {9'd93,-10'd107};
ram[6134] = {9'd96,-10'd104};
ram[6135] = {9'd99,-10'd101};
ram[6136] = {-9'd98,-10'd98};
ram[6137] = {-9'd95,-10'd95};
ram[6138] = {-9'd92,-10'd92};
ram[6139] = {-9'd88,-10'd88};
ram[6140] = {-9'd85,-10'd85};
ram[6141] = {-9'd82,-10'd82};
ram[6142] = {-9'd79,-10'd79};
ram[6143] = {-9'd76,-10'd76};
ram[6144] = {-9'd76,-10'd76};
ram[6145] = {-9'd73,-10'd73};
ram[6146] = {-9'd70,-10'd70};
ram[6147] = {-9'd66,-10'd66};
ram[6148] = {-9'd63,-10'd63};
ram[6149] = {-9'd60,-10'd60};
ram[6150] = {-9'd57,-10'd57};
ram[6151] = {-9'd54,-10'd54};
ram[6152] = {-9'd51,-10'd51};
ram[6153] = {-9'd48,-10'd48};
ram[6154] = {-9'd44,-10'd44};
ram[6155] = {-9'd41,-10'd41};
ram[6156] = {-9'd38,-10'd38};
ram[6157] = {-9'd35,-10'd35};
ram[6158] = {-9'd32,-10'd32};
ram[6159] = {-9'd29,-10'd29};
ram[6160] = {-9'd26,-10'd26};
ram[6161] = {-9'd22,-10'd22};
ram[6162] = {-9'd19,-10'd19};
ram[6163] = {-9'd16,-10'd16};
ram[6164] = {-9'd13,-10'd13};
ram[6165] = {-9'd10,-10'd10};
ram[6166] = {-9'd7,-10'd7};
ram[6167] = {-9'd4,-10'd4};
ram[6168] = {9'd0,10'd0};
ram[6169] = {9'd3,10'd3};
ram[6170] = {9'd6,10'd6};
ram[6171] = {9'd9,10'd9};
ram[6172] = {9'd12,10'd12};
ram[6173] = {9'd15,10'd15};
ram[6174] = {9'd18,10'd18};
ram[6175] = {9'd21,10'd21};
ram[6176] = {9'd25,10'd25};
ram[6177] = {9'd28,10'd28};
ram[6178] = {9'd31,10'd31};
ram[6179] = {9'd34,10'd34};
ram[6180] = {9'd37,10'd37};
ram[6181] = {9'd40,10'd40};
ram[6182] = {9'd43,10'd43};
ram[6183] = {9'd47,10'd47};
ram[6184] = {9'd50,10'd50};
ram[6185] = {9'd53,10'd53};
ram[6186] = {9'd56,10'd56};
ram[6187] = {9'd59,10'd59};
ram[6188] = {9'd62,10'd62};
ram[6189] = {9'd65,10'd65};
ram[6190] = {9'd69,10'd69};
ram[6191] = {9'd72,10'd72};
ram[6192] = {9'd75,10'd75};
ram[6193] = {9'd78,10'd78};
ram[6194] = {9'd81,10'd81};
ram[6195] = {9'd84,10'd84};
ram[6196] = {9'd87,10'd87};
ram[6197] = {9'd91,10'd91};
ram[6198] = {9'd94,10'd94};
ram[6199] = {9'd97,10'd97};
ram[6200] = {-9'd100,10'd100};
ram[6201] = {-9'd97,10'd103};
ram[6202] = {-9'd94,10'd106};
ram[6203] = {-9'd91,10'd109};
ram[6204] = {-9'd88,10'd113};
ram[6205] = {-9'd85,10'd116};
ram[6206] = {-9'd81,10'd119};
ram[6207] = {-9'd78,10'd122};
ram[6208] = {-9'd75,10'd125};
ram[6209] = {-9'd72,10'd128};
ram[6210] = {-9'd69,10'd131};
ram[6211] = {-9'd66,10'd135};
ram[6212] = {-9'd63,10'd138};
ram[6213] = {-9'd59,10'd141};
ram[6214] = {-9'd56,10'd144};
ram[6215] = {-9'd53,10'd147};
ram[6216] = {-9'd50,10'd150};
ram[6217] = {-9'd47,10'd153};
ram[6218] = {-9'd44,10'd157};
ram[6219] = {-9'd41,10'd160};
ram[6220] = {-9'd37,10'd163};
ram[6221] = {-9'd34,10'd166};
ram[6222] = {-9'd31,10'd169};
ram[6223] = {-9'd28,10'd172};
ram[6224] = {-9'd25,10'd175};
ram[6225] = {-9'd22,10'd179};
ram[6226] = {-9'd19,10'd182};
ram[6227] = {-9'd15,10'd185};
ram[6228] = {-9'd12,10'd188};
ram[6229] = {-9'd9,10'd191};
ram[6230] = {-9'd6,10'd194};
ram[6231] = {-9'd3,10'd197};
ram[6232] = {9'd0,10'd201};
ram[6233] = {9'd3,10'd204};
ram[6234] = {9'd7,10'd207};
ram[6235] = {9'd10,10'd210};
ram[6236] = {9'd13,10'd213};
ram[6237] = {9'd16,10'd216};
ram[6238] = {9'd19,10'd219};
ram[6239] = {9'd22,10'd223};
ram[6240] = {9'd25,10'd226};
ram[6241] = {9'd29,10'd229};
ram[6242] = {9'd32,10'd232};
ram[6243] = {9'd35,10'd235};
ram[6244] = {9'd38,10'd238};
ram[6245] = {9'd41,10'd241};
ram[6246] = {9'd44,10'd245};
ram[6247] = {9'd47,10'd248};
ram[6248] = {9'd51,10'd251};
ram[6249] = {9'd54,10'd254};
ram[6250] = {9'd57,10'd257};
ram[6251] = {9'd60,10'd260};
ram[6252] = {9'd63,10'd263};
ram[6253] = {9'd66,10'd267};
ram[6254] = {9'd69,10'd270};
ram[6255] = {9'd73,10'd273};
ram[6256] = {9'd76,10'd276};
ram[6257] = {9'd79,10'd279};
ram[6258] = {9'd82,10'd282};
ram[6259] = {9'd85,10'd285};
ram[6260] = {9'd88,10'd289};
ram[6261] = {9'd91,10'd292};
ram[6262] = {9'd95,10'd295};
ram[6263] = {9'd98,10'd298};
ram[6264] = {-9'd99,10'd301};
ram[6265] = {-9'd96,10'd304};
ram[6266] = {-9'd93,10'd307};
ram[6267] = {-9'd90,10'd311};
ram[6268] = {-9'd87,10'd314};
ram[6269] = {-9'd84,10'd317};
ram[6270] = {-9'd81,10'd320};
ram[6271] = {-9'd77,10'd323};
ram[6272] = {-9'd77,10'd323};
ram[6273] = {-9'd74,10'd326};
ram[6274] = {-9'd71,10'd329};
ram[6275] = {-9'd68,10'd333};
ram[6276] = {-9'd65,10'd336};
ram[6277] = {-9'd62,10'd339};
ram[6278] = {-9'd59,10'd342};
ram[6279] = {-9'd55,10'd345};
ram[6280] = {-9'd52,10'd348};
ram[6281] = {-9'd49,10'd351};
ram[6282] = {-9'd46,10'd354};
ram[6283] = {-9'd43,10'd358};
ram[6284] = {-9'd40,10'd361};
ram[6285] = {-9'd37,10'd364};
ram[6286] = {-9'd33,10'd367};
ram[6287] = {-9'd30,10'd370};
ram[6288] = {-9'd27,10'd373};
ram[6289] = {-9'd24,10'd376};
ram[6290] = {-9'd21,10'd380};
ram[6291] = {-9'd18,10'd383};
ram[6292] = {-9'd15,10'd386};
ram[6293] = {-9'd11,10'd389};
ram[6294] = {-9'd8,10'd392};
ram[6295] = {-9'd5,10'd395};
ram[6296] = {-9'd2,10'd398};
ram[6297] = {9'd1,-10'd399};
ram[6298] = {9'd4,-10'd396};
ram[6299] = {9'd7,-10'd393};
ram[6300] = {9'd10,-10'd390};
ram[6301] = {9'd14,-10'd387};
ram[6302] = {9'd17,-10'd384};
ram[6303] = {9'd20,-10'd381};
ram[6304] = {9'd23,-10'd377};
ram[6305] = {9'd26,-10'd374};
ram[6306] = {9'd29,-10'd371};
ram[6307] = {9'd32,-10'd368};
ram[6308] = {9'd36,-10'd365};
ram[6309] = {9'd39,-10'd362};
ram[6310] = {9'd42,-10'd359};
ram[6311] = {9'd45,-10'd355};
ram[6312] = {9'd48,-10'd352};
ram[6313] = {9'd51,-10'd349};
ram[6314] = {9'd54,-10'd346};
ram[6315] = {9'd58,-10'd343};
ram[6316] = {9'd61,-10'd340};
ram[6317] = {9'd64,-10'd337};
ram[6318] = {9'd67,-10'd334};
ram[6319] = {9'd70,-10'd330};
ram[6320] = {9'd73,-10'd327};
ram[6321] = {9'd76,-10'd324};
ram[6322] = {9'd80,-10'd321};
ram[6323] = {9'd83,-10'd318};
ram[6324] = {9'd86,-10'd315};
ram[6325] = {9'd89,-10'd312};
ram[6326] = {9'd92,-10'd308};
ram[6327] = {9'd95,-10'd305};
ram[6328] = {9'd98,-10'd302};
ram[6329] = {-9'd99,-10'd299};
ram[6330] = {-9'd96,-10'd296};
ram[6331] = {-9'd92,-10'd293};
ram[6332] = {-9'd89,-10'd290};
ram[6333] = {-9'd86,-10'd286};
ram[6334] = {-9'd83,-10'd283};
ram[6335] = {-9'd80,-10'd280};
ram[6336] = {-9'd77,-10'd277};
ram[6337] = {-9'd74,-10'd274};
ram[6338] = {-9'd70,-10'd271};
ram[6339] = {-9'd67,-10'd268};
ram[6340] = {-9'd64,-10'd264};
ram[6341] = {-9'd61,-10'd261};
ram[6342] = {-9'd58,-10'd258};
ram[6343] = {-9'd55,-10'd255};
ram[6344] = {-9'd52,-10'd252};
ram[6345] = {-9'd48,-10'd249};
ram[6346] = {-9'd45,-10'd246};
ram[6347] = {-9'd42,-10'd242};
ram[6348] = {-9'd39,-10'd239};
ram[6349] = {-9'd36,-10'd236};
ram[6350] = {-9'd33,-10'd233};
ram[6351] = {-9'd30,-10'd230};
ram[6352] = {-9'd26,-10'd227};
ram[6353] = {-9'd23,-10'd224};
ram[6354] = {-9'd20,-10'd220};
ram[6355] = {-9'd17,-10'd217};
ram[6356] = {-9'd14,-10'd214};
ram[6357] = {-9'd11,-10'd211};
ram[6358] = {-9'd8,-10'd208};
ram[6359] = {-9'd4,-10'd205};
ram[6360] = {-9'd1,-10'd202};
ram[6361] = {9'd2,-10'd198};
ram[6362] = {9'd5,-10'd195};
ram[6363] = {9'd8,-10'd192};
ram[6364] = {9'd11,-10'd189};
ram[6365] = {9'd14,-10'd186};
ram[6366] = {9'd18,-10'd183};
ram[6367] = {9'd21,-10'd180};
ram[6368] = {9'd24,-10'd176};
ram[6369] = {9'd27,-10'd173};
ram[6370] = {9'd30,-10'd170};
ram[6371] = {9'd33,-10'd167};
ram[6372] = {9'd36,-10'd164};
ram[6373] = {9'd40,-10'd161};
ram[6374] = {9'd43,-10'd158};
ram[6375] = {9'd46,-10'd154};
ram[6376] = {9'd49,-10'd151};
ram[6377] = {9'd52,-10'd148};
ram[6378] = {9'd55,-10'd145};
ram[6379] = {9'd58,-10'd142};
ram[6380] = {9'd62,-10'd139};
ram[6381] = {9'd65,-10'd136};
ram[6382] = {9'd68,-10'd132};
ram[6383] = {9'd71,-10'd129};
ram[6384] = {9'd74,-10'd126};
ram[6385] = {9'd77,-10'd123};
ram[6386] = {9'd80,-10'd120};
ram[6387] = {9'd84,-10'd117};
ram[6388] = {9'd87,-10'd114};
ram[6389] = {9'd90,-10'd110};
ram[6390] = {9'd93,-10'd107};
ram[6391] = {9'd96,-10'd104};
ram[6392] = {9'd99,-10'd101};
ram[6393] = {-9'd98,-10'd98};
ram[6394] = {-9'd95,-10'd95};
ram[6395] = {-9'd92,-10'd92};
ram[6396] = {-9'd88,-10'd88};
ram[6397] = {-9'd85,-10'd85};
ram[6398] = {-9'd82,-10'd82};
ram[6399] = {-9'd79,-10'd79};
ram[6400] = {-9'd79,-10'd79};
ram[6401] = {-9'd76,-10'd76};
ram[6402] = {-9'd73,-10'd73};
ram[6403] = {-9'd70,-10'd70};
ram[6404] = {-9'd66,-10'd66};
ram[6405] = {-9'd63,-10'd63};
ram[6406] = {-9'd60,-10'd60};
ram[6407] = {-9'd57,-10'd57};
ram[6408] = {-9'd54,-10'd54};
ram[6409] = {-9'd51,-10'd51};
ram[6410] = {-9'd48,-10'd48};
ram[6411] = {-9'd44,-10'd44};
ram[6412] = {-9'd41,-10'd41};
ram[6413] = {-9'd38,-10'd38};
ram[6414] = {-9'd35,-10'd35};
ram[6415] = {-9'd32,-10'd32};
ram[6416] = {-9'd29,-10'd29};
ram[6417] = {-9'd26,-10'd26};
ram[6418] = {-9'd22,-10'd22};
ram[6419] = {-9'd19,-10'd19};
ram[6420] = {-9'd16,-10'd16};
ram[6421] = {-9'd13,-10'd13};
ram[6422] = {-9'd10,-10'd10};
ram[6423] = {-9'd7,-10'd7};
ram[6424] = {-9'd4,-10'd4};
ram[6425] = {9'd0,10'd0};
ram[6426] = {9'd3,10'd3};
ram[6427] = {9'd6,10'd6};
ram[6428] = {9'd9,10'd9};
ram[6429] = {9'd12,10'd12};
ram[6430] = {9'd15,10'd15};
ram[6431] = {9'd18,10'd18};
ram[6432] = {9'd21,10'd21};
ram[6433] = {9'd25,10'd25};
ram[6434] = {9'd28,10'd28};
ram[6435] = {9'd31,10'd31};
ram[6436] = {9'd34,10'd34};
ram[6437] = {9'd37,10'd37};
ram[6438] = {9'd40,10'd40};
ram[6439] = {9'd43,10'd43};
ram[6440] = {9'd47,10'd47};
ram[6441] = {9'd50,10'd50};
ram[6442] = {9'd53,10'd53};
ram[6443] = {9'd56,10'd56};
ram[6444] = {9'd59,10'd59};
ram[6445] = {9'd62,10'd62};
ram[6446] = {9'd65,10'd65};
ram[6447] = {9'd69,10'd69};
ram[6448] = {9'd72,10'd72};
ram[6449] = {9'd75,10'd75};
ram[6450] = {9'd78,10'd78};
ram[6451] = {9'd81,10'd81};
ram[6452] = {9'd84,10'd84};
ram[6453] = {9'd87,10'd87};
ram[6454] = {9'd91,10'd91};
ram[6455] = {9'd94,10'd94};
ram[6456] = {9'd97,10'd97};
ram[6457] = {-9'd100,10'd100};
ram[6458] = {-9'd97,10'd103};
ram[6459] = {-9'd94,10'd106};
ram[6460] = {-9'd91,10'd109};
ram[6461] = {-9'd88,10'd113};
ram[6462] = {-9'd85,10'd116};
ram[6463] = {-9'd81,10'd119};
ram[6464] = {-9'd78,10'd122};
ram[6465] = {-9'd75,10'd125};
ram[6466] = {-9'd72,10'd128};
ram[6467] = {-9'd69,10'd131};
ram[6468] = {-9'd66,10'd135};
ram[6469] = {-9'd63,10'd138};
ram[6470] = {-9'd59,10'd141};
ram[6471] = {-9'd56,10'd144};
ram[6472] = {-9'd53,10'd147};
ram[6473] = {-9'd50,10'd150};
ram[6474] = {-9'd47,10'd153};
ram[6475] = {-9'd44,10'd157};
ram[6476] = {-9'd41,10'd160};
ram[6477] = {-9'd37,10'd163};
ram[6478] = {-9'd34,10'd166};
ram[6479] = {-9'd31,10'd169};
ram[6480] = {-9'd28,10'd172};
ram[6481] = {-9'd25,10'd175};
ram[6482] = {-9'd22,10'd179};
ram[6483] = {-9'd19,10'd182};
ram[6484] = {-9'd15,10'd185};
ram[6485] = {-9'd12,10'd188};
ram[6486] = {-9'd9,10'd191};
ram[6487] = {-9'd6,10'd194};
ram[6488] = {-9'd3,10'd197};
ram[6489] = {9'd0,10'd201};
ram[6490] = {9'd3,10'd204};
ram[6491] = {9'd7,10'd207};
ram[6492] = {9'd10,10'd210};
ram[6493] = {9'd13,10'd213};
ram[6494] = {9'd16,10'd216};
ram[6495] = {9'd19,10'd219};
ram[6496] = {9'd22,10'd223};
ram[6497] = {9'd25,10'd226};
ram[6498] = {9'd29,10'd229};
ram[6499] = {9'd32,10'd232};
ram[6500] = {9'd35,10'd235};
ram[6501] = {9'd38,10'd238};
ram[6502] = {9'd41,10'd241};
ram[6503] = {9'd44,10'd245};
ram[6504] = {9'd47,10'd248};
ram[6505] = {9'd51,10'd251};
ram[6506] = {9'd54,10'd254};
ram[6507] = {9'd57,10'd257};
ram[6508] = {9'd60,10'd260};
ram[6509] = {9'd63,10'd263};
ram[6510] = {9'd66,10'd267};
ram[6511] = {9'd69,10'd270};
ram[6512] = {9'd73,10'd273};
ram[6513] = {9'd76,10'd276};
ram[6514] = {9'd79,10'd279};
ram[6515] = {9'd82,10'd282};
ram[6516] = {9'd85,10'd285};
ram[6517] = {9'd88,10'd289};
ram[6518] = {9'd91,10'd292};
ram[6519] = {9'd95,10'd295};
ram[6520] = {9'd98,10'd298};
ram[6521] = {-9'd99,10'd301};
ram[6522] = {-9'd96,10'd304};
ram[6523] = {-9'd93,10'd307};
ram[6524] = {-9'd90,10'd311};
ram[6525] = {-9'd87,10'd314};
ram[6526] = {-9'd84,10'd317};
ram[6527] = {-9'd81,10'd320};
ram[6528] = {-9'd81,10'd320};
ram[6529] = {-9'd77,10'd323};
ram[6530] = {-9'd74,10'd326};
ram[6531] = {-9'd71,10'd329};
ram[6532] = {-9'd68,10'd333};
ram[6533] = {-9'd65,10'd336};
ram[6534] = {-9'd62,10'd339};
ram[6535] = {-9'd59,10'd342};
ram[6536] = {-9'd55,10'd345};
ram[6537] = {-9'd52,10'd348};
ram[6538] = {-9'd49,10'd351};
ram[6539] = {-9'd46,10'd354};
ram[6540] = {-9'd43,10'd358};
ram[6541] = {-9'd40,10'd361};
ram[6542] = {-9'd37,10'd364};
ram[6543] = {-9'd33,10'd367};
ram[6544] = {-9'd30,10'd370};
ram[6545] = {-9'd27,10'd373};
ram[6546] = {-9'd24,10'd376};
ram[6547] = {-9'd21,10'd380};
ram[6548] = {-9'd18,10'd383};
ram[6549] = {-9'd15,10'd386};
ram[6550] = {-9'd11,10'd389};
ram[6551] = {-9'd8,10'd392};
ram[6552] = {-9'd5,10'd395};
ram[6553] = {-9'd2,10'd398};
ram[6554] = {9'd1,-10'd399};
ram[6555] = {9'd4,-10'd396};
ram[6556] = {9'd7,-10'd393};
ram[6557] = {9'd10,-10'd390};
ram[6558] = {9'd14,-10'd387};
ram[6559] = {9'd17,-10'd384};
ram[6560] = {9'd20,-10'd381};
ram[6561] = {9'd23,-10'd377};
ram[6562] = {9'd26,-10'd374};
ram[6563] = {9'd29,-10'd371};
ram[6564] = {9'd32,-10'd368};
ram[6565] = {9'd36,-10'd365};
ram[6566] = {9'd39,-10'd362};
ram[6567] = {9'd42,-10'd359};
ram[6568] = {9'd45,-10'd355};
ram[6569] = {9'd48,-10'd352};
ram[6570] = {9'd51,-10'd349};
ram[6571] = {9'd54,-10'd346};
ram[6572] = {9'd58,-10'd343};
ram[6573] = {9'd61,-10'd340};
ram[6574] = {9'd64,-10'd337};
ram[6575] = {9'd67,-10'd334};
ram[6576] = {9'd70,-10'd330};
ram[6577] = {9'd73,-10'd327};
ram[6578] = {9'd76,-10'd324};
ram[6579] = {9'd80,-10'd321};
ram[6580] = {9'd83,-10'd318};
ram[6581] = {9'd86,-10'd315};
ram[6582] = {9'd89,-10'd312};
ram[6583] = {9'd92,-10'd308};
ram[6584] = {9'd95,-10'd305};
ram[6585] = {9'd98,-10'd302};
ram[6586] = {-9'd99,-10'd299};
ram[6587] = {-9'd96,-10'd296};
ram[6588] = {-9'd92,-10'd293};
ram[6589] = {-9'd89,-10'd290};
ram[6590] = {-9'd86,-10'd286};
ram[6591] = {-9'd83,-10'd283};
ram[6592] = {-9'd80,-10'd280};
ram[6593] = {-9'd77,-10'd277};
ram[6594] = {-9'd74,-10'd274};
ram[6595] = {-9'd70,-10'd271};
ram[6596] = {-9'd67,-10'd268};
ram[6597] = {-9'd64,-10'd264};
ram[6598] = {-9'd61,-10'd261};
ram[6599] = {-9'd58,-10'd258};
ram[6600] = {-9'd55,-10'd255};
ram[6601] = {-9'd52,-10'd252};
ram[6602] = {-9'd48,-10'd249};
ram[6603] = {-9'd45,-10'd246};
ram[6604] = {-9'd42,-10'd242};
ram[6605] = {-9'd39,-10'd239};
ram[6606] = {-9'd36,-10'd236};
ram[6607] = {-9'd33,-10'd233};
ram[6608] = {-9'd30,-10'd230};
ram[6609] = {-9'd26,-10'd227};
ram[6610] = {-9'd23,-10'd224};
ram[6611] = {-9'd20,-10'd220};
ram[6612] = {-9'd17,-10'd217};
ram[6613] = {-9'd14,-10'd214};
ram[6614] = {-9'd11,-10'd211};
ram[6615] = {-9'd8,-10'd208};
ram[6616] = {-9'd4,-10'd205};
ram[6617] = {-9'd1,-10'd202};
ram[6618] = {9'd2,-10'd198};
ram[6619] = {9'd5,-10'd195};
ram[6620] = {9'd8,-10'd192};
ram[6621] = {9'd11,-10'd189};
ram[6622] = {9'd14,-10'd186};
ram[6623] = {9'd18,-10'd183};
ram[6624] = {9'd21,-10'd180};
ram[6625] = {9'd24,-10'd176};
ram[6626] = {9'd27,-10'd173};
ram[6627] = {9'd30,-10'd170};
ram[6628] = {9'd33,-10'd167};
ram[6629] = {9'd36,-10'd164};
ram[6630] = {9'd40,-10'd161};
ram[6631] = {9'd43,-10'd158};
ram[6632] = {9'd46,-10'd154};
ram[6633] = {9'd49,-10'd151};
ram[6634] = {9'd52,-10'd148};
ram[6635] = {9'd55,-10'd145};
ram[6636] = {9'd58,-10'd142};
ram[6637] = {9'd62,-10'd139};
ram[6638] = {9'd65,-10'd136};
ram[6639] = {9'd68,-10'd132};
ram[6640] = {9'd71,-10'd129};
ram[6641] = {9'd74,-10'd126};
ram[6642] = {9'd77,-10'd123};
ram[6643] = {9'd80,-10'd120};
ram[6644] = {9'd84,-10'd117};
ram[6645] = {9'd87,-10'd114};
ram[6646] = {9'd90,-10'd110};
ram[6647] = {9'd93,-10'd107};
ram[6648] = {9'd96,-10'd104};
ram[6649] = {9'd99,-10'd101};
ram[6650] = {-9'd98,-10'd98};
ram[6651] = {-9'd95,-10'd95};
ram[6652] = {-9'd92,-10'd92};
ram[6653] = {-9'd88,-10'd88};
ram[6654] = {-9'd85,-10'd85};
ram[6655] = {-9'd82,-10'd82};
ram[6656] = {-9'd82,-10'd82};
ram[6657] = {-9'd79,-10'd79};
ram[6658] = {-9'd76,-10'd76};
ram[6659] = {-9'd73,-10'd73};
ram[6660] = {-9'd70,-10'd70};
ram[6661] = {-9'd66,-10'd66};
ram[6662] = {-9'd63,-10'd63};
ram[6663] = {-9'd60,-10'd60};
ram[6664] = {-9'd57,-10'd57};
ram[6665] = {-9'd54,-10'd54};
ram[6666] = {-9'd51,-10'd51};
ram[6667] = {-9'd48,-10'd48};
ram[6668] = {-9'd44,-10'd44};
ram[6669] = {-9'd41,-10'd41};
ram[6670] = {-9'd38,-10'd38};
ram[6671] = {-9'd35,-10'd35};
ram[6672] = {-9'd32,-10'd32};
ram[6673] = {-9'd29,-10'd29};
ram[6674] = {-9'd26,-10'd26};
ram[6675] = {-9'd22,-10'd22};
ram[6676] = {-9'd19,-10'd19};
ram[6677] = {-9'd16,-10'd16};
ram[6678] = {-9'd13,-10'd13};
ram[6679] = {-9'd10,-10'd10};
ram[6680] = {-9'd7,-10'd7};
ram[6681] = {-9'd4,-10'd4};
ram[6682] = {9'd0,10'd0};
ram[6683] = {9'd3,10'd3};
ram[6684] = {9'd6,10'd6};
ram[6685] = {9'd9,10'd9};
ram[6686] = {9'd12,10'd12};
ram[6687] = {9'd15,10'd15};
ram[6688] = {9'd18,10'd18};
ram[6689] = {9'd21,10'd21};
ram[6690] = {9'd25,10'd25};
ram[6691] = {9'd28,10'd28};
ram[6692] = {9'd31,10'd31};
ram[6693] = {9'd34,10'd34};
ram[6694] = {9'd37,10'd37};
ram[6695] = {9'd40,10'd40};
ram[6696] = {9'd43,10'd43};
ram[6697] = {9'd47,10'd47};
ram[6698] = {9'd50,10'd50};
ram[6699] = {9'd53,10'd53};
ram[6700] = {9'd56,10'd56};
ram[6701] = {9'd59,10'd59};
ram[6702] = {9'd62,10'd62};
ram[6703] = {9'd65,10'd65};
ram[6704] = {9'd69,10'd69};
ram[6705] = {9'd72,10'd72};
ram[6706] = {9'd75,10'd75};
ram[6707] = {9'd78,10'd78};
ram[6708] = {9'd81,10'd81};
ram[6709] = {9'd84,10'd84};
ram[6710] = {9'd87,10'd87};
ram[6711] = {9'd91,10'd91};
ram[6712] = {9'd94,10'd94};
ram[6713] = {9'd97,10'd97};
ram[6714] = {-9'd100,10'd100};
ram[6715] = {-9'd97,10'd103};
ram[6716] = {-9'd94,10'd106};
ram[6717] = {-9'd91,10'd109};
ram[6718] = {-9'd88,10'd113};
ram[6719] = {-9'd85,10'd116};
ram[6720] = {-9'd81,10'd119};
ram[6721] = {-9'd78,10'd122};
ram[6722] = {-9'd75,10'd125};
ram[6723] = {-9'd72,10'd128};
ram[6724] = {-9'd69,10'd131};
ram[6725] = {-9'd66,10'd135};
ram[6726] = {-9'd63,10'd138};
ram[6727] = {-9'd59,10'd141};
ram[6728] = {-9'd56,10'd144};
ram[6729] = {-9'd53,10'd147};
ram[6730] = {-9'd50,10'd150};
ram[6731] = {-9'd47,10'd153};
ram[6732] = {-9'd44,10'd157};
ram[6733] = {-9'd41,10'd160};
ram[6734] = {-9'd37,10'd163};
ram[6735] = {-9'd34,10'd166};
ram[6736] = {-9'd31,10'd169};
ram[6737] = {-9'd28,10'd172};
ram[6738] = {-9'd25,10'd175};
ram[6739] = {-9'd22,10'd179};
ram[6740] = {-9'd19,10'd182};
ram[6741] = {-9'd15,10'd185};
ram[6742] = {-9'd12,10'd188};
ram[6743] = {-9'd9,10'd191};
ram[6744] = {-9'd6,10'd194};
ram[6745] = {-9'd3,10'd197};
ram[6746] = {9'd0,10'd201};
ram[6747] = {9'd3,10'd204};
ram[6748] = {9'd7,10'd207};
ram[6749] = {9'd10,10'd210};
ram[6750] = {9'd13,10'd213};
ram[6751] = {9'd16,10'd216};
ram[6752] = {9'd19,10'd219};
ram[6753] = {9'd22,10'd223};
ram[6754] = {9'd25,10'd226};
ram[6755] = {9'd29,10'd229};
ram[6756] = {9'd32,10'd232};
ram[6757] = {9'd35,10'd235};
ram[6758] = {9'd38,10'd238};
ram[6759] = {9'd41,10'd241};
ram[6760] = {9'd44,10'd245};
ram[6761] = {9'd47,10'd248};
ram[6762] = {9'd51,10'd251};
ram[6763] = {9'd54,10'd254};
ram[6764] = {9'd57,10'd257};
ram[6765] = {9'd60,10'd260};
ram[6766] = {9'd63,10'd263};
ram[6767] = {9'd66,10'd267};
ram[6768] = {9'd69,10'd270};
ram[6769] = {9'd73,10'd273};
ram[6770] = {9'd76,10'd276};
ram[6771] = {9'd79,10'd279};
ram[6772] = {9'd82,10'd282};
ram[6773] = {9'd85,10'd285};
ram[6774] = {9'd88,10'd289};
ram[6775] = {9'd91,10'd292};
ram[6776] = {9'd95,10'd295};
ram[6777] = {9'd98,10'd298};
ram[6778] = {-9'd99,10'd301};
ram[6779] = {-9'd96,10'd304};
ram[6780] = {-9'd93,10'd307};
ram[6781] = {-9'd90,10'd311};
ram[6782] = {-9'd87,10'd314};
ram[6783] = {-9'd84,10'd317};
ram[6784] = {-9'd84,10'd317};
ram[6785] = {-9'd81,10'd320};
ram[6786] = {-9'd77,10'd323};
ram[6787] = {-9'd74,10'd326};
ram[6788] = {-9'd71,10'd329};
ram[6789] = {-9'd68,10'd333};
ram[6790] = {-9'd65,10'd336};
ram[6791] = {-9'd62,10'd339};
ram[6792] = {-9'd59,10'd342};
ram[6793] = {-9'd55,10'd345};
ram[6794] = {-9'd52,10'd348};
ram[6795] = {-9'd49,10'd351};
ram[6796] = {-9'd46,10'd354};
ram[6797] = {-9'd43,10'd358};
ram[6798] = {-9'd40,10'd361};
ram[6799] = {-9'd37,10'd364};
ram[6800] = {-9'd33,10'd367};
ram[6801] = {-9'd30,10'd370};
ram[6802] = {-9'd27,10'd373};
ram[6803] = {-9'd24,10'd376};
ram[6804] = {-9'd21,10'd380};
ram[6805] = {-9'd18,10'd383};
ram[6806] = {-9'd15,10'd386};
ram[6807] = {-9'd11,10'd389};
ram[6808] = {-9'd8,10'd392};
ram[6809] = {-9'd5,10'd395};
ram[6810] = {-9'd2,10'd398};
ram[6811] = {9'd1,-10'd399};
ram[6812] = {9'd4,-10'd396};
ram[6813] = {9'd7,-10'd393};
ram[6814] = {9'd10,-10'd390};
ram[6815] = {9'd14,-10'd387};
ram[6816] = {9'd17,-10'd384};
ram[6817] = {9'd20,-10'd381};
ram[6818] = {9'd23,-10'd377};
ram[6819] = {9'd26,-10'd374};
ram[6820] = {9'd29,-10'd371};
ram[6821] = {9'd32,-10'd368};
ram[6822] = {9'd36,-10'd365};
ram[6823] = {9'd39,-10'd362};
ram[6824] = {9'd42,-10'd359};
ram[6825] = {9'd45,-10'd355};
ram[6826] = {9'd48,-10'd352};
ram[6827] = {9'd51,-10'd349};
ram[6828] = {9'd54,-10'd346};
ram[6829] = {9'd58,-10'd343};
ram[6830] = {9'd61,-10'd340};
ram[6831] = {9'd64,-10'd337};
ram[6832] = {9'd67,-10'd334};
ram[6833] = {9'd70,-10'd330};
ram[6834] = {9'd73,-10'd327};
ram[6835] = {9'd76,-10'd324};
ram[6836] = {9'd80,-10'd321};
ram[6837] = {9'd83,-10'd318};
ram[6838] = {9'd86,-10'd315};
ram[6839] = {9'd89,-10'd312};
ram[6840] = {9'd92,-10'd308};
ram[6841] = {9'd95,-10'd305};
ram[6842] = {9'd98,-10'd302};
ram[6843] = {-9'd99,-10'd299};
ram[6844] = {-9'd96,-10'd296};
ram[6845] = {-9'd92,-10'd293};
ram[6846] = {-9'd89,-10'd290};
ram[6847] = {-9'd86,-10'd286};
ram[6848] = {-9'd83,-10'd283};
ram[6849] = {-9'd80,-10'd280};
ram[6850] = {-9'd77,-10'd277};
ram[6851] = {-9'd74,-10'd274};
ram[6852] = {-9'd70,-10'd271};
ram[6853] = {-9'd67,-10'd268};
ram[6854] = {-9'd64,-10'd264};
ram[6855] = {-9'd61,-10'd261};
ram[6856] = {-9'd58,-10'd258};
ram[6857] = {-9'd55,-10'd255};
ram[6858] = {-9'd52,-10'd252};
ram[6859] = {-9'd48,-10'd249};
ram[6860] = {-9'd45,-10'd246};
ram[6861] = {-9'd42,-10'd242};
ram[6862] = {-9'd39,-10'd239};
ram[6863] = {-9'd36,-10'd236};
ram[6864] = {-9'd33,-10'd233};
ram[6865] = {-9'd30,-10'd230};
ram[6866] = {-9'd26,-10'd227};
ram[6867] = {-9'd23,-10'd224};
ram[6868] = {-9'd20,-10'd220};
ram[6869] = {-9'd17,-10'd217};
ram[6870] = {-9'd14,-10'd214};
ram[6871] = {-9'd11,-10'd211};
ram[6872] = {-9'd8,-10'd208};
ram[6873] = {-9'd4,-10'd205};
ram[6874] = {-9'd1,-10'd202};
ram[6875] = {9'd2,-10'd198};
ram[6876] = {9'd5,-10'd195};
ram[6877] = {9'd8,-10'd192};
ram[6878] = {9'd11,-10'd189};
ram[6879] = {9'd14,-10'd186};
ram[6880] = {9'd18,-10'd183};
ram[6881] = {9'd21,-10'd180};
ram[6882] = {9'd24,-10'd176};
ram[6883] = {9'd27,-10'd173};
ram[6884] = {9'd30,-10'd170};
ram[6885] = {9'd33,-10'd167};
ram[6886] = {9'd36,-10'd164};
ram[6887] = {9'd40,-10'd161};
ram[6888] = {9'd43,-10'd158};
ram[6889] = {9'd46,-10'd154};
ram[6890] = {9'd49,-10'd151};
ram[6891] = {9'd52,-10'd148};
ram[6892] = {9'd55,-10'd145};
ram[6893] = {9'd58,-10'd142};
ram[6894] = {9'd62,-10'd139};
ram[6895] = {9'd65,-10'd136};
ram[6896] = {9'd68,-10'd132};
ram[6897] = {9'd71,-10'd129};
ram[6898] = {9'd74,-10'd126};
ram[6899] = {9'd77,-10'd123};
ram[6900] = {9'd80,-10'd120};
ram[6901] = {9'd84,-10'd117};
ram[6902] = {9'd87,-10'd114};
ram[6903] = {9'd90,-10'd110};
ram[6904] = {9'd93,-10'd107};
ram[6905] = {9'd96,-10'd104};
ram[6906] = {9'd99,-10'd101};
ram[6907] = {-9'd98,-10'd98};
ram[6908] = {-9'd95,-10'd95};
ram[6909] = {-9'd92,-10'd92};
ram[6910] = {-9'd88,-10'd88};
ram[6911] = {-9'd85,-10'd85};
ram[6912] = {-9'd85,-10'd85};
ram[6913] = {-9'd82,-10'd82};
ram[6914] = {-9'd79,-10'd79};
ram[6915] = {-9'd76,-10'd76};
ram[6916] = {-9'd73,-10'd73};
ram[6917] = {-9'd70,-10'd70};
ram[6918] = {-9'd66,-10'd66};
ram[6919] = {-9'd63,-10'd63};
ram[6920] = {-9'd60,-10'd60};
ram[6921] = {-9'd57,-10'd57};
ram[6922] = {-9'd54,-10'd54};
ram[6923] = {-9'd51,-10'd51};
ram[6924] = {-9'd48,-10'd48};
ram[6925] = {-9'd44,-10'd44};
ram[6926] = {-9'd41,-10'd41};
ram[6927] = {-9'd38,-10'd38};
ram[6928] = {-9'd35,-10'd35};
ram[6929] = {-9'd32,-10'd32};
ram[6930] = {-9'd29,-10'd29};
ram[6931] = {-9'd26,-10'd26};
ram[6932] = {-9'd22,-10'd22};
ram[6933] = {-9'd19,-10'd19};
ram[6934] = {-9'd16,-10'd16};
ram[6935] = {-9'd13,-10'd13};
ram[6936] = {-9'd10,-10'd10};
ram[6937] = {-9'd7,-10'd7};
ram[6938] = {-9'd4,-10'd4};
ram[6939] = {9'd0,10'd0};
ram[6940] = {9'd3,10'd3};
ram[6941] = {9'd6,10'd6};
ram[6942] = {9'd9,10'd9};
ram[6943] = {9'd12,10'd12};
ram[6944] = {9'd15,10'd15};
ram[6945] = {9'd18,10'd18};
ram[6946] = {9'd21,10'd21};
ram[6947] = {9'd25,10'd25};
ram[6948] = {9'd28,10'd28};
ram[6949] = {9'd31,10'd31};
ram[6950] = {9'd34,10'd34};
ram[6951] = {9'd37,10'd37};
ram[6952] = {9'd40,10'd40};
ram[6953] = {9'd43,10'd43};
ram[6954] = {9'd47,10'd47};
ram[6955] = {9'd50,10'd50};
ram[6956] = {9'd53,10'd53};
ram[6957] = {9'd56,10'd56};
ram[6958] = {9'd59,10'd59};
ram[6959] = {9'd62,10'd62};
ram[6960] = {9'd65,10'd65};
ram[6961] = {9'd69,10'd69};
ram[6962] = {9'd72,10'd72};
ram[6963] = {9'd75,10'd75};
ram[6964] = {9'd78,10'd78};
ram[6965] = {9'd81,10'd81};
ram[6966] = {9'd84,10'd84};
ram[6967] = {9'd87,10'd87};
ram[6968] = {9'd91,10'd91};
ram[6969] = {9'd94,10'd94};
ram[6970] = {9'd97,10'd97};
ram[6971] = {-9'd100,10'd100};
ram[6972] = {-9'd97,10'd103};
ram[6973] = {-9'd94,10'd106};
ram[6974] = {-9'd91,10'd109};
ram[6975] = {-9'd88,10'd113};
ram[6976] = {-9'd85,10'd116};
ram[6977] = {-9'd81,10'd119};
ram[6978] = {-9'd78,10'd122};
ram[6979] = {-9'd75,10'd125};
ram[6980] = {-9'd72,10'd128};
ram[6981] = {-9'd69,10'd131};
ram[6982] = {-9'd66,10'd135};
ram[6983] = {-9'd63,10'd138};
ram[6984] = {-9'd59,10'd141};
ram[6985] = {-9'd56,10'd144};
ram[6986] = {-9'd53,10'd147};
ram[6987] = {-9'd50,10'd150};
ram[6988] = {-9'd47,10'd153};
ram[6989] = {-9'd44,10'd157};
ram[6990] = {-9'd41,10'd160};
ram[6991] = {-9'd37,10'd163};
ram[6992] = {-9'd34,10'd166};
ram[6993] = {-9'd31,10'd169};
ram[6994] = {-9'd28,10'd172};
ram[6995] = {-9'd25,10'd175};
ram[6996] = {-9'd22,10'd179};
ram[6997] = {-9'd19,10'd182};
ram[6998] = {-9'd15,10'd185};
ram[6999] = {-9'd12,10'd188};
ram[7000] = {-9'd9,10'd191};
ram[7001] = {-9'd6,10'd194};
ram[7002] = {-9'd3,10'd197};
ram[7003] = {9'd0,10'd201};
ram[7004] = {9'd3,10'd204};
ram[7005] = {9'd7,10'd207};
ram[7006] = {9'd10,10'd210};
ram[7007] = {9'd13,10'd213};
ram[7008] = {9'd16,10'd216};
ram[7009] = {9'd19,10'd219};
ram[7010] = {9'd22,10'd223};
ram[7011] = {9'd25,10'd226};
ram[7012] = {9'd29,10'd229};
ram[7013] = {9'd32,10'd232};
ram[7014] = {9'd35,10'd235};
ram[7015] = {9'd38,10'd238};
ram[7016] = {9'd41,10'd241};
ram[7017] = {9'd44,10'd245};
ram[7018] = {9'd47,10'd248};
ram[7019] = {9'd51,10'd251};
ram[7020] = {9'd54,10'd254};
ram[7021] = {9'd57,10'd257};
ram[7022] = {9'd60,10'd260};
ram[7023] = {9'd63,10'd263};
ram[7024] = {9'd66,10'd267};
ram[7025] = {9'd69,10'd270};
ram[7026] = {9'd73,10'd273};
ram[7027] = {9'd76,10'd276};
ram[7028] = {9'd79,10'd279};
ram[7029] = {9'd82,10'd282};
ram[7030] = {9'd85,10'd285};
ram[7031] = {9'd88,10'd289};
ram[7032] = {9'd91,10'd292};
ram[7033] = {9'd95,10'd295};
ram[7034] = {9'd98,10'd298};
ram[7035] = {-9'd99,10'd301};
ram[7036] = {-9'd96,10'd304};
ram[7037] = {-9'd93,10'd307};
ram[7038] = {-9'd90,10'd311};
ram[7039] = {-9'd87,10'd314};
ram[7040] = {-9'd87,10'd314};
ram[7041] = {-9'd84,10'd317};
ram[7042] = {-9'd81,10'd320};
ram[7043] = {-9'd77,10'd323};
ram[7044] = {-9'd74,10'd326};
ram[7045] = {-9'd71,10'd329};
ram[7046] = {-9'd68,10'd333};
ram[7047] = {-9'd65,10'd336};
ram[7048] = {-9'd62,10'd339};
ram[7049] = {-9'd59,10'd342};
ram[7050] = {-9'd55,10'd345};
ram[7051] = {-9'd52,10'd348};
ram[7052] = {-9'd49,10'd351};
ram[7053] = {-9'd46,10'd354};
ram[7054] = {-9'd43,10'd358};
ram[7055] = {-9'd40,10'd361};
ram[7056] = {-9'd37,10'd364};
ram[7057] = {-9'd33,10'd367};
ram[7058] = {-9'd30,10'd370};
ram[7059] = {-9'd27,10'd373};
ram[7060] = {-9'd24,10'd376};
ram[7061] = {-9'd21,10'd380};
ram[7062] = {-9'd18,10'd383};
ram[7063] = {-9'd15,10'd386};
ram[7064] = {-9'd11,10'd389};
ram[7065] = {-9'd8,10'd392};
ram[7066] = {-9'd5,10'd395};
ram[7067] = {-9'd2,10'd398};
ram[7068] = {9'd1,-10'd399};
ram[7069] = {9'd4,-10'd396};
ram[7070] = {9'd7,-10'd393};
ram[7071] = {9'd10,-10'd390};
ram[7072] = {9'd14,-10'd387};
ram[7073] = {9'd17,-10'd384};
ram[7074] = {9'd20,-10'd381};
ram[7075] = {9'd23,-10'd377};
ram[7076] = {9'd26,-10'd374};
ram[7077] = {9'd29,-10'd371};
ram[7078] = {9'd32,-10'd368};
ram[7079] = {9'd36,-10'd365};
ram[7080] = {9'd39,-10'd362};
ram[7081] = {9'd42,-10'd359};
ram[7082] = {9'd45,-10'd355};
ram[7083] = {9'd48,-10'd352};
ram[7084] = {9'd51,-10'd349};
ram[7085] = {9'd54,-10'd346};
ram[7086] = {9'd58,-10'd343};
ram[7087] = {9'd61,-10'd340};
ram[7088] = {9'd64,-10'd337};
ram[7089] = {9'd67,-10'd334};
ram[7090] = {9'd70,-10'd330};
ram[7091] = {9'd73,-10'd327};
ram[7092] = {9'd76,-10'd324};
ram[7093] = {9'd80,-10'd321};
ram[7094] = {9'd83,-10'd318};
ram[7095] = {9'd86,-10'd315};
ram[7096] = {9'd89,-10'd312};
ram[7097] = {9'd92,-10'd308};
ram[7098] = {9'd95,-10'd305};
ram[7099] = {9'd98,-10'd302};
ram[7100] = {-9'd99,-10'd299};
ram[7101] = {-9'd96,-10'd296};
ram[7102] = {-9'd92,-10'd293};
ram[7103] = {-9'd89,-10'd290};
ram[7104] = {-9'd86,-10'd286};
ram[7105] = {-9'd83,-10'd283};
ram[7106] = {-9'd80,-10'd280};
ram[7107] = {-9'd77,-10'd277};
ram[7108] = {-9'd74,-10'd274};
ram[7109] = {-9'd70,-10'd271};
ram[7110] = {-9'd67,-10'd268};
ram[7111] = {-9'd64,-10'd264};
ram[7112] = {-9'd61,-10'd261};
ram[7113] = {-9'd58,-10'd258};
ram[7114] = {-9'd55,-10'd255};
ram[7115] = {-9'd52,-10'd252};
ram[7116] = {-9'd48,-10'd249};
ram[7117] = {-9'd45,-10'd246};
ram[7118] = {-9'd42,-10'd242};
ram[7119] = {-9'd39,-10'd239};
ram[7120] = {-9'd36,-10'd236};
ram[7121] = {-9'd33,-10'd233};
ram[7122] = {-9'd30,-10'd230};
ram[7123] = {-9'd26,-10'd227};
ram[7124] = {-9'd23,-10'd224};
ram[7125] = {-9'd20,-10'd220};
ram[7126] = {-9'd17,-10'd217};
ram[7127] = {-9'd14,-10'd214};
ram[7128] = {-9'd11,-10'd211};
ram[7129] = {-9'd8,-10'd208};
ram[7130] = {-9'd4,-10'd205};
ram[7131] = {-9'd1,-10'd202};
ram[7132] = {9'd2,-10'd198};
ram[7133] = {9'd5,-10'd195};
ram[7134] = {9'd8,-10'd192};
ram[7135] = {9'd11,-10'd189};
ram[7136] = {9'd14,-10'd186};
ram[7137] = {9'd18,-10'd183};
ram[7138] = {9'd21,-10'd180};
ram[7139] = {9'd24,-10'd176};
ram[7140] = {9'd27,-10'd173};
ram[7141] = {9'd30,-10'd170};
ram[7142] = {9'd33,-10'd167};
ram[7143] = {9'd36,-10'd164};
ram[7144] = {9'd40,-10'd161};
ram[7145] = {9'd43,-10'd158};
ram[7146] = {9'd46,-10'd154};
ram[7147] = {9'd49,-10'd151};
ram[7148] = {9'd52,-10'd148};
ram[7149] = {9'd55,-10'd145};
ram[7150] = {9'd58,-10'd142};
ram[7151] = {9'd62,-10'd139};
ram[7152] = {9'd65,-10'd136};
ram[7153] = {9'd68,-10'd132};
ram[7154] = {9'd71,-10'd129};
ram[7155] = {9'd74,-10'd126};
ram[7156] = {9'd77,-10'd123};
ram[7157] = {9'd80,-10'd120};
ram[7158] = {9'd84,-10'd117};
ram[7159] = {9'd87,-10'd114};
ram[7160] = {9'd90,-10'd110};
ram[7161] = {9'd93,-10'd107};
ram[7162] = {9'd96,-10'd104};
ram[7163] = {9'd99,-10'd101};
ram[7164] = {-9'd98,-10'd98};
ram[7165] = {-9'd95,-10'd95};
ram[7166] = {-9'd92,-10'd92};
ram[7167] = {-9'd88,-10'd88};
ram[7168] = {-9'd88,-10'd88};
ram[7169] = {-9'd85,-10'd85};
ram[7170] = {-9'd82,-10'd82};
ram[7171] = {-9'd79,-10'd79};
ram[7172] = {-9'd76,-10'd76};
ram[7173] = {-9'd73,-10'd73};
ram[7174] = {-9'd70,-10'd70};
ram[7175] = {-9'd66,-10'd66};
ram[7176] = {-9'd63,-10'd63};
ram[7177] = {-9'd60,-10'd60};
ram[7178] = {-9'd57,-10'd57};
ram[7179] = {-9'd54,-10'd54};
ram[7180] = {-9'd51,-10'd51};
ram[7181] = {-9'd48,-10'd48};
ram[7182] = {-9'd44,-10'd44};
ram[7183] = {-9'd41,-10'd41};
ram[7184] = {-9'd38,-10'd38};
ram[7185] = {-9'd35,-10'd35};
ram[7186] = {-9'd32,-10'd32};
ram[7187] = {-9'd29,-10'd29};
ram[7188] = {-9'd26,-10'd26};
ram[7189] = {-9'd22,-10'd22};
ram[7190] = {-9'd19,-10'd19};
ram[7191] = {-9'd16,-10'd16};
ram[7192] = {-9'd13,-10'd13};
ram[7193] = {-9'd10,-10'd10};
ram[7194] = {-9'd7,-10'd7};
ram[7195] = {-9'd4,-10'd4};
ram[7196] = {9'd0,10'd0};
ram[7197] = {9'd3,10'd3};
ram[7198] = {9'd6,10'd6};
ram[7199] = {9'd9,10'd9};
ram[7200] = {9'd12,10'd12};
ram[7201] = {9'd15,10'd15};
ram[7202] = {9'd18,10'd18};
ram[7203] = {9'd21,10'd21};
ram[7204] = {9'd25,10'd25};
ram[7205] = {9'd28,10'd28};
ram[7206] = {9'd31,10'd31};
ram[7207] = {9'd34,10'd34};
ram[7208] = {9'd37,10'd37};
ram[7209] = {9'd40,10'd40};
ram[7210] = {9'd43,10'd43};
ram[7211] = {9'd47,10'd47};
ram[7212] = {9'd50,10'd50};
ram[7213] = {9'd53,10'd53};
ram[7214] = {9'd56,10'd56};
ram[7215] = {9'd59,10'd59};
ram[7216] = {9'd62,10'd62};
ram[7217] = {9'd65,10'd65};
ram[7218] = {9'd69,10'd69};
ram[7219] = {9'd72,10'd72};
ram[7220] = {9'd75,10'd75};
ram[7221] = {9'd78,10'd78};
ram[7222] = {9'd81,10'd81};
ram[7223] = {9'd84,10'd84};
ram[7224] = {9'd87,10'd87};
ram[7225] = {9'd91,10'd91};
ram[7226] = {9'd94,10'd94};
ram[7227] = {9'd97,10'd97};
ram[7228] = {-9'd100,10'd100};
ram[7229] = {-9'd97,10'd103};
ram[7230] = {-9'd94,10'd106};
ram[7231] = {-9'd91,10'd109};
ram[7232] = {-9'd88,10'd113};
ram[7233] = {-9'd85,10'd116};
ram[7234] = {-9'd81,10'd119};
ram[7235] = {-9'd78,10'd122};
ram[7236] = {-9'd75,10'd125};
ram[7237] = {-9'd72,10'd128};
ram[7238] = {-9'd69,10'd131};
ram[7239] = {-9'd66,10'd135};
ram[7240] = {-9'd63,10'd138};
ram[7241] = {-9'd59,10'd141};
ram[7242] = {-9'd56,10'd144};
ram[7243] = {-9'd53,10'd147};
ram[7244] = {-9'd50,10'd150};
ram[7245] = {-9'd47,10'd153};
ram[7246] = {-9'd44,10'd157};
ram[7247] = {-9'd41,10'd160};
ram[7248] = {-9'd37,10'd163};
ram[7249] = {-9'd34,10'd166};
ram[7250] = {-9'd31,10'd169};
ram[7251] = {-9'd28,10'd172};
ram[7252] = {-9'd25,10'd175};
ram[7253] = {-9'd22,10'd179};
ram[7254] = {-9'd19,10'd182};
ram[7255] = {-9'd15,10'd185};
ram[7256] = {-9'd12,10'd188};
ram[7257] = {-9'd9,10'd191};
ram[7258] = {-9'd6,10'd194};
ram[7259] = {-9'd3,10'd197};
ram[7260] = {9'd0,10'd201};
ram[7261] = {9'd3,10'd204};
ram[7262] = {9'd7,10'd207};
ram[7263] = {9'd10,10'd210};
ram[7264] = {9'd13,10'd213};
ram[7265] = {9'd16,10'd216};
ram[7266] = {9'd19,10'd219};
ram[7267] = {9'd22,10'd223};
ram[7268] = {9'd25,10'd226};
ram[7269] = {9'd29,10'd229};
ram[7270] = {9'd32,10'd232};
ram[7271] = {9'd35,10'd235};
ram[7272] = {9'd38,10'd238};
ram[7273] = {9'd41,10'd241};
ram[7274] = {9'd44,10'd245};
ram[7275] = {9'd47,10'd248};
ram[7276] = {9'd51,10'd251};
ram[7277] = {9'd54,10'd254};
ram[7278] = {9'd57,10'd257};
ram[7279] = {9'd60,10'd260};
ram[7280] = {9'd63,10'd263};
ram[7281] = {9'd66,10'd267};
ram[7282] = {9'd69,10'd270};
ram[7283] = {9'd73,10'd273};
ram[7284] = {9'd76,10'd276};
ram[7285] = {9'd79,10'd279};
ram[7286] = {9'd82,10'd282};
ram[7287] = {9'd85,10'd285};
ram[7288] = {9'd88,10'd289};
ram[7289] = {9'd91,10'd292};
ram[7290] = {9'd95,10'd295};
ram[7291] = {9'd98,10'd298};
ram[7292] = {-9'd99,10'd301};
ram[7293] = {-9'd96,10'd304};
ram[7294] = {-9'd93,10'd307};
ram[7295] = {-9'd90,10'd311};
ram[7296] = {-9'd90,10'd311};
ram[7297] = {-9'd87,10'd314};
ram[7298] = {-9'd84,10'd317};
ram[7299] = {-9'd81,10'd320};
ram[7300] = {-9'd77,10'd323};
ram[7301] = {-9'd74,10'd326};
ram[7302] = {-9'd71,10'd329};
ram[7303] = {-9'd68,10'd333};
ram[7304] = {-9'd65,10'd336};
ram[7305] = {-9'd62,10'd339};
ram[7306] = {-9'd59,10'd342};
ram[7307] = {-9'd55,10'd345};
ram[7308] = {-9'd52,10'd348};
ram[7309] = {-9'd49,10'd351};
ram[7310] = {-9'd46,10'd354};
ram[7311] = {-9'd43,10'd358};
ram[7312] = {-9'd40,10'd361};
ram[7313] = {-9'd37,10'd364};
ram[7314] = {-9'd33,10'd367};
ram[7315] = {-9'd30,10'd370};
ram[7316] = {-9'd27,10'd373};
ram[7317] = {-9'd24,10'd376};
ram[7318] = {-9'd21,10'd380};
ram[7319] = {-9'd18,10'd383};
ram[7320] = {-9'd15,10'd386};
ram[7321] = {-9'd11,10'd389};
ram[7322] = {-9'd8,10'd392};
ram[7323] = {-9'd5,10'd395};
ram[7324] = {-9'd2,10'd398};
ram[7325] = {9'd1,-10'd399};
ram[7326] = {9'd4,-10'd396};
ram[7327] = {9'd7,-10'd393};
ram[7328] = {9'd10,-10'd390};
ram[7329] = {9'd14,-10'd387};
ram[7330] = {9'd17,-10'd384};
ram[7331] = {9'd20,-10'd381};
ram[7332] = {9'd23,-10'd377};
ram[7333] = {9'd26,-10'd374};
ram[7334] = {9'd29,-10'd371};
ram[7335] = {9'd32,-10'd368};
ram[7336] = {9'd36,-10'd365};
ram[7337] = {9'd39,-10'd362};
ram[7338] = {9'd42,-10'd359};
ram[7339] = {9'd45,-10'd355};
ram[7340] = {9'd48,-10'd352};
ram[7341] = {9'd51,-10'd349};
ram[7342] = {9'd54,-10'd346};
ram[7343] = {9'd58,-10'd343};
ram[7344] = {9'd61,-10'd340};
ram[7345] = {9'd64,-10'd337};
ram[7346] = {9'd67,-10'd334};
ram[7347] = {9'd70,-10'd330};
ram[7348] = {9'd73,-10'd327};
ram[7349] = {9'd76,-10'd324};
ram[7350] = {9'd80,-10'd321};
ram[7351] = {9'd83,-10'd318};
ram[7352] = {9'd86,-10'd315};
ram[7353] = {9'd89,-10'd312};
ram[7354] = {9'd92,-10'd308};
ram[7355] = {9'd95,-10'd305};
ram[7356] = {9'd98,-10'd302};
ram[7357] = {-9'd99,-10'd299};
ram[7358] = {-9'd96,-10'd296};
ram[7359] = {-9'd92,-10'd293};
ram[7360] = {-9'd89,-10'd290};
ram[7361] = {-9'd86,-10'd286};
ram[7362] = {-9'd83,-10'd283};
ram[7363] = {-9'd80,-10'd280};
ram[7364] = {-9'd77,-10'd277};
ram[7365] = {-9'd74,-10'd274};
ram[7366] = {-9'd70,-10'd271};
ram[7367] = {-9'd67,-10'd268};
ram[7368] = {-9'd64,-10'd264};
ram[7369] = {-9'd61,-10'd261};
ram[7370] = {-9'd58,-10'd258};
ram[7371] = {-9'd55,-10'd255};
ram[7372] = {-9'd52,-10'd252};
ram[7373] = {-9'd48,-10'd249};
ram[7374] = {-9'd45,-10'd246};
ram[7375] = {-9'd42,-10'd242};
ram[7376] = {-9'd39,-10'd239};
ram[7377] = {-9'd36,-10'd236};
ram[7378] = {-9'd33,-10'd233};
ram[7379] = {-9'd30,-10'd230};
ram[7380] = {-9'd26,-10'd227};
ram[7381] = {-9'd23,-10'd224};
ram[7382] = {-9'd20,-10'd220};
ram[7383] = {-9'd17,-10'd217};
ram[7384] = {-9'd14,-10'd214};
ram[7385] = {-9'd11,-10'd211};
ram[7386] = {-9'd8,-10'd208};
ram[7387] = {-9'd4,-10'd205};
ram[7388] = {-9'd1,-10'd202};
ram[7389] = {9'd2,-10'd198};
ram[7390] = {9'd5,-10'd195};
ram[7391] = {9'd8,-10'd192};
ram[7392] = {9'd11,-10'd189};
ram[7393] = {9'd14,-10'd186};
ram[7394] = {9'd18,-10'd183};
ram[7395] = {9'd21,-10'd180};
ram[7396] = {9'd24,-10'd176};
ram[7397] = {9'd27,-10'd173};
ram[7398] = {9'd30,-10'd170};
ram[7399] = {9'd33,-10'd167};
ram[7400] = {9'd36,-10'd164};
ram[7401] = {9'd40,-10'd161};
ram[7402] = {9'd43,-10'd158};
ram[7403] = {9'd46,-10'd154};
ram[7404] = {9'd49,-10'd151};
ram[7405] = {9'd52,-10'd148};
ram[7406] = {9'd55,-10'd145};
ram[7407] = {9'd58,-10'd142};
ram[7408] = {9'd62,-10'd139};
ram[7409] = {9'd65,-10'd136};
ram[7410] = {9'd68,-10'd132};
ram[7411] = {9'd71,-10'd129};
ram[7412] = {9'd74,-10'd126};
ram[7413] = {9'd77,-10'd123};
ram[7414] = {9'd80,-10'd120};
ram[7415] = {9'd84,-10'd117};
ram[7416] = {9'd87,-10'd114};
ram[7417] = {9'd90,-10'd110};
ram[7418] = {9'd93,-10'd107};
ram[7419] = {9'd96,-10'd104};
ram[7420] = {9'd99,-10'd101};
ram[7421] = {-9'd98,-10'd98};
ram[7422] = {-9'd95,-10'd95};
ram[7423] = {-9'd92,-10'd92};
ram[7424] = {-9'd92,-10'd92};
ram[7425] = {-9'd88,-10'd88};
ram[7426] = {-9'd85,-10'd85};
ram[7427] = {-9'd82,-10'd82};
ram[7428] = {-9'd79,-10'd79};
ram[7429] = {-9'd76,-10'd76};
ram[7430] = {-9'd73,-10'd73};
ram[7431] = {-9'd70,-10'd70};
ram[7432] = {-9'd66,-10'd66};
ram[7433] = {-9'd63,-10'd63};
ram[7434] = {-9'd60,-10'd60};
ram[7435] = {-9'd57,-10'd57};
ram[7436] = {-9'd54,-10'd54};
ram[7437] = {-9'd51,-10'd51};
ram[7438] = {-9'd48,-10'd48};
ram[7439] = {-9'd44,-10'd44};
ram[7440] = {-9'd41,-10'd41};
ram[7441] = {-9'd38,-10'd38};
ram[7442] = {-9'd35,-10'd35};
ram[7443] = {-9'd32,-10'd32};
ram[7444] = {-9'd29,-10'd29};
ram[7445] = {-9'd26,-10'd26};
ram[7446] = {-9'd22,-10'd22};
ram[7447] = {-9'd19,-10'd19};
ram[7448] = {-9'd16,-10'd16};
ram[7449] = {-9'd13,-10'd13};
ram[7450] = {-9'd10,-10'd10};
ram[7451] = {-9'd7,-10'd7};
ram[7452] = {-9'd4,-10'd4};
ram[7453] = {9'd0,10'd0};
ram[7454] = {9'd3,10'd3};
ram[7455] = {9'd6,10'd6};
ram[7456] = {9'd9,10'd9};
ram[7457] = {9'd12,10'd12};
ram[7458] = {9'd15,10'd15};
ram[7459] = {9'd18,10'd18};
ram[7460] = {9'd21,10'd21};
ram[7461] = {9'd25,10'd25};
ram[7462] = {9'd28,10'd28};
ram[7463] = {9'd31,10'd31};
ram[7464] = {9'd34,10'd34};
ram[7465] = {9'd37,10'd37};
ram[7466] = {9'd40,10'd40};
ram[7467] = {9'd43,10'd43};
ram[7468] = {9'd47,10'd47};
ram[7469] = {9'd50,10'd50};
ram[7470] = {9'd53,10'd53};
ram[7471] = {9'd56,10'd56};
ram[7472] = {9'd59,10'd59};
ram[7473] = {9'd62,10'd62};
ram[7474] = {9'd65,10'd65};
ram[7475] = {9'd69,10'd69};
ram[7476] = {9'd72,10'd72};
ram[7477] = {9'd75,10'd75};
ram[7478] = {9'd78,10'd78};
ram[7479] = {9'd81,10'd81};
ram[7480] = {9'd84,10'd84};
ram[7481] = {9'd87,10'd87};
ram[7482] = {9'd91,10'd91};
ram[7483] = {9'd94,10'd94};
ram[7484] = {9'd97,10'd97};
ram[7485] = {-9'd100,10'd100};
ram[7486] = {-9'd97,10'd103};
ram[7487] = {-9'd94,10'd106};
ram[7488] = {-9'd91,10'd109};
ram[7489] = {-9'd88,10'd113};
ram[7490] = {-9'd85,10'd116};
ram[7491] = {-9'd81,10'd119};
ram[7492] = {-9'd78,10'd122};
ram[7493] = {-9'd75,10'd125};
ram[7494] = {-9'd72,10'd128};
ram[7495] = {-9'd69,10'd131};
ram[7496] = {-9'd66,10'd135};
ram[7497] = {-9'd63,10'd138};
ram[7498] = {-9'd59,10'd141};
ram[7499] = {-9'd56,10'd144};
ram[7500] = {-9'd53,10'd147};
ram[7501] = {-9'd50,10'd150};
ram[7502] = {-9'd47,10'd153};
ram[7503] = {-9'd44,10'd157};
ram[7504] = {-9'd41,10'd160};
ram[7505] = {-9'd37,10'd163};
ram[7506] = {-9'd34,10'd166};
ram[7507] = {-9'd31,10'd169};
ram[7508] = {-9'd28,10'd172};
ram[7509] = {-9'd25,10'd175};
ram[7510] = {-9'd22,10'd179};
ram[7511] = {-9'd19,10'd182};
ram[7512] = {-9'd15,10'd185};
ram[7513] = {-9'd12,10'd188};
ram[7514] = {-9'd9,10'd191};
ram[7515] = {-9'd6,10'd194};
ram[7516] = {-9'd3,10'd197};
ram[7517] = {9'd0,10'd201};
ram[7518] = {9'd3,10'd204};
ram[7519] = {9'd7,10'd207};
ram[7520] = {9'd10,10'd210};
ram[7521] = {9'd13,10'd213};
ram[7522] = {9'd16,10'd216};
ram[7523] = {9'd19,10'd219};
ram[7524] = {9'd22,10'd223};
ram[7525] = {9'd25,10'd226};
ram[7526] = {9'd29,10'd229};
ram[7527] = {9'd32,10'd232};
ram[7528] = {9'd35,10'd235};
ram[7529] = {9'd38,10'd238};
ram[7530] = {9'd41,10'd241};
ram[7531] = {9'd44,10'd245};
ram[7532] = {9'd47,10'd248};
ram[7533] = {9'd51,10'd251};
ram[7534] = {9'd54,10'd254};
ram[7535] = {9'd57,10'd257};
ram[7536] = {9'd60,10'd260};
ram[7537] = {9'd63,10'd263};
ram[7538] = {9'd66,10'd267};
ram[7539] = {9'd69,10'd270};
ram[7540] = {9'd73,10'd273};
ram[7541] = {9'd76,10'd276};
ram[7542] = {9'd79,10'd279};
ram[7543] = {9'd82,10'd282};
ram[7544] = {9'd85,10'd285};
ram[7545] = {9'd88,10'd289};
ram[7546] = {9'd91,10'd292};
ram[7547] = {9'd95,10'd295};
ram[7548] = {9'd98,10'd298};
ram[7549] = {-9'd99,10'd301};
ram[7550] = {-9'd96,10'd304};
ram[7551] = {-9'd93,10'd307};
ram[7552] = {-9'd93,10'd307};
ram[7553] = {-9'd90,10'd311};
ram[7554] = {-9'd87,10'd314};
ram[7555] = {-9'd84,10'd317};
ram[7556] = {-9'd81,10'd320};
ram[7557] = {-9'd77,10'd323};
ram[7558] = {-9'd74,10'd326};
ram[7559] = {-9'd71,10'd329};
ram[7560] = {-9'd68,10'd333};
ram[7561] = {-9'd65,10'd336};
ram[7562] = {-9'd62,10'd339};
ram[7563] = {-9'd59,10'd342};
ram[7564] = {-9'd55,10'd345};
ram[7565] = {-9'd52,10'd348};
ram[7566] = {-9'd49,10'd351};
ram[7567] = {-9'd46,10'd354};
ram[7568] = {-9'd43,10'd358};
ram[7569] = {-9'd40,10'd361};
ram[7570] = {-9'd37,10'd364};
ram[7571] = {-9'd33,10'd367};
ram[7572] = {-9'd30,10'd370};
ram[7573] = {-9'd27,10'd373};
ram[7574] = {-9'd24,10'd376};
ram[7575] = {-9'd21,10'd380};
ram[7576] = {-9'd18,10'd383};
ram[7577] = {-9'd15,10'd386};
ram[7578] = {-9'd11,10'd389};
ram[7579] = {-9'd8,10'd392};
ram[7580] = {-9'd5,10'd395};
ram[7581] = {-9'd2,10'd398};
ram[7582] = {9'd1,-10'd399};
ram[7583] = {9'd4,-10'd396};
ram[7584] = {9'd7,-10'd393};
ram[7585] = {9'd10,-10'd390};
ram[7586] = {9'd14,-10'd387};
ram[7587] = {9'd17,-10'd384};
ram[7588] = {9'd20,-10'd381};
ram[7589] = {9'd23,-10'd377};
ram[7590] = {9'd26,-10'd374};
ram[7591] = {9'd29,-10'd371};
ram[7592] = {9'd32,-10'd368};
ram[7593] = {9'd36,-10'd365};
ram[7594] = {9'd39,-10'd362};
ram[7595] = {9'd42,-10'd359};
ram[7596] = {9'd45,-10'd355};
ram[7597] = {9'd48,-10'd352};
ram[7598] = {9'd51,-10'd349};
ram[7599] = {9'd54,-10'd346};
ram[7600] = {9'd58,-10'd343};
ram[7601] = {9'd61,-10'd340};
ram[7602] = {9'd64,-10'd337};
ram[7603] = {9'd67,-10'd334};
ram[7604] = {9'd70,-10'd330};
ram[7605] = {9'd73,-10'd327};
ram[7606] = {9'd76,-10'd324};
ram[7607] = {9'd80,-10'd321};
ram[7608] = {9'd83,-10'd318};
ram[7609] = {9'd86,-10'd315};
ram[7610] = {9'd89,-10'd312};
ram[7611] = {9'd92,-10'd308};
ram[7612] = {9'd95,-10'd305};
ram[7613] = {9'd98,-10'd302};
ram[7614] = {-9'd99,-10'd299};
ram[7615] = {-9'd96,-10'd296};
ram[7616] = {-9'd92,-10'd293};
ram[7617] = {-9'd89,-10'd290};
ram[7618] = {-9'd86,-10'd286};
ram[7619] = {-9'd83,-10'd283};
ram[7620] = {-9'd80,-10'd280};
ram[7621] = {-9'd77,-10'd277};
ram[7622] = {-9'd74,-10'd274};
ram[7623] = {-9'd70,-10'd271};
ram[7624] = {-9'd67,-10'd268};
ram[7625] = {-9'd64,-10'd264};
ram[7626] = {-9'd61,-10'd261};
ram[7627] = {-9'd58,-10'd258};
ram[7628] = {-9'd55,-10'd255};
ram[7629] = {-9'd52,-10'd252};
ram[7630] = {-9'd48,-10'd249};
ram[7631] = {-9'd45,-10'd246};
ram[7632] = {-9'd42,-10'd242};
ram[7633] = {-9'd39,-10'd239};
ram[7634] = {-9'd36,-10'd236};
ram[7635] = {-9'd33,-10'd233};
ram[7636] = {-9'd30,-10'd230};
ram[7637] = {-9'd26,-10'd227};
ram[7638] = {-9'd23,-10'd224};
ram[7639] = {-9'd20,-10'd220};
ram[7640] = {-9'd17,-10'd217};
ram[7641] = {-9'd14,-10'd214};
ram[7642] = {-9'd11,-10'd211};
ram[7643] = {-9'd8,-10'd208};
ram[7644] = {-9'd4,-10'd205};
ram[7645] = {-9'd1,-10'd202};
ram[7646] = {9'd2,-10'd198};
ram[7647] = {9'd5,-10'd195};
ram[7648] = {9'd8,-10'd192};
ram[7649] = {9'd11,-10'd189};
ram[7650] = {9'd14,-10'd186};
ram[7651] = {9'd18,-10'd183};
ram[7652] = {9'd21,-10'd180};
ram[7653] = {9'd24,-10'd176};
ram[7654] = {9'd27,-10'd173};
ram[7655] = {9'd30,-10'd170};
ram[7656] = {9'd33,-10'd167};
ram[7657] = {9'd36,-10'd164};
ram[7658] = {9'd40,-10'd161};
ram[7659] = {9'd43,-10'd158};
ram[7660] = {9'd46,-10'd154};
ram[7661] = {9'd49,-10'd151};
ram[7662] = {9'd52,-10'd148};
ram[7663] = {9'd55,-10'd145};
ram[7664] = {9'd58,-10'd142};
ram[7665] = {9'd62,-10'd139};
ram[7666] = {9'd65,-10'd136};
ram[7667] = {9'd68,-10'd132};
ram[7668] = {9'd71,-10'd129};
ram[7669] = {9'd74,-10'd126};
ram[7670] = {9'd77,-10'd123};
ram[7671] = {9'd80,-10'd120};
ram[7672] = {9'd84,-10'd117};
ram[7673] = {9'd87,-10'd114};
ram[7674] = {9'd90,-10'd110};
ram[7675] = {9'd93,-10'd107};
ram[7676] = {9'd96,-10'd104};
ram[7677] = {9'd99,-10'd101};
ram[7678] = {-9'd98,-10'd98};
ram[7679] = {-9'd95,-10'd95};
ram[7680] = {-9'd95,-10'd95};
ram[7681] = {-9'd92,-10'd92};
ram[7682] = {-9'd88,-10'd88};
ram[7683] = {-9'd85,-10'd85};
ram[7684] = {-9'd82,-10'd82};
ram[7685] = {-9'd79,-10'd79};
ram[7686] = {-9'd76,-10'd76};
ram[7687] = {-9'd73,-10'd73};
ram[7688] = {-9'd70,-10'd70};
ram[7689] = {-9'd66,-10'd66};
ram[7690] = {-9'd63,-10'd63};
ram[7691] = {-9'd60,-10'd60};
ram[7692] = {-9'd57,-10'd57};
ram[7693] = {-9'd54,-10'd54};
ram[7694] = {-9'd51,-10'd51};
ram[7695] = {-9'd48,-10'd48};
ram[7696] = {-9'd44,-10'd44};
ram[7697] = {-9'd41,-10'd41};
ram[7698] = {-9'd38,-10'd38};
ram[7699] = {-9'd35,-10'd35};
ram[7700] = {-9'd32,-10'd32};
ram[7701] = {-9'd29,-10'd29};
ram[7702] = {-9'd26,-10'd26};
ram[7703] = {-9'd22,-10'd22};
ram[7704] = {-9'd19,-10'd19};
ram[7705] = {-9'd16,-10'd16};
ram[7706] = {-9'd13,-10'd13};
ram[7707] = {-9'd10,-10'd10};
ram[7708] = {-9'd7,-10'd7};
ram[7709] = {-9'd4,-10'd4};
ram[7710] = {9'd0,10'd0};
ram[7711] = {9'd3,10'd3};
ram[7712] = {9'd6,10'd6};
ram[7713] = {9'd9,10'd9};
ram[7714] = {9'd12,10'd12};
ram[7715] = {9'd15,10'd15};
ram[7716] = {9'd18,10'd18};
ram[7717] = {9'd21,10'd21};
ram[7718] = {9'd25,10'd25};
ram[7719] = {9'd28,10'd28};
ram[7720] = {9'd31,10'd31};
ram[7721] = {9'd34,10'd34};
ram[7722] = {9'd37,10'd37};
ram[7723] = {9'd40,10'd40};
ram[7724] = {9'd43,10'd43};
ram[7725] = {9'd47,10'd47};
ram[7726] = {9'd50,10'd50};
ram[7727] = {9'd53,10'd53};
ram[7728] = {9'd56,10'd56};
ram[7729] = {9'd59,10'd59};
ram[7730] = {9'd62,10'd62};
ram[7731] = {9'd65,10'd65};
ram[7732] = {9'd69,10'd69};
ram[7733] = {9'd72,10'd72};
ram[7734] = {9'd75,10'd75};
ram[7735] = {9'd78,10'd78};
ram[7736] = {9'd81,10'd81};
ram[7737] = {9'd84,10'd84};
ram[7738] = {9'd87,10'd87};
ram[7739] = {9'd91,10'd91};
ram[7740] = {9'd94,10'd94};
ram[7741] = {9'd97,10'd97};
ram[7742] = {-9'd100,10'd100};
ram[7743] = {-9'd97,10'd103};
ram[7744] = {-9'd94,10'd106};
ram[7745] = {-9'd91,10'd109};
ram[7746] = {-9'd88,10'd113};
ram[7747] = {-9'd85,10'd116};
ram[7748] = {-9'd81,10'd119};
ram[7749] = {-9'd78,10'd122};
ram[7750] = {-9'd75,10'd125};
ram[7751] = {-9'd72,10'd128};
ram[7752] = {-9'd69,10'd131};
ram[7753] = {-9'd66,10'd135};
ram[7754] = {-9'd63,10'd138};
ram[7755] = {-9'd59,10'd141};
ram[7756] = {-9'd56,10'd144};
ram[7757] = {-9'd53,10'd147};
ram[7758] = {-9'd50,10'd150};
ram[7759] = {-9'd47,10'd153};
ram[7760] = {-9'd44,10'd157};
ram[7761] = {-9'd41,10'd160};
ram[7762] = {-9'd37,10'd163};
ram[7763] = {-9'd34,10'd166};
ram[7764] = {-9'd31,10'd169};
ram[7765] = {-9'd28,10'd172};
ram[7766] = {-9'd25,10'd175};
ram[7767] = {-9'd22,10'd179};
ram[7768] = {-9'd19,10'd182};
ram[7769] = {-9'd15,10'd185};
ram[7770] = {-9'd12,10'd188};
ram[7771] = {-9'd9,10'd191};
ram[7772] = {-9'd6,10'd194};
ram[7773] = {-9'd3,10'd197};
ram[7774] = {9'd0,10'd201};
ram[7775] = {9'd3,10'd204};
ram[7776] = {9'd7,10'd207};
ram[7777] = {9'd10,10'd210};
ram[7778] = {9'd13,10'd213};
ram[7779] = {9'd16,10'd216};
ram[7780] = {9'd19,10'd219};
ram[7781] = {9'd22,10'd223};
ram[7782] = {9'd25,10'd226};
ram[7783] = {9'd29,10'd229};
ram[7784] = {9'd32,10'd232};
ram[7785] = {9'd35,10'd235};
ram[7786] = {9'd38,10'd238};
ram[7787] = {9'd41,10'd241};
ram[7788] = {9'd44,10'd245};
ram[7789] = {9'd47,10'd248};
ram[7790] = {9'd51,10'd251};
ram[7791] = {9'd54,10'd254};
ram[7792] = {9'd57,10'd257};
ram[7793] = {9'd60,10'd260};
ram[7794] = {9'd63,10'd263};
ram[7795] = {9'd66,10'd267};
ram[7796] = {9'd69,10'd270};
ram[7797] = {9'd73,10'd273};
ram[7798] = {9'd76,10'd276};
ram[7799] = {9'd79,10'd279};
ram[7800] = {9'd82,10'd282};
ram[7801] = {9'd85,10'd285};
ram[7802] = {9'd88,10'd289};
ram[7803] = {9'd91,10'd292};
ram[7804] = {9'd95,10'd295};
ram[7805] = {9'd98,10'd298};
ram[7806] = {-9'd99,10'd301};
ram[7807] = {-9'd96,10'd304};
ram[7808] = {-9'd96,10'd304};
ram[7809] = {-9'd93,10'd307};
ram[7810] = {-9'd90,10'd311};
ram[7811] = {-9'd87,10'd314};
ram[7812] = {-9'd84,10'd317};
ram[7813] = {-9'd81,10'd320};
ram[7814] = {-9'd77,10'd323};
ram[7815] = {-9'd74,10'd326};
ram[7816] = {-9'd71,10'd329};
ram[7817] = {-9'd68,10'd333};
ram[7818] = {-9'd65,10'd336};
ram[7819] = {-9'd62,10'd339};
ram[7820] = {-9'd59,10'd342};
ram[7821] = {-9'd55,10'd345};
ram[7822] = {-9'd52,10'd348};
ram[7823] = {-9'd49,10'd351};
ram[7824] = {-9'd46,10'd354};
ram[7825] = {-9'd43,10'd358};
ram[7826] = {-9'd40,10'd361};
ram[7827] = {-9'd37,10'd364};
ram[7828] = {-9'd33,10'd367};
ram[7829] = {-9'd30,10'd370};
ram[7830] = {-9'd27,10'd373};
ram[7831] = {-9'd24,10'd376};
ram[7832] = {-9'd21,10'd380};
ram[7833] = {-9'd18,10'd383};
ram[7834] = {-9'd15,10'd386};
ram[7835] = {-9'd11,10'd389};
ram[7836] = {-9'd8,10'd392};
ram[7837] = {-9'd5,10'd395};
ram[7838] = {-9'd2,10'd398};
ram[7839] = {9'd1,-10'd399};
ram[7840] = {9'd4,-10'd396};
ram[7841] = {9'd7,-10'd393};
ram[7842] = {9'd10,-10'd390};
ram[7843] = {9'd14,-10'd387};
ram[7844] = {9'd17,-10'd384};
ram[7845] = {9'd20,-10'd381};
ram[7846] = {9'd23,-10'd377};
ram[7847] = {9'd26,-10'd374};
ram[7848] = {9'd29,-10'd371};
ram[7849] = {9'd32,-10'd368};
ram[7850] = {9'd36,-10'd365};
ram[7851] = {9'd39,-10'd362};
ram[7852] = {9'd42,-10'd359};
ram[7853] = {9'd45,-10'd355};
ram[7854] = {9'd48,-10'd352};
ram[7855] = {9'd51,-10'd349};
ram[7856] = {9'd54,-10'd346};
ram[7857] = {9'd58,-10'd343};
ram[7858] = {9'd61,-10'd340};
ram[7859] = {9'd64,-10'd337};
ram[7860] = {9'd67,-10'd334};
ram[7861] = {9'd70,-10'd330};
ram[7862] = {9'd73,-10'd327};
ram[7863] = {9'd76,-10'd324};
ram[7864] = {9'd80,-10'd321};
ram[7865] = {9'd83,-10'd318};
ram[7866] = {9'd86,-10'd315};
ram[7867] = {9'd89,-10'd312};
ram[7868] = {9'd92,-10'd308};
ram[7869] = {9'd95,-10'd305};
ram[7870] = {9'd98,-10'd302};
ram[7871] = {-9'd99,-10'd299};
ram[7872] = {-9'd96,-10'd296};
ram[7873] = {-9'd92,-10'd293};
ram[7874] = {-9'd89,-10'd290};
ram[7875] = {-9'd86,-10'd286};
ram[7876] = {-9'd83,-10'd283};
ram[7877] = {-9'd80,-10'd280};
ram[7878] = {-9'd77,-10'd277};
ram[7879] = {-9'd74,-10'd274};
ram[7880] = {-9'd70,-10'd271};
ram[7881] = {-9'd67,-10'd268};
ram[7882] = {-9'd64,-10'd264};
ram[7883] = {-9'd61,-10'd261};
ram[7884] = {-9'd58,-10'd258};
ram[7885] = {-9'd55,-10'd255};
ram[7886] = {-9'd52,-10'd252};
ram[7887] = {-9'd48,-10'd249};
ram[7888] = {-9'd45,-10'd246};
ram[7889] = {-9'd42,-10'd242};
ram[7890] = {-9'd39,-10'd239};
ram[7891] = {-9'd36,-10'd236};
ram[7892] = {-9'd33,-10'd233};
ram[7893] = {-9'd30,-10'd230};
ram[7894] = {-9'd26,-10'd227};
ram[7895] = {-9'd23,-10'd224};
ram[7896] = {-9'd20,-10'd220};
ram[7897] = {-9'd17,-10'd217};
ram[7898] = {-9'd14,-10'd214};
ram[7899] = {-9'd11,-10'd211};
ram[7900] = {-9'd8,-10'd208};
ram[7901] = {-9'd4,-10'd205};
ram[7902] = {-9'd1,-10'd202};
ram[7903] = {9'd2,-10'd198};
ram[7904] = {9'd5,-10'd195};
ram[7905] = {9'd8,-10'd192};
ram[7906] = {9'd11,-10'd189};
ram[7907] = {9'd14,-10'd186};
ram[7908] = {9'd18,-10'd183};
ram[7909] = {9'd21,-10'd180};
ram[7910] = {9'd24,-10'd176};
ram[7911] = {9'd27,-10'd173};
ram[7912] = {9'd30,-10'd170};
ram[7913] = {9'd33,-10'd167};
ram[7914] = {9'd36,-10'd164};
ram[7915] = {9'd40,-10'd161};
ram[7916] = {9'd43,-10'd158};
ram[7917] = {9'd46,-10'd154};
ram[7918] = {9'd49,-10'd151};
ram[7919] = {9'd52,-10'd148};
ram[7920] = {9'd55,-10'd145};
ram[7921] = {9'd58,-10'd142};
ram[7922] = {9'd62,-10'd139};
ram[7923] = {9'd65,-10'd136};
ram[7924] = {9'd68,-10'd132};
ram[7925] = {9'd71,-10'd129};
ram[7926] = {9'd74,-10'd126};
ram[7927] = {9'd77,-10'd123};
ram[7928] = {9'd80,-10'd120};
ram[7929] = {9'd84,-10'd117};
ram[7930] = {9'd87,-10'd114};
ram[7931] = {9'd90,-10'd110};
ram[7932] = {9'd93,-10'd107};
ram[7933] = {9'd96,-10'd104};
ram[7934] = {9'd99,-10'd101};
ram[7935] = {-9'd98,-10'd98};
ram[7936] = {-9'd98,-10'd98};
ram[7937] = {-9'd95,-10'd95};
ram[7938] = {-9'd92,-10'd92};
ram[7939] = {-9'd88,-10'd88};
ram[7940] = {-9'd85,-10'd85};
ram[7941] = {-9'd82,-10'd82};
ram[7942] = {-9'd79,-10'd79};
ram[7943] = {-9'd76,-10'd76};
ram[7944] = {-9'd73,-10'd73};
ram[7945] = {-9'd70,-10'd70};
ram[7946] = {-9'd66,-10'd66};
ram[7947] = {-9'd63,-10'd63};
ram[7948] = {-9'd60,-10'd60};
ram[7949] = {-9'd57,-10'd57};
ram[7950] = {-9'd54,-10'd54};
ram[7951] = {-9'd51,-10'd51};
ram[7952] = {-9'd48,-10'd48};
ram[7953] = {-9'd44,-10'd44};
ram[7954] = {-9'd41,-10'd41};
ram[7955] = {-9'd38,-10'd38};
ram[7956] = {-9'd35,-10'd35};
ram[7957] = {-9'd32,-10'd32};
ram[7958] = {-9'd29,-10'd29};
ram[7959] = {-9'd26,-10'd26};
ram[7960] = {-9'd22,-10'd22};
ram[7961] = {-9'd19,-10'd19};
ram[7962] = {-9'd16,-10'd16};
ram[7963] = {-9'd13,-10'd13};
ram[7964] = {-9'd10,-10'd10};
ram[7965] = {-9'd7,-10'd7};
ram[7966] = {-9'd4,-10'd4};
ram[7967] = {9'd0,10'd0};
ram[7968] = {9'd3,10'd3};
ram[7969] = {9'd6,10'd6};
ram[7970] = {9'd9,10'd9};
ram[7971] = {9'd12,10'd12};
ram[7972] = {9'd15,10'd15};
ram[7973] = {9'd18,10'd18};
ram[7974] = {9'd21,10'd21};
ram[7975] = {9'd25,10'd25};
ram[7976] = {9'd28,10'd28};
ram[7977] = {9'd31,10'd31};
ram[7978] = {9'd34,10'd34};
ram[7979] = {9'd37,10'd37};
ram[7980] = {9'd40,10'd40};
ram[7981] = {9'd43,10'd43};
ram[7982] = {9'd47,10'd47};
ram[7983] = {9'd50,10'd50};
ram[7984] = {9'd53,10'd53};
ram[7985] = {9'd56,10'd56};
ram[7986] = {9'd59,10'd59};
ram[7987] = {9'd62,10'd62};
ram[7988] = {9'd65,10'd65};
ram[7989] = {9'd69,10'd69};
ram[7990] = {9'd72,10'd72};
ram[7991] = {9'd75,10'd75};
ram[7992] = {9'd78,10'd78};
ram[7993] = {9'd81,10'd81};
ram[7994] = {9'd84,10'd84};
ram[7995] = {9'd87,10'd87};
ram[7996] = {9'd91,10'd91};
ram[7997] = {9'd94,10'd94};
ram[7998] = {9'd97,10'd97};
ram[7999] = {-9'd100,10'd100};
ram[8000] = {-9'd97,10'd103};
ram[8001] = {-9'd94,10'd106};
ram[8002] = {-9'd91,10'd109};
ram[8003] = {-9'd88,10'd113};
ram[8004] = {-9'd85,10'd116};
ram[8005] = {-9'd81,10'd119};
ram[8006] = {-9'd78,10'd122};
ram[8007] = {-9'd75,10'd125};
ram[8008] = {-9'd72,10'd128};
ram[8009] = {-9'd69,10'd131};
ram[8010] = {-9'd66,10'd135};
ram[8011] = {-9'd63,10'd138};
ram[8012] = {-9'd59,10'd141};
ram[8013] = {-9'd56,10'd144};
ram[8014] = {-9'd53,10'd147};
ram[8015] = {-9'd50,10'd150};
ram[8016] = {-9'd47,10'd153};
ram[8017] = {-9'd44,10'd157};
ram[8018] = {-9'd41,10'd160};
ram[8019] = {-9'd37,10'd163};
ram[8020] = {-9'd34,10'd166};
ram[8021] = {-9'd31,10'd169};
ram[8022] = {-9'd28,10'd172};
ram[8023] = {-9'd25,10'd175};
ram[8024] = {-9'd22,10'd179};
ram[8025] = {-9'd19,10'd182};
ram[8026] = {-9'd15,10'd185};
ram[8027] = {-9'd12,10'd188};
ram[8028] = {-9'd9,10'd191};
ram[8029] = {-9'd6,10'd194};
ram[8030] = {-9'd3,10'd197};
ram[8031] = {9'd0,10'd201};
ram[8032] = {9'd3,10'd204};
ram[8033] = {9'd7,10'd207};
ram[8034] = {9'd10,10'd210};
ram[8035] = {9'd13,10'd213};
ram[8036] = {9'd16,10'd216};
ram[8037] = {9'd19,10'd219};
ram[8038] = {9'd22,10'd223};
ram[8039] = {9'd25,10'd226};
ram[8040] = {9'd29,10'd229};
ram[8041] = {9'd32,10'd232};
ram[8042] = {9'd35,10'd235};
ram[8043] = {9'd38,10'd238};
ram[8044] = {9'd41,10'd241};
ram[8045] = {9'd44,10'd245};
ram[8046] = {9'd47,10'd248};
ram[8047] = {9'd51,10'd251};
ram[8048] = {9'd54,10'd254};
ram[8049] = {9'd57,10'd257};
ram[8050] = {9'd60,10'd260};
ram[8051] = {9'd63,10'd263};
ram[8052] = {9'd66,10'd267};
ram[8053] = {9'd69,10'd270};
ram[8054] = {9'd73,10'd273};
ram[8055] = {9'd76,10'd276};
ram[8056] = {9'd79,10'd279};
ram[8057] = {9'd82,10'd282};
ram[8058] = {9'd85,10'd285};
ram[8059] = {9'd88,10'd289};
ram[8060] = {9'd91,10'd292};
ram[8061] = {9'd95,10'd295};
ram[8062] = {9'd98,10'd298};
ram[8063] = {-9'd99,10'd301};
ram[8064] = {-9'd99,10'd301};
ram[8065] = {-9'd96,10'd304};
ram[8066] = {-9'd93,10'd307};
ram[8067] = {-9'd90,10'd311};
ram[8068] = {-9'd87,10'd314};
ram[8069] = {-9'd84,10'd317};
ram[8070] = {-9'd81,10'd320};
ram[8071] = {-9'd77,10'd323};
ram[8072] = {-9'd74,10'd326};
ram[8073] = {-9'd71,10'd329};
ram[8074] = {-9'd68,10'd333};
ram[8075] = {-9'd65,10'd336};
ram[8076] = {-9'd62,10'd339};
ram[8077] = {-9'd59,10'd342};
ram[8078] = {-9'd55,10'd345};
ram[8079] = {-9'd52,10'd348};
ram[8080] = {-9'd49,10'd351};
ram[8081] = {-9'd46,10'd354};
ram[8082] = {-9'd43,10'd358};
ram[8083] = {-9'd40,10'd361};
ram[8084] = {-9'd37,10'd364};
ram[8085] = {-9'd33,10'd367};
ram[8086] = {-9'd30,10'd370};
ram[8087] = {-9'd27,10'd373};
ram[8088] = {-9'd24,10'd376};
ram[8089] = {-9'd21,10'd380};
ram[8090] = {-9'd18,10'd383};
ram[8091] = {-9'd15,10'd386};
ram[8092] = {-9'd11,10'd389};
ram[8093] = {-9'd8,10'd392};
ram[8094] = {-9'd5,10'd395};
ram[8095] = {-9'd2,10'd398};
ram[8096] = {9'd1,-10'd399};
ram[8097] = {9'd4,-10'd396};
ram[8098] = {9'd7,-10'd393};
ram[8099] = {9'd10,-10'd390};
ram[8100] = {9'd14,-10'd387};
ram[8101] = {9'd17,-10'd384};
ram[8102] = {9'd20,-10'd381};
ram[8103] = {9'd23,-10'd377};
ram[8104] = {9'd26,-10'd374};
ram[8105] = {9'd29,-10'd371};
ram[8106] = {9'd32,-10'd368};
ram[8107] = {9'd36,-10'd365};
ram[8108] = {9'd39,-10'd362};
ram[8109] = {9'd42,-10'd359};
ram[8110] = {9'd45,-10'd355};
ram[8111] = {9'd48,-10'd352};
ram[8112] = {9'd51,-10'd349};
ram[8113] = {9'd54,-10'd346};
ram[8114] = {9'd58,-10'd343};
ram[8115] = {9'd61,-10'd340};
ram[8116] = {9'd64,-10'd337};
ram[8117] = {9'd67,-10'd334};
ram[8118] = {9'd70,-10'd330};
ram[8119] = {9'd73,-10'd327};
ram[8120] = {9'd76,-10'd324};
ram[8121] = {9'd80,-10'd321};
ram[8122] = {9'd83,-10'd318};
ram[8123] = {9'd86,-10'd315};
ram[8124] = {9'd89,-10'd312};
ram[8125] = {9'd92,-10'd308};
ram[8126] = {9'd95,-10'd305};
ram[8127] = {9'd98,-10'd302};
ram[8128] = {-9'd99,-10'd299};
ram[8129] = {-9'd96,-10'd296};
ram[8130] = {-9'd92,-10'd293};
ram[8131] = {-9'd89,-10'd290};
ram[8132] = {-9'd86,-10'd286};
ram[8133] = {-9'd83,-10'd283};
ram[8134] = {-9'd80,-10'd280};
ram[8135] = {-9'd77,-10'd277};
ram[8136] = {-9'd74,-10'd274};
ram[8137] = {-9'd70,-10'd271};
ram[8138] = {-9'd67,-10'd268};
ram[8139] = {-9'd64,-10'd264};
ram[8140] = {-9'd61,-10'd261};
ram[8141] = {-9'd58,-10'd258};
ram[8142] = {-9'd55,-10'd255};
ram[8143] = {-9'd52,-10'd252};
ram[8144] = {-9'd48,-10'd249};
ram[8145] = {-9'd45,-10'd246};
ram[8146] = {-9'd42,-10'd242};
ram[8147] = {-9'd39,-10'd239};
ram[8148] = {-9'd36,-10'd236};
ram[8149] = {-9'd33,-10'd233};
ram[8150] = {-9'd30,-10'd230};
ram[8151] = {-9'd26,-10'd227};
ram[8152] = {-9'd23,-10'd224};
ram[8153] = {-9'd20,-10'd220};
ram[8154] = {-9'd17,-10'd217};
ram[8155] = {-9'd14,-10'd214};
ram[8156] = {-9'd11,-10'd211};
ram[8157] = {-9'd8,-10'd208};
ram[8158] = {-9'd4,-10'd205};
ram[8159] = {-9'd1,-10'd202};
ram[8160] = {9'd2,-10'd198};
ram[8161] = {9'd5,-10'd195};
ram[8162] = {9'd8,-10'd192};
ram[8163] = {9'd11,-10'd189};
ram[8164] = {9'd14,-10'd186};
ram[8165] = {9'd18,-10'd183};
ram[8166] = {9'd21,-10'd180};
ram[8167] = {9'd24,-10'd176};
ram[8168] = {9'd27,-10'd173};
ram[8169] = {9'd30,-10'd170};
ram[8170] = {9'd33,-10'd167};
ram[8171] = {9'd36,-10'd164};
ram[8172] = {9'd40,-10'd161};
ram[8173] = {9'd43,-10'd158};
ram[8174] = {9'd46,-10'd154};
ram[8175] = {9'd49,-10'd151};
ram[8176] = {9'd52,-10'd148};
ram[8177] = {9'd55,-10'd145};
ram[8178] = {9'd58,-10'd142};
ram[8179] = {9'd62,-10'd139};
ram[8180] = {9'd65,-10'd136};
ram[8181] = {9'd68,-10'd132};
ram[8182] = {9'd71,-10'd129};
ram[8183] = {9'd74,-10'd126};
ram[8184] = {9'd77,-10'd123};
ram[8185] = {9'd80,-10'd120};
ram[8186] = {9'd84,-10'd117};
ram[8187] = {9'd87,-10'd114};
ram[8188] = {9'd90,-10'd110};
ram[8189] = {9'd93,-10'd107};
ram[8190] = {9'd96,-10'd104};
ram[8191] = {9'd99,-10'd101};
ram[8192] = {9'd99,-10'd101};
ram[8193] = {-9'd98,-10'd98};
ram[8194] = {-9'd95,-10'd95};
ram[8195] = {-9'd92,-10'd92};
ram[8196] = {-9'd88,-10'd88};
ram[8197] = {-9'd85,-10'd85};
ram[8198] = {-9'd82,-10'd82};
ram[8199] = {-9'd79,-10'd79};
ram[8200] = {-9'd76,-10'd76};
ram[8201] = {-9'd73,-10'd73};
ram[8202] = {-9'd70,-10'd70};
ram[8203] = {-9'd66,-10'd66};
ram[8204] = {-9'd63,-10'd63};
ram[8205] = {-9'd60,-10'd60};
ram[8206] = {-9'd57,-10'd57};
ram[8207] = {-9'd54,-10'd54};
ram[8208] = {-9'd51,-10'd51};
ram[8209] = {-9'd48,-10'd48};
ram[8210] = {-9'd44,-10'd44};
ram[8211] = {-9'd41,-10'd41};
ram[8212] = {-9'd38,-10'd38};
ram[8213] = {-9'd35,-10'd35};
ram[8214] = {-9'd32,-10'd32};
ram[8215] = {-9'd29,-10'd29};
ram[8216] = {-9'd26,-10'd26};
ram[8217] = {-9'd22,-10'd22};
ram[8218] = {-9'd19,-10'd19};
ram[8219] = {-9'd16,-10'd16};
ram[8220] = {-9'd13,-10'd13};
ram[8221] = {-9'd10,-10'd10};
ram[8222] = {-9'd7,-10'd7};
ram[8223] = {-9'd4,-10'd4};
ram[8224] = {9'd0,10'd0};
ram[8225] = {9'd3,10'd3};
ram[8226] = {9'd6,10'd6};
ram[8227] = {9'd9,10'd9};
ram[8228] = {9'd12,10'd12};
ram[8229] = {9'd15,10'd15};
ram[8230] = {9'd18,10'd18};
ram[8231] = {9'd21,10'd21};
ram[8232] = {9'd25,10'd25};
ram[8233] = {9'd28,10'd28};
ram[8234] = {9'd31,10'd31};
ram[8235] = {9'd34,10'd34};
ram[8236] = {9'd37,10'd37};
ram[8237] = {9'd40,10'd40};
ram[8238] = {9'd43,10'd43};
ram[8239] = {9'd47,10'd47};
ram[8240] = {9'd50,10'd50};
ram[8241] = {9'd53,10'd53};
ram[8242] = {9'd56,10'd56};
ram[8243] = {9'd59,10'd59};
ram[8244] = {9'd62,10'd62};
ram[8245] = {9'd65,10'd65};
ram[8246] = {9'd69,10'd69};
ram[8247] = {9'd72,10'd72};
ram[8248] = {9'd75,10'd75};
ram[8249] = {9'd78,10'd78};
ram[8250] = {9'd81,10'd81};
ram[8251] = {9'd84,10'd84};
ram[8252] = {9'd87,10'd87};
ram[8253] = {9'd91,10'd91};
ram[8254] = {9'd94,10'd94};
ram[8255] = {9'd97,10'd97};
ram[8256] = {-9'd100,10'd100};
ram[8257] = {-9'd97,10'd103};
ram[8258] = {-9'd94,10'd106};
ram[8259] = {-9'd91,10'd109};
ram[8260] = {-9'd88,10'd113};
ram[8261] = {-9'd85,10'd116};
ram[8262] = {-9'd81,10'd119};
ram[8263] = {-9'd78,10'd122};
ram[8264] = {-9'd75,10'd125};
ram[8265] = {-9'd72,10'd128};
ram[8266] = {-9'd69,10'd131};
ram[8267] = {-9'd66,10'd135};
ram[8268] = {-9'd63,10'd138};
ram[8269] = {-9'd59,10'd141};
ram[8270] = {-9'd56,10'd144};
ram[8271] = {-9'd53,10'd147};
ram[8272] = {-9'd50,10'd150};
ram[8273] = {-9'd47,10'd153};
ram[8274] = {-9'd44,10'd157};
ram[8275] = {-9'd41,10'd160};
ram[8276] = {-9'd37,10'd163};
ram[8277] = {-9'd34,10'd166};
ram[8278] = {-9'd31,10'd169};
ram[8279] = {-9'd28,10'd172};
ram[8280] = {-9'd25,10'd175};
ram[8281] = {-9'd22,10'd179};
ram[8282] = {-9'd19,10'd182};
ram[8283] = {-9'd15,10'd185};
ram[8284] = {-9'd12,10'd188};
ram[8285] = {-9'd9,10'd191};
ram[8286] = {-9'd6,10'd194};
ram[8287] = {-9'd3,10'd197};
ram[8288] = {9'd0,10'd201};
ram[8289] = {9'd3,10'd204};
ram[8290] = {9'd7,10'd207};
ram[8291] = {9'd10,10'd210};
ram[8292] = {9'd13,10'd213};
ram[8293] = {9'd16,10'd216};
ram[8294] = {9'd19,10'd219};
ram[8295] = {9'd22,10'd223};
ram[8296] = {9'd25,10'd226};
ram[8297] = {9'd29,10'd229};
ram[8298] = {9'd32,10'd232};
ram[8299] = {9'd35,10'd235};
ram[8300] = {9'd38,10'd238};
ram[8301] = {9'd41,10'd241};
ram[8302] = {9'd44,10'd245};
ram[8303] = {9'd47,10'd248};
ram[8304] = {9'd51,10'd251};
ram[8305] = {9'd54,10'd254};
ram[8306] = {9'd57,10'd257};
ram[8307] = {9'd60,10'd260};
ram[8308] = {9'd63,10'd263};
ram[8309] = {9'd66,10'd267};
ram[8310] = {9'd69,10'd270};
ram[8311] = {9'd73,10'd273};
ram[8312] = {9'd76,10'd276};
ram[8313] = {9'd79,10'd279};
ram[8314] = {9'd82,10'd282};
ram[8315] = {9'd85,10'd285};
ram[8316] = {9'd88,10'd289};
ram[8317] = {9'd91,10'd292};
ram[8318] = {9'd95,10'd295};
ram[8319] = {9'd98,10'd298};
ram[8320] = {9'd98,10'd298};
ram[8321] = {-9'd99,10'd301};
ram[8322] = {-9'd96,10'd304};
ram[8323] = {-9'd93,10'd307};
ram[8324] = {-9'd90,10'd311};
ram[8325] = {-9'd87,10'd314};
ram[8326] = {-9'd84,10'd317};
ram[8327] = {-9'd81,10'd320};
ram[8328] = {-9'd77,10'd323};
ram[8329] = {-9'd74,10'd326};
ram[8330] = {-9'd71,10'd329};
ram[8331] = {-9'd68,10'd333};
ram[8332] = {-9'd65,10'd336};
ram[8333] = {-9'd62,10'd339};
ram[8334] = {-9'd59,10'd342};
ram[8335] = {-9'd55,10'd345};
ram[8336] = {-9'd52,10'd348};
ram[8337] = {-9'd49,10'd351};
ram[8338] = {-9'd46,10'd354};
ram[8339] = {-9'd43,10'd358};
ram[8340] = {-9'd40,10'd361};
ram[8341] = {-9'd37,10'd364};
ram[8342] = {-9'd33,10'd367};
ram[8343] = {-9'd30,10'd370};
ram[8344] = {-9'd27,10'd373};
ram[8345] = {-9'd24,10'd376};
ram[8346] = {-9'd21,10'd380};
ram[8347] = {-9'd18,10'd383};
ram[8348] = {-9'd15,10'd386};
ram[8349] = {-9'd11,10'd389};
ram[8350] = {-9'd8,10'd392};
ram[8351] = {-9'd5,10'd395};
ram[8352] = {-9'd2,10'd398};
ram[8353] = {9'd1,-10'd399};
ram[8354] = {9'd4,-10'd396};
ram[8355] = {9'd7,-10'd393};
ram[8356] = {9'd10,-10'd390};
ram[8357] = {9'd14,-10'd387};
ram[8358] = {9'd17,-10'd384};
ram[8359] = {9'd20,-10'd381};
ram[8360] = {9'd23,-10'd377};
ram[8361] = {9'd26,-10'd374};
ram[8362] = {9'd29,-10'd371};
ram[8363] = {9'd32,-10'd368};
ram[8364] = {9'd36,-10'd365};
ram[8365] = {9'd39,-10'd362};
ram[8366] = {9'd42,-10'd359};
ram[8367] = {9'd45,-10'd355};
ram[8368] = {9'd48,-10'd352};
ram[8369] = {9'd51,-10'd349};
ram[8370] = {9'd54,-10'd346};
ram[8371] = {9'd58,-10'd343};
ram[8372] = {9'd61,-10'd340};
ram[8373] = {9'd64,-10'd337};
ram[8374] = {9'd67,-10'd334};
ram[8375] = {9'd70,-10'd330};
ram[8376] = {9'd73,-10'd327};
ram[8377] = {9'd76,-10'd324};
ram[8378] = {9'd80,-10'd321};
ram[8379] = {9'd83,-10'd318};
ram[8380] = {9'd86,-10'd315};
ram[8381] = {9'd89,-10'd312};
ram[8382] = {9'd92,-10'd308};
ram[8383] = {9'd95,-10'd305};
ram[8384] = {9'd98,-10'd302};
ram[8385] = {-9'd99,-10'd299};
ram[8386] = {-9'd96,-10'd296};
ram[8387] = {-9'd92,-10'd293};
ram[8388] = {-9'd89,-10'd290};
ram[8389] = {-9'd86,-10'd286};
ram[8390] = {-9'd83,-10'd283};
ram[8391] = {-9'd80,-10'd280};
ram[8392] = {-9'd77,-10'd277};
ram[8393] = {-9'd74,-10'd274};
ram[8394] = {-9'd70,-10'd271};
ram[8395] = {-9'd67,-10'd268};
ram[8396] = {-9'd64,-10'd264};
ram[8397] = {-9'd61,-10'd261};
ram[8398] = {-9'd58,-10'd258};
ram[8399] = {-9'd55,-10'd255};
ram[8400] = {-9'd52,-10'd252};
ram[8401] = {-9'd48,-10'd249};
ram[8402] = {-9'd45,-10'd246};
ram[8403] = {-9'd42,-10'd242};
ram[8404] = {-9'd39,-10'd239};
ram[8405] = {-9'd36,-10'd236};
ram[8406] = {-9'd33,-10'd233};
ram[8407] = {-9'd30,-10'd230};
ram[8408] = {-9'd26,-10'd227};
ram[8409] = {-9'd23,-10'd224};
ram[8410] = {-9'd20,-10'd220};
ram[8411] = {-9'd17,-10'd217};
ram[8412] = {-9'd14,-10'd214};
ram[8413] = {-9'd11,-10'd211};
ram[8414] = {-9'd8,-10'd208};
ram[8415] = {-9'd4,-10'd205};
ram[8416] = {-9'd1,-10'd202};
ram[8417] = {9'd2,-10'd198};
ram[8418] = {9'd5,-10'd195};
ram[8419] = {9'd8,-10'd192};
ram[8420] = {9'd11,-10'd189};
ram[8421] = {9'd14,-10'd186};
ram[8422] = {9'd18,-10'd183};
ram[8423] = {9'd21,-10'd180};
ram[8424] = {9'd24,-10'd176};
ram[8425] = {9'd27,-10'd173};
ram[8426] = {9'd30,-10'd170};
ram[8427] = {9'd33,-10'd167};
ram[8428] = {9'd36,-10'd164};
ram[8429] = {9'd40,-10'd161};
ram[8430] = {9'd43,-10'd158};
ram[8431] = {9'd46,-10'd154};
ram[8432] = {9'd49,-10'd151};
ram[8433] = {9'd52,-10'd148};
ram[8434] = {9'd55,-10'd145};
ram[8435] = {9'd58,-10'd142};
ram[8436] = {9'd62,-10'd139};
ram[8437] = {9'd65,-10'd136};
ram[8438] = {9'd68,-10'd132};
ram[8439] = {9'd71,-10'd129};
ram[8440] = {9'd74,-10'd126};
ram[8441] = {9'd77,-10'd123};
ram[8442] = {9'd80,-10'd120};
ram[8443] = {9'd84,-10'd117};
ram[8444] = {9'd87,-10'd114};
ram[8445] = {9'd90,-10'd110};
ram[8446] = {9'd93,-10'd107};
ram[8447] = {9'd96,-10'd104};
ram[8448] = {9'd96,-10'd104};
ram[8449] = {9'd99,-10'd101};
ram[8450] = {-9'd98,-10'd98};
ram[8451] = {-9'd95,-10'd95};
ram[8452] = {-9'd92,-10'd92};
ram[8453] = {-9'd88,-10'd88};
ram[8454] = {-9'd85,-10'd85};
ram[8455] = {-9'd82,-10'd82};
ram[8456] = {-9'd79,-10'd79};
ram[8457] = {-9'd76,-10'd76};
ram[8458] = {-9'd73,-10'd73};
ram[8459] = {-9'd70,-10'd70};
ram[8460] = {-9'd66,-10'd66};
ram[8461] = {-9'd63,-10'd63};
ram[8462] = {-9'd60,-10'd60};
ram[8463] = {-9'd57,-10'd57};
ram[8464] = {-9'd54,-10'd54};
ram[8465] = {-9'd51,-10'd51};
ram[8466] = {-9'd48,-10'd48};
ram[8467] = {-9'd44,-10'd44};
ram[8468] = {-9'd41,-10'd41};
ram[8469] = {-9'd38,-10'd38};
ram[8470] = {-9'd35,-10'd35};
ram[8471] = {-9'd32,-10'd32};
ram[8472] = {-9'd29,-10'd29};
ram[8473] = {-9'd26,-10'd26};
ram[8474] = {-9'd22,-10'd22};
ram[8475] = {-9'd19,-10'd19};
ram[8476] = {-9'd16,-10'd16};
ram[8477] = {-9'd13,-10'd13};
ram[8478] = {-9'd10,-10'd10};
ram[8479] = {-9'd7,-10'd7};
ram[8480] = {-9'd4,-10'd4};
ram[8481] = {9'd0,10'd0};
ram[8482] = {9'd3,10'd3};
ram[8483] = {9'd6,10'd6};
ram[8484] = {9'd9,10'd9};
ram[8485] = {9'd12,10'd12};
ram[8486] = {9'd15,10'd15};
ram[8487] = {9'd18,10'd18};
ram[8488] = {9'd21,10'd21};
ram[8489] = {9'd25,10'd25};
ram[8490] = {9'd28,10'd28};
ram[8491] = {9'd31,10'd31};
ram[8492] = {9'd34,10'd34};
ram[8493] = {9'd37,10'd37};
ram[8494] = {9'd40,10'd40};
ram[8495] = {9'd43,10'd43};
ram[8496] = {9'd47,10'd47};
ram[8497] = {9'd50,10'd50};
ram[8498] = {9'd53,10'd53};
ram[8499] = {9'd56,10'd56};
ram[8500] = {9'd59,10'd59};
ram[8501] = {9'd62,10'd62};
ram[8502] = {9'd65,10'd65};
ram[8503] = {9'd69,10'd69};
ram[8504] = {9'd72,10'd72};
ram[8505] = {9'd75,10'd75};
ram[8506] = {9'd78,10'd78};
ram[8507] = {9'd81,10'd81};
ram[8508] = {9'd84,10'd84};
ram[8509] = {9'd87,10'd87};
ram[8510] = {9'd91,10'd91};
ram[8511] = {9'd94,10'd94};
ram[8512] = {9'd97,10'd97};
ram[8513] = {-9'd100,10'd100};
ram[8514] = {-9'd97,10'd103};
ram[8515] = {-9'd94,10'd106};
ram[8516] = {-9'd91,10'd109};
ram[8517] = {-9'd88,10'd113};
ram[8518] = {-9'd85,10'd116};
ram[8519] = {-9'd81,10'd119};
ram[8520] = {-9'd78,10'd122};
ram[8521] = {-9'd75,10'd125};
ram[8522] = {-9'd72,10'd128};
ram[8523] = {-9'd69,10'd131};
ram[8524] = {-9'd66,10'd135};
ram[8525] = {-9'd63,10'd138};
ram[8526] = {-9'd59,10'd141};
ram[8527] = {-9'd56,10'd144};
ram[8528] = {-9'd53,10'd147};
ram[8529] = {-9'd50,10'd150};
ram[8530] = {-9'd47,10'd153};
ram[8531] = {-9'd44,10'd157};
ram[8532] = {-9'd41,10'd160};
ram[8533] = {-9'd37,10'd163};
ram[8534] = {-9'd34,10'd166};
ram[8535] = {-9'd31,10'd169};
ram[8536] = {-9'd28,10'd172};
ram[8537] = {-9'd25,10'd175};
ram[8538] = {-9'd22,10'd179};
ram[8539] = {-9'd19,10'd182};
ram[8540] = {-9'd15,10'd185};
ram[8541] = {-9'd12,10'd188};
ram[8542] = {-9'd9,10'd191};
ram[8543] = {-9'd6,10'd194};
ram[8544] = {-9'd3,10'd197};
ram[8545] = {9'd0,10'd201};
ram[8546] = {9'd3,10'd204};
ram[8547] = {9'd7,10'd207};
ram[8548] = {9'd10,10'd210};
ram[8549] = {9'd13,10'd213};
ram[8550] = {9'd16,10'd216};
ram[8551] = {9'd19,10'd219};
ram[8552] = {9'd22,10'd223};
ram[8553] = {9'd25,10'd226};
ram[8554] = {9'd29,10'd229};
ram[8555] = {9'd32,10'd232};
ram[8556] = {9'd35,10'd235};
ram[8557] = {9'd38,10'd238};
ram[8558] = {9'd41,10'd241};
ram[8559] = {9'd44,10'd245};
ram[8560] = {9'd47,10'd248};
ram[8561] = {9'd51,10'd251};
ram[8562] = {9'd54,10'd254};
ram[8563] = {9'd57,10'd257};
ram[8564] = {9'd60,10'd260};
ram[8565] = {9'd63,10'd263};
ram[8566] = {9'd66,10'd267};
ram[8567] = {9'd69,10'd270};
ram[8568] = {9'd73,10'd273};
ram[8569] = {9'd76,10'd276};
ram[8570] = {9'd79,10'd279};
ram[8571] = {9'd82,10'd282};
ram[8572] = {9'd85,10'd285};
ram[8573] = {9'd88,10'd289};
ram[8574] = {9'd91,10'd292};
ram[8575] = {9'd95,10'd295};
ram[8576] = {9'd95,10'd295};
ram[8577] = {9'd98,10'd298};
ram[8578] = {-9'd99,10'd301};
ram[8579] = {-9'd96,10'd304};
ram[8580] = {-9'd93,10'd307};
ram[8581] = {-9'd90,10'd311};
ram[8582] = {-9'd87,10'd314};
ram[8583] = {-9'd84,10'd317};
ram[8584] = {-9'd81,10'd320};
ram[8585] = {-9'd77,10'd323};
ram[8586] = {-9'd74,10'd326};
ram[8587] = {-9'd71,10'd329};
ram[8588] = {-9'd68,10'd333};
ram[8589] = {-9'd65,10'd336};
ram[8590] = {-9'd62,10'd339};
ram[8591] = {-9'd59,10'd342};
ram[8592] = {-9'd55,10'd345};
ram[8593] = {-9'd52,10'd348};
ram[8594] = {-9'd49,10'd351};
ram[8595] = {-9'd46,10'd354};
ram[8596] = {-9'd43,10'd358};
ram[8597] = {-9'd40,10'd361};
ram[8598] = {-9'd37,10'd364};
ram[8599] = {-9'd33,10'd367};
ram[8600] = {-9'd30,10'd370};
ram[8601] = {-9'd27,10'd373};
ram[8602] = {-9'd24,10'd376};
ram[8603] = {-9'd21,10'd380};
ram[8604] = {-9'd18,10'd383};
ram[8605] = {-9'd15,10'd386};
ram[8606] = {-9'd11,10'd389};
ram[8607] = {-9'd8,10'd392};
ram[8608] = {-9'd5,10'd395};
ram[8609] = {-9'd2,10'd398};
ram[8610] = {9'd1,-10'd399};
ram[8611] = {9'd4,-10'd396};
ram[8612] = {9'd7,-10'd393};
ram[8613] = {9'd10,-10'd390};
ram[8614] = {9'd14,-10'd387};
ram[8615] = {9'd17,-10'd384};
ram[8616] = {9'd20,-10'd381};
ram[8617] = {9'd23,-10'd377};
ram[8618] = {9'd26,-10'd374};
ram[8619] = {9'd29,-10'd371};
ram[8620] = {9'd32,-10'd368};
ram[8621] = {9'd36,-10'd365};
ram[8622] = {9'd39,-10'd362};
ram[8623] = {9'd42,-10'd359};
ram[8624] = {9'd45,-10'd355};
ram[8625] = {9'd48,-10'd352};
ram[8626] = {9'd51,-10'd349};
ram[8627] = {9'd54,-10'd346};
ram[8628] = {9'd58,-10'd343};
ram[8629] = {9'd61,-10'd340};
ram[8630] = {9'd64,-10'd337};
ram[8631] = {9'd67,-10'd334};
ram[8632] = {9'd70,-10'd330};
ram[8633] = {9'd73,-10'd327};
ram[8634] = {9'd76,-10'd324};
ram[8635] = {9'd80,-10'd321};
ram[8636] = {9'd83,-10'd318};
ram[8637] = {9'd86,-10'd315};
ram[8638] = {9'd89,-10'd312};
ram[8639] = {9'd92,-10'd308};
ram[8640] = {9'd95,-10'd305};
ram[8641] = {9'd98,-10'd302};
ram[8642] = {-9'd99,-10'd299};
ram[8643] = {-9'd96,-10'd296};
ram[8644] = {-9'd92,-10'd293};
ram[8645] = {-9'd89,-10'd290};
ram[8646] = {-9'd86,-10'd286};
ram[8647] = {-9'd83,-10'd283};
ram[8648] = {-9'd80,-10'd280};
ram[8649] = {-9'd77,-10'd277};
ram[8650] = {-9'd74,-10'd274};
ram[8651] = {-9'd70,-10'd271};
ram[8652] = {-9'd67,-10'd268};
ram[8653] = {-9'd64,-10'd264};
ram[8654] = {-9'd61,-10'd261};
ram[8655] = {-9'd58,-10'd258};
ram[8656] = {-9'd55,-10'd255};
ram[8657] = {-9'd52,-10'd252};
ram[8658] = {-9'd48,-10'd249};
ram[8659] = {-9'd45,-10'd246};
ram[8660] = {-9'd42,-10'd242};
ram[8661] = {-9'd39,-10'd239};
ram[8662] = {-9'd36,-10'd236};
ram[8663] = {-9'd33,-10'd233};
ram[8664] = {-9'd30,-10'd230};
ram[8665] = {-9'd26,-10'd227};
ram[8666] = {-9'd23,-10'd224};
ram[8667] = {-9'd20,-10'd220};
ram[8668] = {-9'd17,-10'd217};
ram[8669] = {-9'd14,-10'd214};
ram[8670] = {-9'd11,-10'd211};
ram[8671] = {-9'd8,-10'd208};
ram[8672] = {-9'd4,-10'd205};
ram[8673] = {-9'd1,-10'd202};
ram[8674] = {9'd2,-10'd198};
ram[8675] = {9'd5,-10'd195};
ram[8676] = {9'd8,-10'd192};
ram[8677] = {9'd11,-10'd189};
ram[8678] = {9'd14,-10'd186};
ram[8679] = {9'd18,-10'd183};
ram[8680] = {9'd21,-10'd180};
ram[8681] = {9'd24,-10'd176};
ram[8682] = {9'd27,-10'd173};
ram[8683] = {9'd30,-10'd170};
ram[8684] = {9'd33,-10'd167};
ram[8685] = {9'd36,-10'd164};
ram[8686] = {9'd40,-10'd161};
ram[8687] = {9'd43,-10'd158};
ram[8688] = {9'd46,-10'd154};
ram[8689] = {9'd49,-10'd151};
ram[8690] = {9'd52,-10'd148};
ram[8691] = {9'd55,-10'd145};
ram[8692] = {9'd58,-10'd142};
ram[8693] = {9'd62,-10'd139};
ram[8694] = {9'd65,-10'd136};
ram[8695] = {9'd68,-10'd132};
ram[8696] = {9'd71,-10'd129};
ram[8697] = {9'd74,-10'd126};
ram[8698] = {9'd77,-10'd123};
ram[8699] = {9'd80,-10'd120};
ram[8700] = {9'd84,-10'd117};
ram[8701] = {9'd87,-10'd114};
ram[8702] = {9'd90,-10'd110};
ram[8703] = {9'd93,-10'd107};
ram[8704] = {9'd93,-10'd107};
ram[8705] = {9'd96,-10'd104};
ram[8706] = {9'd99,-10'd101};
ram[8707] = {-9'd98,-10'd98};
ram[8708] = {-9'd95,-10'd95};
ram[8709] = {-9'd92,-10'd92};
ram[8710] = {-9'd88,-10'd88};
ram[8711] = {-9'd85,-10'd85};
ram[8712] = {-9'd82,-10'd82};
ram[8713] = {-9'd79,-10'd79};
ram[8714] = {-9'd76,-10'd76};
ram[8715] = {-9'd73,-10'd73};
ram[8716] = {-9'd70,-10'd70};
ram[8717] = {-9'd66,-10'd66};
ram[8718] = {-9'd63,-10'd63};
ram[8719] = {-9'd60,-10'd60};
ram[8720] = {-9'd57,-10'd57};
ram[8721] = {-9'd54,-10'd54};
ram[8722] = {-9'd51,-10'd51};
ram[8723] = {-9'd48,-10'd48};
ram[8724] = {-9'd44,-10'd44};
ram[8725] = {-9'd41,-10'd41};
ram[8726] = {-9'd38,-10'd38};
ram[8727] = {-9'd35,-10'd35};
ram[8728] = {-9'd32,-10'd32};
ram[8729] = {-9'd29,-10'd29};
ram[8730] = {-9'd26,-10'd26};
ram[8731] = {-9'd22,-10'd22};
ram[8732] = {-9'd19,-10'd19};
ram[8733] = {-9'd16,-10'd16};
ram[8734] = {-9'd13,-10'd13};
ram[8735] = {-9'd10,-10'd10};
ram[8736] = {-9'd7,-10'd7};
ram[8737] = {-9'd4,-10'd4};
ram[8738] = {9'd0,10'd0};
ram[8739] = {9'd3,10'd3};
ram[8740] = {9'd6,10'd6};
ram[8741] = {9'd9,10'd9};
ram[8742] = {9'd12,10'd12};
ram[8743] = {9'd15,10'd15};
ram[8744] = {9'd18,10'd18};
ram[8745] = {9'd21,10'd21};
ram[8746] = {9'd25,10'd25};
ram[8747] = {9'd28,10'd28};
ram[8748] = {9'd31,10'd31};
ram[8749] = {9'd34,10'd34};
ram[8750] = {9'd37,10'd37};
ram[8751] = {9'd40,10'd40};
ram[8752] = {9'd43,10'd43};
ram[8753] = {9'd47,10'd47};
ram[8754] = {9'd50,10'd50};
ram[8755] = {9'd53,10'd53};
ram[8756] = {9'd56,10'd56};
ram[8757] = {9'd59,10'd59};
ram[8758] = {9'd62,10'd62};
ram[8759] = {9'd65,10'd65};
ram[8760] = {9'd69,10'd69};
ram[8761] = {9'd72,10'd72};
ram[8762] = {9'd75,10'd75};
ram[8763] = {9'd78,10'd78};
ram[8764] = {9'd81,10'd81};
ram[8765] = {9'd84,10'd84};
ram[8766] = {9'd87,10'd87};
ram[8767] = {9'd91,10'd91};
ram[8768] = {9'd94,10'd94};
ram[8769] = {9'd97,10'd97};
ram[8770] = {-9'd100,10'd100};
ram[8771] = {-9'd97,10'd103};
ram[8772] = {-9'd94,10'd106};
ram[8773] = {-9'd91,10'd109};
ram[8774] = {-9'd88,10'd113};
ram[8775] = {-9'd85,10'd116};
ram[8776] = {-9'd81,10'd119};
ram[8777] = {-9'd78,10'd122};
ram[8778] = {-9'd75,10'd125};
ram[8779] = {-9'd72,10'd128};
ram[8780] = {-9'd69,10'd131};
ram[8781] = {-9'd66,10'd135};
ram[8782] = {-9'd63,10'd138};
ram[8783] = {-9'd59,10'd141};
ram[8784] = {-9'd56,10'd144};
ram[8785] = {-9'd53,10'd147};
ram[8786] = {-9'd50,10'd150};
ram[8787] = {-9'd47,10'd153};
ram[8788] = {-9'd44,10'd157};
ram[8789] = {-9'd41,10'd160};
ram[8790] = {-9'd37,10'd163};
ram[8791] = {-9'd34,10'd166};
ram[8792] = {-9'd31,10'd169};
ram[8793] = {-9'd28,10'd172};
ram[8794] = {-9'd25,10'd175};
ram[8795] = {-9'd22,10'd179};
ram[8796] = {-9'd19,10'd182};
ram[8797] = {-9'd15,10'd185};
ram[8798] = {-9'd12,10'd188};
ram[8799] = {-9'd9,10'd191};
ram[8800] = {-9'd6,10'd194};
ram[8801] = {-9'd3,10'd197};
ram[8802] = {9'd0,10'd201};
ram[8803] = {9'd3,10'd204};
ram[8804] = {9'd7,10'd207};
ram[8805] = {9'd10,10'd210};
ram[8806] = {9'd13,10'd213};
ram[8807] = {9'd16,10'd216};
ram[8808] = {9'd19,10'd219};
ram[8809] = {9'd22,10'd223};
ram[8810] = {9'd25,10'd226};
ram[8811] = {9'd29,10'd229};
ram[8812] = {9'd32,10'd232};
ram[8813] = {9'd35,10'd235};
ram[8814] = {9'd38,10'd238};
ram[8815] = {9'd41,10'd241};
ram[8816] = {9'd44,10'd245};
ram[8817] = {9'd47,10'd248};
ram[8818] = {9'd51,10'd251};
ram[8819] = {9'd54,10'd254};
ram[8820] = {9'd57,10'd257};
ram[8821] = {9'd60,10'd260};
ram[8822] = {9'd63,10'd263};
ram[8823] = {9'd66,10'd267};
ram[8824] = {9'd69,10'd270};
ram[8825] = {9'd73,10'd273};
ram[8826] = {9'd76,10'd276};
ram[8827] = {9'd79,10'd279};
ram[8828] = {9'd82,10'd282};
ram[8829] = {9'd85,10'd285};
ram[8830] = {9'd88,10'd289};
ram[8831] = {9'd91,10'd292};
ram[8832] = {9'd91,10'd292};
ram[8833] = {9'd95,10'd295};
ram[8834] = {9'd98,10'd298};
ram[8835] = {-9'd99,10'd301};
ram[8836] = {-9'd96,10'd304};
ram[8837] = {-9'd93,10'd307};
ram[8838] = {-9'd90,10'd311};
ram[8839] = {-9'd87,10'd314};
ram[8840] = {-9'd84,10'd317};
ram[8841] = {-9'd81,10'd320};
ram[8842] = {-9'd77,10'd323};
ram[8843] = {-9'd74,10'd326};
ram[8844] = {-9'd71,10'd329};
ram[8845] = {-9'd68,10'd333};
ram[8846] = {-9'd65,10'd336};
ram[8847] = {-9'd62,10'd339};
ram[8848] = {-9'd59,10'd342};
ram[8849] = {-9'd55,10'd345};
ram[8850] = {-9'd52,10'd348};
ram[8851] = {-9'd49,10'd351};
ram[8852] = {-9'd46,10'd354};
ram[8853] = {-9'd43,10'd358};
ram[8854] = {-9'd40,10'd361};
ram[8855] = {-9'd37,10'd364};
ram[8856] = {-9'd33,10'd367};
ram[8857] = {-9'd30,10'd370};
ram[8858] = {-9'd27,10'd373};
ram[8859] = {-9'd24,10'd376};
ram[8860] = {-9'd21,10'd380};
ram[8861] = {-9'd18,10'd383};
ram[8862] = {-9'd15,10'd386};
ram[8863] = {-9'd11,10'd389};
ram[8864] = {-9'd8,10'd392};
ram[8865] = {-9'd5,10'd395};
ram[8866] = {-9'd2,10'd398};
ram[8867] = {9'd1,-10'd399};
ram[8868] = {9'd4,-10'd396};
ram[8869] = {9'd7,-10'd393};
ram[8870] = {9'd10,-10'd390};
ram[8871] = {9'd14,-10'd387};
ram[8872] = {9'd17,-10'd384};
ram[8873] = {9'd20,-10'd381};
ram[8874] = {9'd23,-10'd377};
ram[8875] = {9'd26,-10'd374};
ram[8876] = {9'd29,-10'd371};
ram[8877] = {9'd32,-10'd368};
ram[8878] = {9'd36,-10'd365};
ram[8879] = {9'd39,-10'd362};
ram[8880] = {9'd42,-10'd359};
ram[8881] = {9'd45,-10'd355};
ram[8882] = {9'd48,-10'd352};
ram[8883] = {9'd51,-10'd349};
ram[8884] = {9'd54,-10'd346};
ram[8885] = {9'd58,-10'd343};
ram[8886] = {9'd61,-10'd340};
ram[8887] = {9'd64,-10'd337};
ram[8888] = {9'd67,-10'd334};
ram[8889] = {9'd70,-10'd330};
ram[8890] = {9'd73,-10'd327};
ram[8891] = {9'd76,-10'd324};
ram[8892] = {9'd80,-10'd321};
ram[8893] = {9'd83,-10'd318};
ram[8894] = {9'd86,-10'd315};
ram[8895] = {9'd89,-10'd312};
ram[8896] = {9'd92,-10'd308};
ram[8897] = {9'd95,-10'd305};
ram[8898] = {9'd98,-10'd302};
ram[8899] = {-9'd99,-10'd299};
ram[8900] = {-9'd96,-10'd296};
ram[8901] = {-9'd92,-10'd293};
ram[8902] = {-9'd89,-10'd290};
ram[8903] = {-9'd86,-10'd286};
ram[8904] = {-9'd83,-10'd283};
ram[8905] = {-9'd80,-10'd280};
ram[8906] = {-9'd77,-10'd277};
ram[8907] = {-9'd74,-10'd274};
ram[8908] = {-9'd70,-10'd271};
ram[8909] = {-9'd67,-10'd268};
ram[8910] = {-9'd64,-10'd264};
ram[8911] = {-9'd61,-10'd261};
ram[8912] = {-9'd58,-10'd258};
ram[8913] = {-9'd55,-10'd255};
ram[8914] = {-9'd52,-10'd252};
ram[8915] = {-9'd48,-10'd249};
ram[8916] = {-9'd45,-10'd246};
ram[8917] = {-9'd42,-10'd242};
ram[8918] = {-9'd39,-10'd239};
ram[8919] = {-9'd36,-10'd236};
ram[8920] = {-9'd33,-10'd233};
ram[8921] = {-9'd30,-10'd230};
ram[8922] = {-9'd26,-10'd227};
ram[8923] = {-9'd23,-10'd224};
ram[8924] = {-9'd20,-10'd220};
ram[8925] = {-9'd17,-10'd217};
ram[8926] = {-9'd14,-10'd214};
ram[8927] = {-9'd11,-10'd211};
ram[8928] = {-9'd8,-10'd208};
ram[8929] = {-9'd4,-10'd205};
ram[8930] = {-9'd1,-10'd202};
ram[8931] = {9'd2,-10'd198};
ram[8932] = {9'd5,-10'd195};
ram[8933] = {9'd8,-10'd192};
ram[8934] = {9'd11,-10'd189};
ram[8935] = {9'd14,-10'd186};
ram[8936] = {9'd18,-10'd183};
ram[8937] = {9'd21,-10'd180};
ram[8938] = {9'd24,-10'd176};
ram[8939] = {9'd27,-10'd173};
ram[8940] = {9'd30,-10'd170};
ram[8941] = {9'd33,-10'd167};
ram[8942] = {9'd36,-10'd164};
ram[8943] = {9'd40,-10'd161};
ram[8944] = {9'd43,-10'd158};
ram[8945] = {9'd46,-10'd154};
ram[8946] = {9'd49,-10'd151};
ram[8947] = {9'd52,-10'd148};
ram[8948] = {9'd55,-10'd145};
ram[8949] = {9'd58,-10'd142};
ram[8950] = {9'd62,-10'd139};
ram[8951] = {9'd65,-10'd136};
ram[8952] = {9'd68,-10'd132};
ram[8953] = {9'd71,-10'd129};
ram[8954] = {9'd74,-10'd126};
ram[8955] = {9'd77,-10'd123};
ram[8956] = {9'd80,-10'd120};
ram[8957] = {9'd84,-10'd117};
ram[8958] = {9'd87,-10'd114};
ram[8959] = {9'd90,-10'd110};
ram[8960] = {9'd90,-10'd110};
ram[8961] = {9'd93,-10'd107};
ram[8962] = {9'd96,-10'd104};
ram[8963] = {9'd99,-10'd101};
ram[8964] = {-9'd98,-10'd98};
ram[8965] = {-9'd95,-10'd95};
ram[8966] = {-9'd92,-10'd92};
ram[8967] = {-9'd88,-10'd88};
ram[8968] = {-9'd85,-10'd85};
ram[8969] = {-9'd82,-10'd82};
ram[8970] = {-9'd79,-10'd79};
ram[8971] = {-9'd76,-10'd76};
ram[8972] = {-9'd73,-10'd73};
ram[8973] = {-9'd70,-10'd70};
ram[8974] = {-9'd66,-10'd66};
ram[8975] = {-9'd63,-10'd63};
ram[8976] = {-9'd60,-10'd60};
ram[8977] = {-9'd57,-10'd57};
ram[8978] = {-9'd54,-10'd54};
ram[8979] = {-9'd51,-10'd51};
ram[8980] = {-9'd48,-10'd48};
ram[8981] = {-9'd44,-10'd44};
ram[8982] = {-9'd41,-10'd41};
ram[8983] = {-9'd38,-10'd38};
ram[8984] = {-9'd35,-10'd35};
ram[8985] = {-9'd32,-10'd32};
ram[8986] = {-9'd29,-10'd29};
ram[8987] = {-9'd26,-10'd26};
ram[8988] = {-9'd22,-10'd22};
ram[8989] = {-9'd19,-10'd19};
ram[8990] = {-9'd16,-10'd16};
ram[8991] = {-9'd13,-10'd13};
ram[8992] = {-9'd10,-10'd10};
ram[8993] = {-9'd7,-10'd7};
ram[8994] = {-9'd4,-10'd4};
ram[8995] = {9'd0,10'd0};
ram[8996] = {9'd3,10'd3};
ram[8997] = {9'd6,10'd6};
ram[8998] = {9'd9,10'd9};
ram[8999] = {9'd12,10'd12};
ram[9000] = {9'd15,10'd15};
ram[9001] = {9'd18,10'd18};
ram[9002] = {9'd21,10'd21};
ram[9003] = {9'd25,10'd25};
ram[9004] = {9'd28,10'd28};
ram[9005] = {9'd31,10'd31};
ram[9006] = {9'd34,10'd34};
ram[9007] = {9'd37,10'd37};
ram[9008] = {9'd40,10'd40};
ram[9009] = {9'd43,10'd43};
ram[9010] = {9'd47,10'd47};
ram[9011] = {9'd50,10'd50};
ram[9012] = {9'd53,10'd53};
ram[9013] = {9'd56,10'd56};
ram[9014] = {9'd59,10'd59};
ram[9015] = {9'd62,10'd62};
ram[9016] = {9'd65,10'd65};
ram[9017] = {9'd69,10'd69};
ram[9018] = {9'd72,10'd72};
ram[9019] = {9'd75,10'd75};
ram[9020] = {9'd78,10'd78};
ram[9021] = {9'd81,10'd81};
ram[9022] = {9'd84,10'd84};
ram[9023] = {9'd87,10'd87};
ram[9024] = {9'd91,10'd91};
ram[9025] = {9'd94,10'd94};
ram[9026] = {9'd97,10'd97};
ram[9027] = {-9'd100,10'd100};
ram[9028] = {-9'd97,10'd103};
ram[9029] = {-9'd94,10'd106};
ram[9030] = {-9'd91,10'd109};
ram[9031] = {-9'd88,10'd113};
ram[9032] = {-9'd85,10'd116};
ram[9033] = {-9'd81,10'd119};
ram[9034] = {-9'd78,10'd122};
ram[9035] = {-9'd75,10'd125};
ram[9036] = {-9'd72,10'd128};
ram[9037] = {-9'd69,10'd131};
ram[9038] = {-9'd66,10'd135};
ram[9039] = {-9'd63,10'd138};
ram[9040] = {-9'd59,10'd141};
ram[9041] = {-9'd56,10'd144};
ram[9042] = {-9'd53,10'd147};
ram[9043] = {-9'd50,10'd150};
ram[9044] = {-9'd47,10'd153};
ram[9045] = {-9'd44,10'd157};
ram[9046] = {-9'd41,10'd160};
ram[9047] = {-9'd37,10'd163};
ram[9048] = {-9'd34,10'd166};
ram[9049] = {-9'd31,10'd169};
ram[9050] = {-9'd28,10'd172};
ram[9051] = {-9'd25,10'd175};
ram[9052] = {-9'd22,10'd179};
ram[9053] = {-9'd19,10'd182};
ram[9054] = {-9'd15,10'd185};
ram[9055] = {-9'd12,10'd188};
ram[9056] = {-9'd9,10'd191};
ram[9057] = {-9'd6,10'd194};
ram[9058] = {-9'd3,10'd197};
ram[9059] = {9'd0,10'd201};
ram[9060] = {9'd3,10'd204};
ram[9061] = {9'd7,10'd207};
ram[9062] = {9'd10,10'd210};
ram[9063] = {9'd13,10'd213};
ram[9064] = {9'd16,10'd216};
ram[9065] = {9'd19,10'd219};
ram[9066] = {9'd22,10'd223};
ram[9067] = {9'd25,10'd226};
ram[9068] = {9'd29,10'd229};
ram[9069] = {9'd32,10'd232};
ram[9070] = {9'd35,10'd235};
ram[9071] = {9'd38,10'd238};
ram[9072] = {9'd41,10'd241};
ram[9073] = {9'd44,10'd245};
ram[9074] = {9'd47,10'd248};
ram[9075] = {9'd51,10'd251};
ram[9076] = {9'd54,10'd254};
ram[9077] = {9'd57,10'd257};
ram[9078] = {9'd60,10'd260};
ram[9079] = {9'd63,10'd263};
ram[9080] = {9'd66,10'd267};
ram[9081] = {9'd69,10'd270};
ram[9082] = {9'd73,10'd273};
ram[9083] = {9'd76,10'd276};
ram[9084] = {9'd79,10'd279};
ram[9085] = {9'd82,10'd282};
ram[9086] = {9'd85,10'd285};
ram[9087] = {9'd88,10'd289};
ram[9088] = {9'd88,10'd289};
ram[9089] = {9'd91,10'd292};
ram[9090] = {9'd95,10'd295};
ram[9091] = {9'd98,10'd298};
ram[9092] = {-9'd99,10'd301};
ram[9093] = {-9'd96,10'd304};
ram[9094] = {-9'd93,10'd307};
ram[9095] = {-9'd90,10'd311};
ram[9096] = {-9'd87,10'd314};
ram[9097] = {-9'd84,10'd317};
ram[9098] = {-9'd81,10'd320};
ram[9099] = {-9'd77,10'd323};
ram[9100] = {-9'd74,10'd326};
ram[9101] = {-9'd71,10'd329};
ram[9102] = {-9'd68,10'd333};
ram[9103] = {-9'd65,10'd336};
ram[9104] = {-9'd62,10'd339};
ram[9105] = {-9'd59,10'd342};
ram[9106] = {-9'd55,10'd345};
ram[9107] = {-9'd52,10'd348};
ram[9108] = {-9'd49,10'd351};
ram[9109] = {-9'd46,10'd354};
ram[9110] = {-9'd43,10'd358};
ram[9111] = {-9'd40,10'd361};
ram[9112] = {-9'd37,10'd364};
ram[9113] = {-9'd33,10'd367};
ram[9114] = {-9'd30,10'd370};
ram[9115] = {-9'd27,10'd373};
ram[9116] = {-9'd24,10'd376};
ram[9117] = {-9'd21,10'd380};
ram[9118] = {-9'd18,10'd383};
ram[9119] = {-9'd15,10'd386};
ram[9120] = {-9'd11,10'd389};
ram[9121] = {-9'd8,10'd392};
ram[9122] = {-9'd5,10'd395};
ram[9123] = {-9'd2,10'd398};
ram[9124] = {9'd1,-10'd399};
ram[9125] = {9'd4,-10'd396};
ram[9126] = {9'd7,-10'd393};
ram[9127] = {9'd10,-10'd390};
ram[9128] = {9'd14,-10'd387};
ram[9129] = {9'd17,-10'd384};
ram[9130] = {9'd20,-10'd381};
ram[9131] = {9'd23,-10'd377};
ram[9132] = {9'd26,-10'd374};
ram[9133] = {9'd29,-10'd371};
ram[9134] = {9'd32,-10'd368};
ram[9135] = {9'd36,-10'd365};
ram[9136] = {9'd39,-10'd362};
ram[9137] = {9'd42,-10'd359};
ram[9138] = {9'd45,-10'd355};
ram[9139] = {9'd48,-10'd352};
ram[9140] = {9'd51,-10'd349};
ram[9141] = {9'd54,-10'd346};
ram[9142] = {9'd58,-10'd343};
ram[9143] = {9'd61,-10'd340};
ram[9144] = {9'd64,-10'd337};
ram[9145] = {9'd67,-10'd334};
ram[9146] = {9'd70,-10'd330};
ram[9147] = {9'd73,-10'd327};
ram[9148] = {9'd76,-10'd324};
ram[9149] = {9'd80,-10'd321};
ram[9150] = {9'd83,-10'd318};
ram[9151] = {9'd86,-10'd315};
ram[9152] = {9'd89,-10'd312};
ram[9153] = {9'd92,-10'd308};
ram[9154] = {9'd95,-10'd305};
ram[9155] = {9'd98,-10'd302};
ram[9156] = {-9'd99,-10'd299};
ram[9157] = {-9'd96,-10'd296};
ram[9158] = {-9'd92,-10'd293};
ram[9159] = {-9'd89,-10'd290};
ram[9160] = {-9'd86,-10'd286};
ram[9161] = {-9'd83,-10'd283};
ram[9162] = {-9'd80,-10'd280};
ram[9163] = {-9'd77,-10'd277};
ram[9164] = {-9'd74,-10'd274};
ram[9165] = {-9'd70,-10'd271};
ram[9166] = {-9'd67,-10'd268};
ram[9167] = {-9'd64,-10'd264};
ram[9168] = {-9'd61,-10'd261};
ram[9169] = {-9'd58,-10'd258};
ram[9170] = {-9'd55,-10'd255};
ram[9171] = {-9'd52,-10'd252};
ram[9172] = {-9'd48,-10'd249};
ram[9173] = {-9'd45,-10'd246};
ram[9174] = {-9'd42,-10'd242};
ram[9175] = {-9'd39,-10'd239};
ram[9176] = {-9'd36,-10'd236};
ram[9177] = {-9'd33,-10'd233};
ram[9178] = {-9'd30,-10'd230};
ram[9179] = {-9'd26,-10'd227};
ram[9180] = {-9'd23,-10'd224};
ram[9181] = {-9'd20,-10'd220};
ram[9182] = {-9'd17,-10'd217};
ram[9183] = {-9'd14,-10'd214};
ram[9184] = {-9'd11,-10'd211};
ram[9185] = {-9'd8,-10'd208};
ram[9186] = {-9'd4,-10'd205};
ram[9187] = {-9'd1,-10'd202};
ram[9188] = {9'd2,-10'd198};
ram[9189] = {9'd5,-10'd195};
ram[9190] = {9'd8,-10'd192};
ram[9191] = {9'd11,-10'd189};
ram[9192] = {9'd14,-10'd186};
ram[9193] = {9'd18,-10'd183};
ram[9194] = {9'd21,-10'd180};
ram[9195] = {9'd24,-10'd176};
ram[9196] = {9'd27,-10'd173};
ram[9197] = {9'd30,-10'd170};
ram[9198] = {9'd33,-10'd167};
ram[9199] = {9'd36,-10'd164};
ram[9200] = {9'd40,-10'd161};
ram[9201] = {9'd43,-10'd158};
ram[9202] = {9'd46,-10'd154};
ram[9203] = {9'd49,-10'd151};
ram[9204] = {9'd52,-10'd148};
ram[9205] = {9'd55,-10'd145};
ram[9206] = {9'd58,-10'd142};
ram[9207] = {9'd62,-10'd139};
ram[9208] = {9'd65,-10'd136};
ram[9209] = {9'd68,-10'd132};
ram[9210] = {9'd71,-10'd129};
ram[9211] = {9'd74,-10'd126};
ram[9212] = {9'd77,-10'd123};
ram[9213] = {9'd80,-10'd120};
ram[9214] = {9'd84,-10'd117};
ram[9215] = {9'd87,-10'd114};
ram[9216] = {9'd87,-10'd114};
ram[9217] = {9'd90,-10'd110};
ram[9218] = {9'd93,-10'd107};
ram[9219] = {9'd96,-10'd104};
ram[9220] = {9'd99,-10'd101};
ram[9221] = {-9'd98,-10'd98};
ram[9222] = {-9'd95,-10'd95};
ram[9223] = {-9'd92,-10'd92};
ram[9224] = {-9'd88,-10'd88};
ram[9225] = {-9'd85,-10'd85};
ram[9226] = {-9'd82,-10'd82};
ram[9227] = {-9'd79,-10'd79};
ram[9228] = {-9'd76,-10'd76};
ram[9229] = {-9'd73,-10'd73};
ram[9230] = {-9'd70,-10'd70};
ram[9231] = {-9'd66,-10'd66};
ram[9232] = {-9'd63,-10'd63};
ram[9233] = {-9'd60,-10'd60};
ram[9234] = {-9'd57,-10'd57};
ram[9235] = {-9'd54,-10'd54};
ram[9236] = {-9'd51,-10'd51};
ram[9237] = {-9'd48,-10'd48};
ram[9238] = {-9'd44,-10'd44};
ram[9239] = {-9'd41,-10'd41};
ram[9240] = {-9'd38,-10'd38};
ram[9241] = {-9'd35,-10'd35};
ram[9242] = {-9'd32,-10'd32};
ram[9243] = {-9'd29,-10'd29};
ram[9244] = {-9'd26,-10'd26};
ram[9245] = {-9'd22,-10'd22};
ram[9246] = {-9'd19,-10'd19};
ram[9247] = {-9'd16,-10'd16};
ram[9248] = {-9'd13,-10'd13};
ram[9249] = {-9'd10,-10'd10};
ram[9250] = {-9'd7,-10'd7};
ram[9251] = {-9'd4,-10'd4};
ram[9252] = {9'd0,10'd0};
ram[9253] = {9'd3,10'd3};
ram[9254] = {9'd6,10'd6};
ram[9255] = {9'd9,10'd9};
ram[9256] = {9'd12,10'd12};
ram[9257] = {9'd15,10'd15};
ram[9258] = {9'd18,10'd18};
ram[9259] = {9'd21,10'd21};
ram[9260] = {9'd25,10'd25};
ram[9261] = {9'd28,10'd28};
ram[9262] = {9'd31,10'd31};
ram[9263] = {9'd34,10'd34};
ram[9264] = {9'd37,10'd37};
ram[9265] = {9'd40,10'd40};
ram[9266] = {9'd43,10'd43};
ram[9267] = {9'd47,10'd47};
ram[9268] = {9'd50,10'd50};
ram[9269] = {9'd53,10'd53};
ram[9270] = {9'd56,10'd56};
ram[9271] = {9'd59,10'd59};
ram[9272] = {9'd62,10'd62};
ram[9273] = {9'd65,10'd65};
ram[9274] = {9'd69,10'd69};
ram[9275] = {9'd72,10'd72};
ram[9276] = {9'd75,10'd75};
ram[9277] = {9'd78,10'd78};
ram[9278] = {9'd81,10'd81};
ram[9279] = {9'd84,10'd84};
ram[9280] = {9'd87,10'd87};
ram[9281] = {9'd91,10'd91};
ram[9282] = {9'd94,10'd94};
ram[9283] = {9'd97,10'd97};
ram[9284] = {-9'd100,10'd100};
ram[9285] = {-9'd97,10'd103};
ram[9286] = {-9'd94,10'd106};
ram[9287] = {-9'd91,10'd109};
ram[9288] = {-9'd88,10'd113};
ram[9289] = {-9'd85,10'd116};
ram[9290] = {-9'd81,10'd119};
ram[9291] = {-9'd78,10'd122};
ram[9292] = {-9'd75,10'd125};
ram[9293] = {-9'd72,10'd128};
ram[9294] = {-9'd69,10'd131};
ram[9295] = {-9'd66,10'd135};
ram[9296] = {-9'd63,10'd138};
ram[9297] = {-9'd59,10'd141};
ram[9298] = {-9'd56,10'd144};
ram[9299] = {-9'd53,10'd147};
ram[9300] = {-9'd50,10'd150};
ram[9301] = {-9'd47,10'd153};
ram[9302] = {-9'd44,10'd157};
ram[9303] = {-9'd41,10'd160};
ram[9304] = {-9'd37,10'd163};
ram[9305] = {-9'd34,10'd166};
ram[9306] = {-9'd31,10'd169};
ram[9307] = {-9'd28,10'd172};
ram[9308] = {-9'd25,10'd175};
ram[9309] = {-9'd22,10'd179};
ram[9310] = {-9'd19,10'd182};
ram[9311] = {-9'd15,10'd185};
ram[9312] = {-9'd12,10'd188};
ram[9313] = {-9'd9,10'd191};
ram[9314] = {-9'd6,10'd194};
ram[9315] = {-9'd3,10'd197};
ram[9316] = {9'd0,10'd201};
ram[9317] = {9'd3,10'd204};
ram[9318] = {9'd7,10'd207};
ram[9319] = {9'd10,10'd210};
ram[9320] = {9'd13,10'd213};
ram[9321] = {9'd16,10'd216};
ram[9322] = {9'd19,10'd219};
ram[9323] = {9'd22,10'd223};
ram[9324] = {9'd25,10'd226};
ram[9325] = {9'd29,10'd229};
ram[9326] = {9'd32,10'd232};
ram[9327] = {9'd35,10'd235};
ram[9328] = {9'd38,10'd238};
ram[9329] = {9'd41,10'd241};
ram[9330] = {9'd44,10'd245};
ram[9331] = {9'd47,10'd248};
ram[9332] = {9'd51,10'd251};
ram[9333] = {9'd54,10'd254};
ram[9334] = {9'd57,10'd257};
ram[9335] = {9'd60,10'd260};
ram[9336] = {9'd63,10'd263};
ram[9337] = {9'd66,10'd267};
ram[9338] = {9'd69,10'd270};
ram[9339] = {9'd73,10'd273};
ram[9340] = {9'd76,10'd276};
ram[9341] = {9'd79,10'd279};
ram[9342] = {9'd82,10'd282};
ram[9343] = {9'd85,10'd285};
ram[9344] = {9'd85,10'd285};
ram[9345] = {9'd88,10'd289};
ram[9346] = {9'd91,10'd292};
ram[9347] = {9'd95,10'd295};
ram[9348] = {9'd98,10'd298};
ram[9349] = {-9'd99,10'd301};
ram[9350] = {-9'd96,10'd304};
ram[9351] = {-9'd93,10'd307};
ram[9352] = {-9'd90,10'd311};
ram[9353] = {-9'd87,10'd314};
ram[9354] = {-9'd84,10'd317};
ram[9355] = {-9'd81,10'd320};
ram[9356] = {-9'd77,10'd323};
ram[9357] = {-9'd74,10'd326};
ram[9358] = {-9'd71,10'd329};
ram[9359] = {-9'd68,10'd333};
ram[9360] = {-9'd65,10'd336};
ram[9361] = {-9'd62,10'd339};
ram[9362] = {-9'd59,10'd342};
ram[9363] = {-9'd55,10'd345};
ram[9364] = {-9'd52,10'd348};
ram[9365] = {-9'd49,10'd351};
ram[9366] = {-9'd46,10'd354};
ram[9367] = {-9'd43,10'd358};
ram[9368] = {-9'd40,10'd361};
ram[9369] = {-9'd37,10'd364};
ram[9370] = {-9'd33,10'd367};
ram[9371] = {-9'd30,10'd370};
ram[9372] = {-9'd27,10'd373};
ram[9373] = {-9'd24,10'd376};
ram[9374] = {-9'd21,10'd380};
ram[9375] = {-9'd18,10'd383};
ram[9376] = {-9'd15,10'd386};
ram[9377] = {-9'd11,10'd389};
ram[9378] = {-9'd8,10'd392};
ram[9379] = {-9'd5,10'd395};
ram[9380] = {-9'd2,10'd398};
ram[9381] = {9'd1,-10'd399};
ram[9382] = {9'd4,-10'd396};
ram[9383] = {9'd7,-10'd393};
ram[9384] = {9'd10,-10'd390};
ram[9385] = {9'd14,-10'd387};
ram[9386] = {9'd17,-10'd384};
ram[9387] = {9'd20,-10'd381};
ram[9388] = {9'd23,-10'd377};
ram[9389] = {9'd26,-10'd374};
ram[9390] = {9'd29,-10'd371};
ram[9391] = {9'd32,-10'd368};
ram[9392] = {9'd36,-10'd365};
ram[9393] = {9'd39,-10'd362};
ram[9394] = {9'd42,-10'd359};
ram[9395] = {9'd45,-10'd355};
ram[9396] = {9'd48,-10'd352};
ram[9397] = {9'd51,-10'd349};
ram[9398] = {9'd54,-10'd346};
ram[9399] = {9'd58,-10'd343};
ram[9400] = {9'd61,-10'd340};
ram[9401] = {9'd64,-10'd337};
ram[9402] = {9'd67,-10'd334};
ram[9403] = {9'd70,-10'd330};
ram[9404] = {9'd73,-10'd327};
ram[9405] = {9'd76,-10'd324};
ram[9406] = {9'd80,-10'd321};
ram[9407] = {9'd83,-10'd318};
ram[9408] = {9'd86,-10'd315};
ram[9409] = {9'd89,-10'd312};
ram[9410] = {9'd92,-10'd308};
ram[9411] = {9'd95,-10'd305};
ram[9412] = {9'd98,-10'd302};
ram[9413] = {-9'd99,-10'd299};
ram[9414] = {-9'd96,-10'd296};
ram[9415] = {-9'd92,-10'd293};
ram[9416] = {-9'd89,-10'd290};
ram[9417] = {-9'd86,-10'd286};
ram[9418] = {-9'd83,-10'd283};
ram[9419] = {-9'd80,-10'd280};
ram[9420] = {-9'd77,-10'd277};
ram[9421] = {-9'd74,-10'd274};
ram[9422] = {-9'd70,-10'd271};
ram[9423] = {-9'd67,-10'd268};
ram[9424] = {-9'd64,-10'd264};
ram[9425] = {-9'd61,-10'd261};
ram[9426] = {-9'd58,-10'd258};
ram[9427] = {-9'd55,-10'd255};
ram[9428] = {-9'd52,-10'd252};
ram[9429] = {-9'd48,-10'd249};
ram[9430] = {-9'd45,-10'd246};
ram[9431] = {-9'd42,-10'd242};
ram[9432] = {-9'd39,-10'd239};
ram[9433] = {-9'd36,-10'd236};
ram[9434] = {-9'd33,-10'd233};
ram[9435] = {-9'd30,-10'd230};
ram[9436] = {-9'd26,-10'd227};
ram[9437] = {-9'd23,-10'd224};
ram[9438] = {-9'd20,-10'd220};
ram[9439] = {-9'd17,-10'd217};
ram[9440] = {-9'd14,-10'd214};
ram[9441] = {-9'd11,-10'd211};
ram[9442] = {-9'd8,-10'd208};
ram[9443] = {-9'd4,-10'd205};
ram[9444] = {-9'd1,-10'd202};
ram[9445] = {9'd2,-10'd198};
ram[9446] = {9'd5,-10'd195};
ram[9447] = {9'd8,-10'd192};
ram[9448] = {9'd11,-10'd189};
ram[9449] = {9'd14,-10'd186};
ram[9450] = {9'd18,-10'd183};
ram[9451] = {9'd21,-10'd180};
ram[9452] = {9'd24,-10'd176};
ram[9453] = {9'd27,-10'd173};
ram[9454] = {9'd30,-10'd170};
ram[9455] = {9'd33,-10'd167};
ram[9456] = {9'd36,-10'd164};
ram[9457] = {9'd40,-10'd161};
ram[9458] = {9'd43,-10'd158};
ram[9459] = {9'd46,-10'd154};
ram[9460] = {9'd49,-10'd151};
ram[9461] = {9'd52,-10'd148};
ram[9462] = {9'd55,-10'd145};
ram[9463] = {9'd58,-10'd142};
ram[9464] = {9'd62,-10'd139};
ram[9465] = {9'd65,-10'd136};
ram[9466] = {9'd68,-10'd132};
ram[9467] = {9'd71,-10'd129};
ram[9468] = {9'd74,-10'd126};
ram[9469] = {9'd77,-10'd123};
ram[9470] = {9'd80,-10'd120};
ram[9471] = {9'd84,-10'd117};
ram[9472] = {9'd84,-10'd117};
ram[9473] = {9'd87,-10'd114};
ram[9474] = {9'd90,-10'd110};
ram[9475] = {9'd93,-10'd107};
ram[9476] = {9'd96,-10'd104};
ram[9477] = {9'd99,-10'd101};
ram[9478] = {-9'd98,-10'd98};
ram[9479] = {-9'd95,-10'd95};
ram[9480] = {-9'd92,-10'd92};
ram[9481] = {-9'd88,-10'd88};
ram[9482] = {-9'd85,-10'd85};
ram[9483] = {-9'd82,-10'd82};
ram[9484] = {-9'd79,-10'd79};
ram[9485] = {-9'd76,-10'd76};
ram[9486] = {-9'd73,-10'd73};
ram[9487] = {-9'd70,-10'd70};
ram[9488] = {-9'd66,-10'd66};
ram[9489] = {-9'd63,-10'd63};
ram[9490] = {-9'd60,-10'd60};
ram[9491] = {-9'd57,-10'd57};
ram[9492] = {-9'd54,-10'd54};
ram[9493] = {-9'd51,-10'd51};
ram[9494] = {-9'd48,-10'd48};
ram[9495] = {-9'd44,-10'd44};
ram[9496] = {-9'd41,-10'd41};
ram[9497] = {-9'd38,-10'd38};
ram[9498] = {-9'd35,-10'd35};
ram[9499] = {-9'd32,-10'd32};
ram[9500] = {-9'd29,-10'd29};
ram[9501] = {-9'd26,-10'd26};
ram[9502] = {-9'd22,-10'd22};
ram[9503] = {-9'd19,-10'd19};
ram[9504] = {-9'd16,-10'd16};
ram[9505] = {-9'd13,-10'd13};
ram[9506] = {-9'd10,-10'd10};
ram[9507] = {-9'd7,-10'd7};
ram[9508] = {-9'd4,-10'd4};
ram[9509] = {9'd0,10'd0};
ram[9510] = {9'd3,10'd3};
ram[9511] = {9'd6,10'd6};
ram[9512] = {9'd9,10'd9};
ram[9513] = {9'd12,10'd12};
ram[9514] = {9'd15,10'd15};
ram[9515] = {9'd18,10'd18};
ram[9516] = {9'd21,10'd21};
ram[9517] = {9'd25,10'd25};
ram[9518] = {9'd28,10'd28};
ram[9519] = {9'd31,10'd31};
ram[9520] = {9'd34,10'd34};
ram[9521] = {9'd37,10'd37};
ram[9522] = {9'd40,10'd40};
ram[9523] = {9'd43,10'd43};
ram[9524] = {9'd47,10'd47};
ram[9525] = {9'd50,10'd50};
ram[9526] = {9'd53,10'd53};
ram[9527] = {9'd56,10'd56};
ram[9528] = {9'd59,10'd59};
ram[9529] = {9'd62,10'd62};
ram[9530] = {9'd65,10'd65};
ram[9531] = {9'd69,10'd69};
ram[9532] = {9'd72,10'd72};
ram[9533] = {9'd75,10'd75};
ram[9534] = {9'd78,10'd78};
ram[9535] = {9'd81,10'd81};
ram[9536] = {9'd84,10'd84};
ram[9537] = {9'd87,10'd87};
ram[9538] = {9'd91,10'd91};
ram[9539] = {9'd94,10'd94};
ram[9540] = {9'd97,10'd97};
ram[9541] = {-9'd100,10'd100};
ram[9542] = {-9'd97,10'd103};
ram[9543] = {-9'd94,10'd106};
ram[9544] = {-9'd91,10'd109};
ram[9545] = {-9'd88,10'd113};
ram[9546] = {-9'd85,10'd116};
ram[9547] = {-9'd81,10'd119};
ram[9548] = {-9'd78,10'd122};
ram[9549] = {-9'd75,10'd125};
ram[9550] = {-9'd72,10'd128};
ram[9551] = {-9'd69,10'd131};
ram[9552] = {-9'd66,10'd135};
ram[9553] = {-9'd63,10'd138};
ram[9554] = {-9'd59,10'd141};
ram[9555] = {-9'd56,10'd144};
ram[9556] = {-9'd53,10'd147};
ram[9557] = {-9'd50,10'd150};
ram[9558] = {-9'd47,10'd153};
ram[9559] = {-9'd44,10'd157};
ram[9560] = {-9'd41,10'd160};
ram[9561] = {-9'd37,10'd163};
ram[9562] = {-9'd34,10'd166};
ram[9563] = {-9'd31,10'd169};
ram[9564] = {-9'd28,10'd172};
ram[9565] = {-9'd25,10'd175};
ram[9566] = {-9'd22,10'd179};
ram[9567] = {-9'd19,10'd182};
ram[9568] = {-9'd15,10'd185};
ram[9569] = {-9'd12,10'd188};
ram[9570] = {-9'd9,10'd191};
ram[9571] = {-9'd6,10'd194};
ram[9572] = {-9'd3,10'd197};
ram[9573] = {9'd0,10'd201};
ram[9574] = {9'd3,10'd204};
ram[9575] = {9'd7,10'd207};
ram[9576] = {9'd10,10'd210};
ram[9577] = {9'd13,10'd213};
ram[9578] = {9'd16,10'd216};
ram[9579] = {9'd19,10'd219};
ram[9580] = {9'd22,10'd223};
ram[9581] = {9'd25,10'd226};
ram[9582] = {9'd29,10'd229};
ram[9583] = {9'd32,10'd232};
ram[9584] = {9'd35,10'd235};
ram[9585] = {9'd38,10'd238};
ram[9586] = {9'd41,10'd241};
ram[9587] = {9'd44,10'd245};
ram[9588] = {9'd47,10'd248};
ram[9589] = {9'd51,10'd251};
ram[9590] = {9'd54,10'd254};
ram[9591] = {9'd57,10'd257};
ram[9592] = {9'd60,10'd260};
ram[9593] = {9'd63,10'd263};
ram[9594] = {9'd66,10'd267};
ram[9595] = {9'd69,10'd270};
ram[9596] = {9'd73,10'd273};
ram[9597] = {9'd76,10'd276};
ram[9598] = {9'd79,10'd279};
ram[9599] = {9'd82,10'd282};
ram[9600] = {9'd82,10'd282};
ram[9601] = {9'd85,10'd285};
ram[9602] = {9'd88,10'd289};
ram[9603] = {9'd91,10'd292};
ram[9604] = {9'd95,10'd295};
ram[9605] = {9'd98,10'd298};
ram[9606] = {-9'd99,10'd301};
ram[9607] = {-9'd96,10'd304};
ram[9608] = {-9'd93,10'd307};
ram[9609] = {-9'd90,10'd311};
ram[9610] = {-9'd87,10'd314};
ram[9611] = {-9'd84,10'd317};
ram[9612] = {-9'd81,10'd320};
ram[9613] = {-9'd77,10'd323};
ram[9614] = {-9'd74,10'd326};
ram[9615] = {-9'd71,10'd329};
ram[9616] = {-9'd68,10'd333};
ram[9617] = {-9'd65,10'd336};
ram[9618] = {-9'd62,10'd339};
ram[9619] = {-9'd59,10'd342};
ram[9620] = {-9'd55,10'd345};
ram[9621] = {-9'd52,10'd348};
ram[9622] = {-9'd49,10'd351};
ram[9623] = {-9'd46,10'd354};
ram[9624] = {-9'd43,10'd358};
ram[9625] = {-9'd40,10'd361};
ram[9626] = {-9'd37,10'd364};
ram[9627] = {-9'd33,10'd367};
ram[9628] = {-9'd30,10'd370};
ram[9629] = {-9'd27,10'd373};
ram[9630] = {-9'd24,10'd376};
ram[9631] = {-9'd21,10'd380};
ram[9632] = {-9'd18,10'd383};
ram[9633] = {-9'd15,10'd386};
ram[9634] = {-9'd11,10'd389};
ram[9635] = {-9'd8,10'd392};
ram[9636] = {-9'd5,10'd395};
ram[9637] = {-9'd2,10'd398};
ram[9638] = {9'd1,-10'd399};
ram[9639] = {9'd4,-10'd396};
ram[9640] = {9'd7,-10'd393};
ram[9641] = {9'd10,-10'd390};
ram[9642] = {9'd14,-10'd387};
ram[9643] = {9'd17,-10'd384};
ram[9644] = {9'd20,-10'd381};
ram[9645] = {9'd23,-10'd377};
ram[9646] = {9'd26,-10'd374};
ram[9647] = {9'd29,-10'd371};
ram[9648] = {9'd32,-10'd368};
ram[9649] = {9'd36,-10'd365};
ram[9650] = {9'd39,-10'd362};
ram[9651] = {9'd42,-10'd359};
ram[9652] = {9'd45,-10'd355};
ram[9653] = {9'd48,-10'd352};
ram[9654] = {9'd51,-10'd349};
ram[9655] = {9'd54,-10'd346};
ram[9656] = {9'd58,-10'd343};
ram[9657] = {9'd61,-10'd340};
ram[9658] = {9'd64,-10'd337};
ram[9659] = {9'd67,-10'd334};
ram[9660] = {9'd70,-10'd330};
ram[9661] = {9'd73,-10'd327};
ram[9662] = {9'd76,-10'd324};
ram[9663] = {9'd80,-10'd321};
ram[9664] = {9'd83,-10'd318};
ram[9665] = {9'd86,-10'd315};
ram[9666] = {9'd89,-10'd312};
ram[9667] = {9'd92,-10'd308};
ram[9668] = {9'd95,-10'd305};
ram[9669] = {9'd98,-10'd302};
ram[9670] = {-9'd99,-10'd299};
ram[9671] = {-9'd96,-10'd296};
ram[9672] = {-9'd92,-10'd293};
ram[9673] = {-9'd89,-10'd290};
ram[9674] = {-9'd86,-10'd286};
ram[9675] = {-9'd83,-10'd283};
ram[9676] = {-9'd80,-10'd280};
ram[9677] = {-9'd77,-10'd277};
ram[9678] = {-9'd74,-10'd274};
ram[9679] = {-9'd70,-10'd271};
ram[9680] = {-9'd67,-10'd268};
ram[9681] = {-9'd64,-10'd264};
ram[9682] = {-9'd61,-10'd261};
ram[9683] = {-9'd58,-10'd258};
ram[9684] = {-9'd55,-10'd255};
ram[9685] = {-9'd52,-10'd252};
ram[9686] = {-9'd48,-10'd249};
ram[9687] = {-9'd45,-10'd246};
ram[9688] = {-9'd42,-10'd242};
ram[9689] = {-9'd39,-10'd239};
ram[9690] = {-9'd36,-10'd236};
ram[9691] = {-9'd33,-10'd233};
ram[9692] = {-9'd30,-10'd230};
ram[9693] = {-9'd26,-10'd227};
ram[9694] = {-9'd23,-10'd224};
ram[9695] = {-9'd20,-10'd220};
ram[9696] = {-9'd17,-10'd217};
ram[9697] = {-9'd14,-10'd214};
ram[9698] = {-9'd11,-10'd211};
ram[9699] = {-9'd8,-10'd208};
ram[9700] = {-9'd4,-10'd205};
ram[9701] = {-9'd1,-10'd202};
ram[9702] = {9'd2,-10'd198};
ram[9703] = {9'd5,-10'd195};
ram[9704] = {9'd8,-10'd192};
ram[9705] = {9'd11,-10'd189};
ram[9706] = {9'd14,-10'd186};
ram[9707] = {9'd18,-10'd183};
ram[9708] = {9'd21,-10'd180};
ram[9709] = {9'd24,-10'd176};
ram[9710] = {9'd27,-10'd173};
ram[9711] = {9'd30,-10'd170};
ram[9712] = {9'd33,-10'd167};
ram[9713] = {9'd36,-10'd164};
ram[9714] = {9'd40,-10'd161};
ram[9715] = {9'd43,-10'd158};
ram[9716] = {9'd46,-10'd154};
ram[9717] = {9'd49,-10'd151};
ram[9718] = {9'd52,-10'd148};
ram[9719] = {9'd55,-10'd145};
ram[9720] = {9'd58,-10'd142};
ram[9721] = {9'd62,-10'd139};
ram[9722] = {9'd65,-10'd136};
ram[9723] = {9'd68,-10'd132};
ram[9724] = {9'd71,-10'd129};
ram[9725] = {9'd74,-10'd126};
ram[9726] = {9'd77,-10'd123};
ram[9727] = {9'd80,-10'd120};
ram[9728] = {9'd80,-10'd120};
ram[9729] = {9'd84,-10'd117};
ram[9730] = {9'd87,-10'd114};
ram[9731] = {9'd90,-10'd110};
ram[9732] = {9'd93,-10'd107};
ram[9733] = {9'd96,-10'd104};
ram[9734] = {9'd99,-10'd101};
ram[9735] = {-9'd98,-10'd98};
ram[9736] = {-9'd95,-10'd95};
ram[9737] = {-9'd92,-10'd92};
ram[9738] = {-9'd88,-10'd88};
ram[9739] = {-9'd85,-10'd85};
ram[9740] = {-9'd82,-10'd82};
ram[9741] = {-9'd79,-10'd79};
ram[9742] = {-9'd76,-10'd76};
ram[9743] = {-9'd73,-10'd73};
ram[9744] = {-9'd70,-10'd70};
ram[9745] = {-9'd66,-10'd66};
ram[9746] = {-9'd63,-10'd63};
ram[9747] = {-9'd60,-10'd60};
ram[9748] = {-9'd57,-10'd57};
ram[9749] = {-9'd54,-10'd54};
ram[9750] = {-9'd51,-10'd51};
ram[9751] = {-9'd48,-10'd48};
ram[9752] = {-9'd44,-10'd44};
ram[9753] = {-9'd41,-10'd41};
ram[9754] = {-9'd38,-10'd38};
ram[9755] = {-9'd35,-10'd35};
ram[9756] = {-9'd32,-10'd32};
ram[9757] = {-9'd29,-10'd29};
ram[9758] = {-9'd26,-10'd26};
ram[9759] = {-9'd22,-10'd22};
ram[9760] = {-9'd19,-10'd19};
ram[9761] = {-9'd16,-10'd16};
ram[9762] = {-9'd13,-10'd13};
ram[9763] = {-9'd10,-10'd10};
ram[9764] = {-9'd7,-10'd7};
ram[9765] = {-9'd4,-10'd4};
ram[9766] = {9'd0,10'd0};
ram[9767] = {9'd3,10'd3};
ram[9768] = {9'd6,10'd6};
ram[9769] = {9'd9,10'd9};
ram[9770] = {9'd12,10'd12};
ram[9771] = {9'd15,10'd15};
ram[9772] = {9'd18,10'd18};
ram[9773] = {9'd21,10'd21};
ram[9774] = {9'd25,10'd25};
ram[9775] = {9'd28,10'd28};
ram[9776] = {9'd31,10'd31};
ram[9777] = {9'd34,10'd34};
ram[9778] = {9'd37,10'd37};
ram[9779] = {9'd40,10'd40};
ram[9780] = {9'd43,10'd43};
ram[9781] = {9'd47,10'd47};
ram[9782] = {9'd50,10'd50};
ram[9783] = {9'd53,10'd53};
ram[9784] = {9'd56,10'd56};
ram[9785] = {9'd59,10'd59};
ram[9786] = {9'd62,10'd62};
ram[9787] = {9'd65,10'd65};
ram[9788] = {9'd69,10'd69};
ram[9789] = {9'd72,10'd72};
ram[9790] = {9'd75,10'd75};
ram[9791] = {9'd78,10'd78};
ram[9792] = {9'd81,10'd81};
ram[9793] = {9'd84,10'd84};
ram[9794] = {9'd87,10'd87};
ram[9795] = {9'd91,10'd91};
ram[9796] = {9'd94,10'd94};
ram[9797] = {9'd97,10'd97};
ram[9798] = {-9'd100,10'd100};
ram[9799] = {-9'd97,10'd103};
ram[9800] = {-9'd94,10'd106};
ram[9801] = {-9'd91,10'd109};
ram[9802] = {-9'd88,10'd113};
ram[9803] = {-9'd85,10'd116};
ram[9804] = {-9'd81,10'd119};
ram[9805] = {-9'd78,10'd122};
ram[9806] = {-9'd75,10'd125};
ram[9807] = {-9'd72,10'd128};
ram[9808] = {-9'd69,10'd131};
ram[9809] = {-9'd66,10'd135};
ram[9810] = {-9'd63,10'd138};
ram[9811] = {-9'd59,10'd141};
ram[9812] = {-9'd56,10'd144};
ram[9813] = {-9'd53,10'd147};
ram[9814] = {-9'd50,10'd150};
ram[9815] = {-9'd47,10'd153};
ram[9816] = {-9'd44,10'd157};
ram[9817] = {-9'd41,10'd160};
ram[9818] = {-9'd37,10'd163};
ram[9819] = {-9'd34,10'd166};
ram[9820] = {-9'd31,10'd169};
ram[9821] = {-9'd28,10'd172};
ram[9822] = {-9'd25,10'd175};
ram[9823] = {-9'd22,10'd179};
ram[9824] = {-9'd19,10'd182};
ram[9825] = {-9'd15,10'd185};
ram[9826] = {-9'd12,10'd188};
ram[9827] = {-9'd9,10'd191};
ram[9828] = {-9'd6,10'd194};
ram[9829] = {-9'd3,10'd197};
ram[9830] = {9'd0,10'd201};
ram[9831] = {9'd3,10'd204};
ram[9832] = {9'd7,10'd207};
ram[9833] = {9'd10,10'd210};
ram[9834] = {9'd13,10'd213};
ram[9835] = {9'd16,10'd216};
ram[9836] = {9'd19,10'd219};
ram[9837] = {9'd22,10'd223};
ram[9838] = {9'd25,10'd226};
ram[9839] = {9'd29,10'd229};
ram[9840] = {9'd32,10'd232};
ram[9841] = {9'd35,10'd235};
ram[9842] = {9'd38,10'd238};
ram[9843] = {9'd41,10'd241};
ram[9844] = {9'd44,10'd245};
ram[9845] = {9'd47,10'd248};
ram[9846] = {9'd51,10'd251};
ram[9847] = {9'd54,10'd254};
ram[9848] = {9'd57,10'd257};
ram[9849] = {9'd60,10'd260};
ram[9850] = {9'd63,10'd263};
ram[9851] = {9'd66,10'd267};
ram[9852] = {9'd69,10'd270};
ram[9853] = {9'd73,10'd273};
ram[9854] = {9'd76,10'd276};
ram[9855] = {9'd79,10'd279};
ram[9856] = {9'd79,10'd279};
ram[9857] = {9'd82,10'd282};
ram[9858] = {9'd85,10'd285};
ram[9859] = {9'd88,10'd289};
ram[9860] = {9'd91,10'd292};
ram[9861] = {9'd95,10'd295};
ram[9862] = {9'd98,10'd298};
ram[9863] = {-9'd99,10'd301};
ram[9864] = {-9'd96,10'd304};
ram[9865] = {-9'd93,10'd307};
ram[9866] = {-9'd90,10'd311};
ram[9867] = {-9'd87,10'd314};
ram[9868] = {-9'd84,10'd317};
ram[9869] = {-9'd81,10'd320};
ram[9870] = {-9'd77,10'd323};
ram[9871] = {-9'd74,10'd326};
ram[9872] = {-9'd71,10'd329};
ram[9873] = {-9'd68,10'd333};
ram[9874] = {-9'd65,10'd336};
ram[9875] = {-9'd62,10'd339};
ram[9876] = {-9'd59,10'd342};
ram[9877] = {-9'd55,10'd345};
ram[9878] = {-9'd52,10'd348};
ram[9879] = {-9'd49,10'd351};
ram[9880] = {-9'd46,10'd354};
ram[9881] = {-9'd43,10'd358};
ram[9882] = {-9'd40,10'd361};
ram[9883] = {-9'd37,10'd364};
ram[9884] = {-9'd33,10'd367};
ram[9885] = {-9'd30,10'd370};
ram[9886] = {-9'd27,10'd373};
ram[9887] = {-9'd24,10'd376};
ram[9888] = {-9'd21,10'd380};
ram[9889] = {-9'd18,10'd383};
ram[9890] = {-9'd15,10'd386};
ram[9891] = {-9'd11,10'd389};
ram[9892] = {-9'd8,10'd392};
ram[9893] = {-9'd5,10'd395};
ram[9894] = {-9'd2,10'd398};
ram[9895] = {9'd1,-10'd399};
ram[9896] = {9'd4,-10'd396};
ram[9897] = {9'd7,-10'd393};
ram[9898] = {9'd10,-10'd390};
ram[9899] = {9'd14,-10'd387};
ram[9900] = {9'd17,-10'd384};
ram[9901] = {9'd20,-10'd381};
ram[9902] = {9'd23,-10'd377};
ram[9903] = {9'd26,-10'd374};
ram[9904] = {9'd29,-10'd371};
ram[9905] = {9'd32,-10'd368};
ram[9906] = {9'd36,-10'd365};
ram[9907] = {9'd39,-10'd362};
ram[9908] = {9'd42,-10'd359};
ram[9909] = {9'd45,-10'd355};
ram[9910] = {9'd48,-10'd352};
ram[9911] = {9'd51,-10'd349};
ram[9912] = {9'd54,-10'd346};
ram[9913] = {9'd58,-10'd343};
ram[9914] = {9'd61,-10'd340};
ram[9915] = {9'd64,-10'd337};
ram[9916] = {9'd67,-10'd334};
ram[9917] = {9'd70,-10'd330};
ram[9918] = {9'd73,-10'd327};
ram[9919] = {9'd76,-10'd324};
ram[9920] = {9'd80,-10'd321};
ram[9921] = {9'd83,-10'd318};
ram[9922] = {9'd86,-10'd315};
ram[9923] = {9'd89,-10'd312};
ram[9924] = {9'd92,-10'd308};
ram[9925] = {9'd95,-10'd305};
ram[9926] = {9'd98,-10'd302};
ram[9927] = {-9'd99,-10'd299};
ram[9928] = {-9'd96,-10'd296};
ram[9929] = {-9'd92,-10'd293};
ram[9930] = {-9'd89,-10'd290};
ram[9931] = {-9'd86,-10'd286};
ram[9932] = {-9'd83,-10'd283};
ram[9933] = {-9'd80,-10'd280};
ram[9934] = {-9'd77,-10'd277};
ram[9935] = {-9'd74,-10'd274};
ram[9936] = {-9'd70,-10'd271};
ram[9937] = {-9'd67,-10'd268};
ram[9938] = {-9'd64,-10'd264};
ram[9939] = {-9'd61,-10'd261};
ram[9940] = {-9'd58,-10'd258};
ram[9941] = {-9'd55,-10'd255};
ram[9942] = {-9'd52,-10'd252};
ram[9943] = {-9'd48,-10'd249};
ram[9944] = {-9'd45,-10'd246};
ram[9945] = {-9'd42,-10'd242};
ram[9946] = {-9'd39,-10'd239};
ram[9947] = {-9'd36,-10'd236};
ram[9948] = {-9'd33,-10'd233};
ram[9949] = {-9'd30,-10'd230};
ram[9950] = {-9'd26,-10'd227};
ram[9951] = {-9'd23,-10'd224};
ram[9952] = {-9'd20,-10'd220};
ram[9953] = {-9'd17,-10'd217};
ram[9954] = {-9'd14,-10'd214};
ram[9955] = {-9'd11,-10'd211};
ram[9956] = {-9'd8,-10'd208};
ram[9957] = {-9'd4,-10'd205};
ram[9958] = {-9'd1,-10'd202};
ram[9959] = {9'd2,-10'd198};
ram[9960] = {9'd5,-10'd195};
ram[9961] = {9'd8,-10'd192};
ram[9962] = {9'd11,-10'd189};
ram[9963] = {9'd14,-10'd186};
ram[9964] = {9'd18,-10'd183};
ram[9965] = {9'd21,-10'd180};
ram[9966] = {9'd24,-10'd176};
ram[9967] = {9'd27,-10'd173};
ram[9968] = {9'd30,-10'd170};
ram[9969] = {9'd33,-10'd167};
ram[9970] = {9'd36,-10'd164};
ram[9971] = {9'd40,-10'd161};
ram[9972] = {9'd43,-10'd158};
ram[9973] = {9'd46,-10'd154};
ram[9974] = {9'd49,-10'd151};
ram[9975] = {9'd52,-10'd148};
ram[9976] = {9'd55,-10'd145};
ram[9977] = {9'd58,-10'd142};
ram[9978] = {9'd62,-10'd139};
ram[9979] = {9'd65,-10'd136};
ram[9980] = {9'd68,-10'd132};
ram[9981] = {9'd71,-10'd129};
ram[9982] = {9'd74,-10'd126};
ram[9983] = {9'd77,-10'd123};
ram[9984] = {9'd77,-10'd123};
ram[9985] = {9'd80,-10'd120};
ram[9986] = {9'd84,-10'd117};
ram[9987] = {9'd87,-10'd114};
ram[9988] = {9'd90,-10'd110};
ram[9989] = {9'd93,-10'd107};
ram[9990] = {9'd96,-10'd104};
ram[9991] = {9'd99,-10'd101};
ram[9992] = {-9'd98,-10'd98};
ram[9993] = {-9'd95,-10'd95};
ram[9994] = {-9'd92,-10'd92};
ram[9995] = {-9'd88,-10'd88};
ram[9996] = {-9'd85,-10'd85};
ram[9997] = {-9'd82,-10'd82};
ram[9998] = {-9'd79,-10'd79};
ram[9999] = {-9'd76,-10'd76};
ram[10000] = {-9'd73,-10'd73};
ram[10001] = {-9'd70,-10'd70};
ram[10002] = {-9'd66,-10'd66};
ram[10003] = {-9'd63,-10'd63};
ram[10004] = {-9'd60,-10'd60};
ram[10005] = {-9'd57,-10'd57};
ram[10006] = {-9'd54,-10'd54};
ram[10007] = {-9'd51,-10'd51};
ram[10008] = {-9'd48,-10'd48};
ram[10009] = {-9'd44,-10'd44};
ram[10010] = {-9'd41,-10'd41};
ram[10011] = {-9'd38,-10'd38};
ram[10012] = {-9'd35,-10'd35};
ram[10013] = {-9'd32,-10'd32};
ram[10014] = {-9'd29,-10'd29};
ram[10015] = {-9'd26,-10'd26};
ram[10016] = {-9'd22,-10'd22};
ram[10017] = {-9'd19,-10'd19};
ram[10018] = {-9'd16,-10'd16};
ram[10019] = {-9'd13,-10'd13};
ram[10020] = {-9'd10,-10'd10};
ram[10021] = {-9'd7,-10'd7};
ram[10022] = {-9'd4,-10'd4};
ram[10023] = {9'd0,10'd0};
ram[10024] = {9'd3,10'd3};
ram[10025] = {9'd6,10'd6};
ram[10026] = {9'd9,10'd9};
ram[10027] = {9'd12,10'd12};
ram[10028] = {9'd15,10'd15};
ram[10029] = {9'd18,10'd18};
ram[10030] = {9'd21,10'd21};
ram[10031] = {9'd25,10'd25};
ram[10032] = {9'd28,10'd28};
ram[10033] = {9'd31,10'd31};
ram[10034] = {9'd34,10'd34};
ram[10035] = {9'd37,10'd37};
ram[10036] = {9'd40,10'd40};
ram[10037] = {9'd43,10'd43};
ram[10038] = {9'd47,10'd47};
ram[10039] = {9'd50,10'd50};
ram[10040] = {9'd53,10'd53};
ram[10041] = {9'd56,10'd56};
ram[10042] = {9'd59,10'd59};
ram[10043] = {9'd62,10'd62};
ram[10044] = {9'd65,10'd65};
ram[10045] = {9'd69,10'd69};
ram[10046] = {9'd72,10'd72};
ram[10047] = {9'd75,10'd75};
ram[10048] = {9'd78,10'd78};
ram[10049] = {9'd81,10'd81};
ram[10050] = {9'd84,10'd84};
ram[10051] = {9'd87,10'd87};
ram[10052] = {9'd91,10'd91};
ram[10053] = {9'd94,10'd94};
ram[10054] = {9'd97,10'd97};
ram[10055] = {-9'd100,10'd100};
ram[10056] = {-9'd97,10'd103};
ram[10057] = {-9'd94,10'd106};
ram[10058] = {-9'd91,10'd109};
ram[10059] = {-9'd88,10'd113};
ram[10060] = {-9'd85,10'd116};
ram[10061] = {-9'd81,10'd119};
ram[10062] = {-9'd78,10'd122};
ram[10063] = {-9'd75,10'd125};
ram[10064] = {-9'd72,10'd128};
ram[10065] = {-9'd69,10'd131};
ram[10066] = {-9'd66,10'd135};
ram[10067] = {-9'd63,10'd138};
ram[10068] = {-9'd59,10'd141};
ram[10069] = {-9'd56,10'd144};
ram[10070] = {-9'd53,10'd147};
ram[10071] = {-9'd50,10'd150};
ram[10072] = {-9'd47,10'd153};
ram[10073] = {-9'd44,10'd157};
ram[10074] = {-9'd41,10'd160};
ram[10075] = {-9'd37,10'd163};
ram[10076] = {-9'd34,10'd166};
ram[10077] = {-9'd31,10'd169};
ram[10078] = {-9'd28,10'd172};
ram[10079] = {-9'd25,10'd175};
ram[10080] = {-9'd22,10'd179};
ram[10081] = {-9'd19,10'd182};
ram[10082] = {-9'd15,10'd185};
ram[10083] = {-9'd12,10'd188};
ram[10084] = {-9'd9,10'd191};
ram[10085] = {-9'd6,10'd194};
ram[10086] = {-9'd3,10'd197};
ram[10087] = {9'd0,10'd201};
ram[10088] = {9'd3,10'd204};
ram[10089] = {9'd7,10'd207};
ram[10090] = {9'd10,10'd210};
ram[10091] = {9'd13,10'd213};
ram[10092] = {9'd16,10'd216};
ram[10093] = {9'd19,10'd219};
ram[10094] = {9'd22,10'd223};
ram[10095] = {9'd25,10'd226};
ram[10096] = {9'd29,10'd229};
ram[10097] = {9'd32,10'd232};
ram[10098] = {9'd35,10'd235};
ram[10099] = {9'd38,10'd238};
ram[10100] = {9'd41,10'd241};
ram[10101] = {9'd44,10'd245};
ram[10102] = {9'd47,10'd248};
ram[10103] = {9'd51,10'd251};
ram[10104] = {9'd54,10'd254};
ram[10105] = {9'd57,10'd257};
ram[10106] = {9'd60,10'd260};
ram[10107] = {9'd63,10'd263};
ram[10108] = {9'd66,10'd267};
ram[10109] = {9'd69,10'd270};
ram[10110] = {9'd73,10'd273};
ram[10111] = {9'd76,10'd276};
ram[10112] = {9'd76,10'd276};
ram[10113] = {9'd79,10'd279};
ram[10114] = {9'd82,10'd282};
ram[10115] = {9'd85,10'd285};
ram[10116] = {9'd88,10'd289};
ram[10117] = {9'd91,10'd292};
ram[10118] = {9'd95,10'd295};
ram[10119] = {9'd98,10'd298};
ram[10120] = {-9'd99,10'd301};
ram[10121] = {-9'd96,10'd304};
ram[10122] = {-9'd93,10'd307};
ram[10123] = {-9'd90,10'd311};
ram[10124] = {-9'd87,10'd314};
ram[10125] = {-9'd84,10'd317};
ram[10126] = {-9'd81,10'd320};
ram[10127] = {-9'd77,10'd323};
ram[10128] = {-9'd74,10'd326};
ram[10129] = {-9'd71,10'd329};
ram[10130] = {-9'd68,10'd333};
ram[10131] = {-9'd65,10'd336};
ram[10132] = {-9'd62,10'd339};
ram[10133] = {-9'd59,10'd342};
ram[10134] = {-9'd55,10'd345};
ram[10135] = {-9'd52,10'd348};
ram[10136] = {-9'd49,10'd351};
ram[10137] = {-9'd46,10'd354};
ram[10138] = {-9'd43,10'd358};
ram[10139] = {-9'd40,10'd361};
ram[10140] = {-9'd37,10'd364};
ram[10141] = {-9'd33,10'd367};
ram[10142] = {-9'd30,10'd370};
ram[10143] = {-9'd27,10'd373};
ram[10144] = {-9'd24,10'd376};
ram[10145] = {-9'd21,10'd380};
ram[10146] = {-9'd18,10'd383};
ram[10147] = {-9'd15,10'd386};
ram[10148] = {-9'd11,10'd389};
ram[10149] = {-9'd8,10'd392};
ram[10150] = {-9'd5,10'd395};
ram[10151] = {-9'd2,10'd398};
ram[10152] = {9'd1,-10'd399};
ram[10153] = {9'd4,-10'd396};
ram[10154] = {9'd7,-10'd393};
ram[10155] = {9'd10,-10'd390};
ram[10156] = {9'd14,-10'd387};
ram[10157] = {9'd17,-10'd384};
ram[10158] = {9'd20,-10'd381};
ram[10159] = {9'd23,-10'd377};
ram[10160] = {9'd26,-10'd374};
ram[10161] = {9'd29,-10'd371};
ram[10162] = {9'd32,-10'd368};
ram[10163] = {9'd36,-10'd365};
ram[10164] = {9'd39,-10'd362};
ram[10165] = {9'd42,-10'd359};
ram[10166] = {9'd45,-10'd355};
ram[10167] = {9'd48,-10'd352};
ram[10168] = {9'd51,-10'd349};
ram[10169] = {9'd54,-10'd346};
ram[10170] = {9'd58,-10'd343};
ram[10171] = {9'd61,-10'd340};
ram[10172] = {9'd64,-10'd337};
ram[10173] = {9'd67,-10'd334};
ram[10174] = {9'd70,-10'd330};
ram[10175] = {9'd73,-10'd327};
ram[10176] = {9'd76,-10'd324};
ram[10177] = {9'd80,-10'd321};
ram[10178] = {9'd83,-10'd318};
ram[10179] = {9'd86,-10'd315};
ram[10180] = {9'd89,-10'd312};
ram[10181] = {9'd92,-10'd308};
ram[10182] = {9'd95,-10'd305};
ram[10183] = {9'd98,-10'd302};
ram[10184] = {-9'd99,-10'd299};
ram[10185] = {-9'd96,-10'd296};
ram[10186] = {-9'd92,-10'd293};
ram[10187] = {-9'd89,-10'd290};
ram[10188] = {-9'd86,-10'd286};
ram[10189] = {-9'd83,-10'd283};
ram[10190] = {-9'd80,-10'd280};
ram[10191] = {-9'd77,-10'd277};
ram[10192] = {-9'd74,-10'd274};
ram[10193] = {-9'd70,-10'd271};
ram[10194] = {-9'd67,-10'd268};
ram[10195] = {-9'd64,-10'd264};
ram[10196] = {-9'd61,-10'd261};
ram[10197] = {-9'd58,-10'd258};
ram[10198] = {-9'd55,-10'd255};
ram[10199] = {-9'd52,-10'd252};
ram[10200] = {-9'd48,-10'd249};
ram[10201] = {-9'd45,-10'd246};
ram[10202] = {-9'd42,-10'd242};
ram[10203] = {-9'd39,-10'd239};
ram[10204] = {-9'd36,-10'd236};
ram[10205] = {-9'd33,-10'd233};
ram[10206] = {-9'd30,-10'd230};
ram[10207] = {-9'd26,-10'd227};
ram[10208] = {-9'd23,-10'd224};
ram[10209] = {-9'd20,-10'd220};
ram[10210] = {-9'd17,-10'd217};
ram[10211] = {-9'd14,-10'd214};
ram[10212] = {-9'd11,-10'd211};
ram[10213] = {-9'd8,-10'd208};
ram[10214] = {-9'd4,-10'd205};
ram[10215] = {-9'd1,-10'd202};
ram[10216] = {9'd2,-10'd198};
ram[10217] = {9'd5,-10'd195};
ram[10218] = {9'd8,-10'd192};
ram[10219] = {9'd11,-10'd189};
ram[10220] = {9'd14,-10'd186};
ram[10221] = {9'd18,-10'd183};
ram[10222] = {9'd21,-10'd180};
ram[10223] = {9'd24,-10'd176};
ram[10224] = {9'd27,-10'd173};
ram[10225] = {9'd30,-10'd170};
ram[10226] = {9'd33,-10'd167};
ram[10227] = {9'd36,-10'd164};
ram[10228] = {9'd40,-10'd161};
ram[10229] = {9'd43,-10'd158};
ram[10230] = {9'd46,-10'd154};
ram[10231] = {9'd49,-10'd151};
ram[10232] = {9'd52,-10'd148};
ram[10233] = {9'd55,-10'd145};
ram[10234] = {9'd58,-10'd142};
ram[10235] = {9'd62,-10'd139};
ram[10236] = {9'd65,-10'd136};
ram[10237] = {9'd68,-10'd132};
ram[10238] = {9'd71,-10'd129};
ram[10239] = {9'd74,-10'd126};
ram[10240] = {9'd74,-10'd126};
ram[10241] = {9'd77,-10'd123};
ram[10242] = {9'd80,-10'd120};
ram[10243] = {9'd84,-10'd117};
ram[10244] = {9'd87,-10'd114};
ram[10245] = {9'd90,-10'd110};
ram[10246] = {9'd93,-10'd107};
ram[10247] = {9'd96,-10'd104};
ram[10248] = {9'd99,-10'd101};
ram[10249] = {-9'd98,-10'd98};
ram[10250] = {-9'd95,-10'd95};
ram[10251] = {-9'd92,-10'd92};
ram[10252] = {-9'd88,-10'd88};
ram[10253] = {-9'd85,-10'd85};
ram[10254] = {-9'd82,-10'd82};
ram[10255] = {-9'd79,-10'd79};
ram[10256] = {-9'd76,-10'd76};
ram[10257] = {-9'd73,-10'd73};
ram[10258] = {-9'd70,-10'd70};
ram[10259] = {-9'd66,-10'd66};
ram[10260] = {-9'd63,-10'd63};
ram[10261] = {-9'd60,-10'd60};
ram[10262] = {-9'd57,-10'd57};
ram[10263] = {-9'd54,-10'd54};
ram[10264] = {-9'd51,-10'd51};
ram[10265] = {-9'd48,-10'd48};
ram[10266] = {-9'd44,-10'd44};
ram[10267] = {-9'd41,-10'd41};
ram[10268] = {-9'd38,-10'd38};
ram[10269] = {-9'd35,-10'd35};
ram[10270] = {-9'd32,-10'd32};
ram[10271] = {-9'd29,-10'd29};
ram[10272] = {-9'd26,-10'd26};
ram[10273] = {-9'd22,-10'd22};
ram[10274] = {-9'd19,-10'd19};
ram[10275] = {-9'd16,-10'd16};
ram[10276] = {-9'd13,-10'd13};
ram[10277] = {-9'd10,-10'd10};
ram[10278] = {-9'd7,-10'd7};
ram[10279] = {-9'd4,-10'd4};
ram[10280] = {9'd0,10'd0};
ram[10281] = {9'd3,10'd3};
ram[10282] = {9'd6,10'd6};
ram[10283] = {9'd9,10'd9};
ram[10284] = {9'd12,10'd12};
ram[10285] = {9'd15,10'd15};
ram[10286] = {9'd18,10'd18};
ram[10287] = {9'd21,10'd21};
ram[10288] = {9'd25,10'd25};
ram[10289] = {9'd28,10'd28};
ram[10290] = {9'd31,10'd31};
ram[10291] = {9'd34,10'd34};
ram[10292] = {9'd37,10'd37};
ram[10293] = {9'd40,10'd40};
ram[10294] = {9'd43,10'd43};
ram[10295] = {9'd47,10'd47};
ram[10296] = {9'd50,10'd50};
ram[10297] = {9'd53,10'd53};
ram[10298] = {9'd56,10'd56};
ram[10299] = {9'd59,10'd59};
ram[10300] = {9'd62,10'd62};
ram[10301] = {9'd65,10'd65};
ram[10302] = {9'd69,10'd69};
ram[10303] = {9'd72,10'd72};
ram[10304] = {9'd75,10'd75};
ram[10305] = {9'd78,10'd78};
ram[10306] = {9'd81,10'd81};
ram[10307] = {9'd84,10'd84};
ram[10308] = {9'd87,10'd87};
ram[10309] = {9'd91,10'd91};
ram[10310] = {9'd94,10'd94};
ram[10311] = {9'd97,10'd97};
ram[10312] = {-9'd100,10'd100};
ram[10313] = {-9'd97,10'd103};
ram[10314] = {-9'd94,10'd106};
ram[10315] = {-9'd91,10'd109};
ram[10316] = {-9'd88,10'd113};
ram[10317] = {-9'd85,10'd116};
ram[10318] = {-9'd81,10'd119};
ram[10319] = {-9'd78,10'd122};
ram[10320] = {-9'd75,10'd125};
ram[10321] = {-9'd72,10'd128};
ram[10322] = {-9'd69,10'd131};
ram[10323] = {-9'd66,10'd135};
ram[10324] = {-9'd63,10'd138};
ram[10325] = {-9'd59,10'd141};
ram[10326] = {-9'd56,10'd144};
ram[10327] = {-9'd53,10'd147};
ram[10328] = {-9'd50,10'd150};
ram[10329] = {-9'd47,10'd153};
ram[10330] = {-9'd44,10'd157};
ram[10331] = {-9'd41,10'd160};
ram[10332] = {-9'd37,10'd163};
ram[10333] = {-9'd34,10'd166};
ram[10334] = {-9'd31,10'd169};
ram[10335] = {-9'd28,10'd172};
ram[10336] = {-9'd25,10'd175};
ram[10337] = {-9'd22,10'd179};
ram[10338] = {-9'd19,10'd182};
ram[10339] = {-9'd15,10'd185};
ram[10340] = {-9'd12,10'd188};
ram[10341] = {-9'd9,10'd191};
ram[10342] = {-9'd6,10'd194};
ram[10343] = {-9'd3,10'd197};
ram[10344] = {9'd0,10'd201};
ram[10345] = {9'd3,10'd204};
ram[10346] = {9'd7,10'd207};
ram[10347] = {9'd10,10'd210};
ram[10348] = {9'd13,10'd213};
ram[10349] = {9'd16,10'd216};
ram[10350] = {9'd19,10'd219};
ram[10351] = {9'd22,10'd223};
ram[10352] = {9'd25,10'd226};
ram[10353] = {9'd29,10'd229};
ram[10354] = {9'd32,10'd232};
ram[10355] = {9'd35,10'd235};
ram[10356] = {9'd38,10'd238};
ram[10357] = {9'd41,10'd241};
ram[10358] = {9'd44,10'd245};
ram[10359] = {9'd47,10'd248};
ram[10360] = {9'd51,10'd251};
ram[10361] = {9'd54,10'd254};
ram[10362] = {9'd57,10'd257};
ram[10363] = {9'd60,10'd260};
ram[10364] = {9'd63,10'd263};
ram[10365] = {9'd66,10'd267};
ram[10366] = {9'd69,10'd270};
ram[10367] = {9'd73,10'd273};
ram[10368] = {9'd73,10'd273};
ram[10369] = {9'd76,10'd276};
ram[10370] = {9'd79,10'd279};
ram[10371] = {9'd82,10'd282};
ram[10372] = {9'd85,10'd285};
ram[10373] = {9'd88,10'd289};
ram[10374] = {9'd91,10'd292};
ram[10375] = {9'd95,10'd295};
ram[10376] = {9'd98,10'd298};
ram[10377] = {-9'd99,10'd301};
ram[10378] = {-9'd96,10'd304};
ram[10379] = {-9'd93,10'd307};
ram[10380] = {-9'd90,10'd311};
ram[10381] = {-9'd87,10'd314};
ram[10382] = {-9'd84,10'd317};
ram[10383] = {-9'd81,10'd320};
ram[10384] = {-9'd77,10'd323};
ram[10385] = {-9'd74,10'd326};
ram[10386] = {-9'd71,10'd329};
ram[10387] = {-9'd68,10'd333};
ram[10388] = {-9'd65,10'd336};
ram[10389] = {-9'd62,10'd339};
ram[10390] = {-9'd59,10'd342};
ram[10391] = {-9'd55,10'd345};
ram[10392] = {-9'd52,10'd348};
ram[10393] = {-9'd49,10'd351};
ram[10394] = {-9'd46,10'd354};
ram[10395] = {-9'd43,10'd358};
ram[10396] = {-9'd40,10'd361};
ram[10397] = {-9'd37,10'd364};
ram[10398] = {-9'd33,10'd367};
ram[10399] = {-9'd30,10'd370};
ram[10400] = {-9'd27,10'd373};
ram[10401] = {-9'd24,10'd376};
ram[10402] = {-9'd21,10'd380};
ram[10403] = {-9'd18,10'd383};
ram[10404] = {-9'd15,10'd386};
ram[10405] = {-9'd11,10'd389};
ram[10406] = {-9'd8,10'd392};
ram[10407] = {-9'd5,10'd395};
ram[10408] = {-9'd2,10'd398};
ram[10409] = {9'd1,-10'd399};
ram[10410] = {9'd4,-10'd396};
ram[10411] = {9'd7,-10'd393};
ram[10412] = {9'd10,-10'd390};
ram[10413] = {9'd14,-10'd387};
ram[10414] = {9'd17,-10'd384};
ram[10415] = {9'd20,-10'd381};
ram[10416] = {9'd23,-10'd377};
ram[10417] = {9'd26,-10'd374};
ram[10418] = {9'd29,-10'd371};
ram[10419] = {9'd32,-10'd368};
ram[10420] = {9'd36,-10'd365};
ram[10421] = {9'd39,-10'd362};
ram[10422] = {9'd42,-10'd359};
ram[10423] = {9'd45,-10'd355};
ram[10424] = {9'd48,-10'd352};
ram[10425] = {9'd51,-10'd349};
ram[10426] = {9'd54,-10'd346};
ram[10427] = {9'd58,-10'd343};
ram[10428] = {9'd61,-10'd340};
ram[10429] = {9'd64,-10'd337};
ram[10430] = {9'd67,-10'd334};
ram[10431] = {9'd70,-10'd330};
ram[10432] = {9'd73,-10'd327};
ram[10433] = {9'd76,-10'd324};
ram[10434] = {9'd80,-10'd321};
ram[10435] = {9'd83,-10'd318};
ram[10436] = {9'd86,-10'd315};
ram[10437] = {9'd89,-10'd312};
ram[10438] = {9'd92,-10'd308};
ram[10439] = {9'd95,-10'd305};
ram[10440] = {9'd98,-10'd302};
ram[10441] = {-9'd99,-10'd299};
ram[10442] = {-9'd96,-10'd296};
ram[10443] = {-9'd92,-10'd293};
ram[10444] = {-9'd89,-10'd290};
ram[10445] = {-9'd86,-10'd286};
ram[10446] = {-9'd83,-10'd283};
ram[10447] = {-9'd80,-10'd280};
ram[10448] = {-9'd77,-10'd277};
ram[10449] = {-9'd74,-10'd274};
ram[10450] = {-9'd70,-10'd271};
ram[10451] = {-9'd67,-10'd268};
ram[10452] = {-9'd64,-10'd264};
ram[10453] = {-9'd61,-10'd261};
ram[10454] = {-9'd58,-10'd258};
ram[10455] = {-9'd55,-10'd255};
ram[10456] = {-9'd52,-10'd252};
ram[10457] = {-9'd48,-10'd249};
ram[10458] = {-9'd45,-10'd246};
ram[10459] = {-9'd42,-10'd242};
ram[10460] = {-9'd39,-10'd239};
ram[10461] = {-9'd36,-10'd236};
ram[10462] = {-9'd33,-10'd233};
ram[10463] = {-9'd30,-10'd230};
ram[10464] = {-9'd26,-10'd227};
ram[10465] = {-9'd23,-10'd224};
ram[10466] = {-9'd20,-10'd220};
ram[10467] = {-9'd17,-10'd217};
ram[10468] = {-9'd14,-10'd214};
ram[10469] = {-9'd11,-10'd211};
ram[10470] = {-9'd8,-10'd208};
ram[10471] = {-9'd4,-10'd205};
ram[10472] = {-9'd1,-10'd202};
ram[10473] = {9'd2,-10'd198};
ram[10474] = {9'd5,-10'd195};
ram[10475] = {9'd8,-10'd192};
ram[10476] = {9'd11,-10'd189};
ram[10477] = {9'd14,-10'd186};
ram[10478] = {9'd18,-10'd183};
ram[10479] = {9'd21,-10'd180};
ram[10480] = {9'd24,-10'd176};
ram[10481] = {9'd27,-10'd173};
ram[10482] = {9'd30,-10'd170};
ram[10483] = {9'd33,-10'd167};
ram[10484] = {9'd36,-10'd164};
ram[10485] = {9'd40,-10'd161};
ram[10486] = {9'd43,-10'd158};
ram[10487] = {9'd46,-10'd154};
ram[10488] = {9'd49,-10'd151};
ram[10489] = {9'd52,-10'd148};
ram[10490] = {9'd55,-10'd145};
ram[10491] = {9'd58,-10'd142};
ram[10492] = {9'd62,-10'd139};
ram[10493] = {9'd65,-10'd136};
ram[10494] = {9'd68,-10'd132};
ram[10495] = {9'd71,-10'd129};
ram[10496] = {9'd71,-10'd129};
ram[10497] = {9'd74,-10'd126};
ram[10498] = {9'd77,-10'd123};
ram[10499] = {9'd80,-10'd120};
ram[10500] = {9'd84,-10'd117};
ram[10501] = {9'd87,-10'd114};
ram[10502] = {9'd90,-10'd110};
ram[10503] = {9'd93,-10'd107};
ram[10504] = {9'd96,-10'd104};
ram[10505] = {9'd99,-10'd101};
ram[10506] = {-9'd98,-10'd98};
ram[10507] = {-9'd95,-10'd95};
ram[10508] = {-9'd92,-10'd92};
ram[10509] = {-9'd88,-10'd88};
ram[10510] = {-9'd85,-10'd85};
ram[10511] = {-9'd82,-10'd82};
ram[10512] = {-9'd79,-10'd79};
ram[10513] = {-9'd76,-10'd76};
ram[10514] = {-9'd73,-10'd73};
ram[10515] = {-9'd70,-10'd70};
ram[10516] = {-9'd66,-10'd66};
ram[10517] = {-9'd63,-10'd63};
ram[10518] = {-9'd60,-10'd60};
ram[10519] = {-9'd57,-10'd57};
ram[10520] = {-9'd54,-10'd54};
ram[10521] = {-9'd51,-10'd51};
ram[10522] = {-9'd48,-10'd48};
ram[10523] = {-9'd44,-10'd44};
ram[10524] = {-9'd41,-10'd41};
ram[10525] = {-9'd38,-10'd38};
ram[10526] = {-9'd35,-10'd35};
ram[10527] = {-9'd32,-10'd32};
ram[10528] = {-9'd29,-10'd29};
ram[10529] = {-9'd26,-10'd26};
ram[10530] = {-9'd22,-10'd22};
ram[10531] = {-9'd19,-10'd19};
ram[10532] = {-9'd16,-10'd16};
ram[10533] = {-9'd13,-10'd13};
ram[10534] = {-9'd10,-10'd10};
ram[10535] = {-9'd7,-10'd7};
ram[10536] = {-9'd4,-10'd4};
ram[10537] = {9'd0,10'd0};
ram[10538] = {9'd3,10'd3};
ram[10539] = {9'd6,10'd6};
ram[10540] = {9'd9,10'd9};
ram[10541] = {9'd12,10'd12};
ram[10542] = {9'd15,10'd15};
ram[10543] = {9'd18,10'd18};
ram[10544] = {9'd21,10'd21};
ram[10545] = {9'd25,10'd25};
ram[10546] = {9'd28,10'd28};
ram[10547] = {9'd31,10'd31};
ram[10548] = {9'd34,10'd34};
ram[10549] = {9'd37,10'd37};
ram[10550] = {9'd40,10'd40};
ram[10551] = {9'd43,10'd43};
ram[10552] = {9'd47,10'd47};
ram[10553] = {9'd50,10'd50};
ram[10554] = {9'd53,10'd53};
ram[10555] = {9'd56,10'd56};
ram[10556] = {9'd59,10'd59};
ram[10557] = {9'd62,10'd62};
ram[10558] = {9'd65,10'd65};
ram[10559] = {9'd69,10'd69};
ram[10560] = {9'd72,10'd72};
ram[10561] = {9'd75,10'd75};
ram[10562] = {9'd78,10'd78};
ram[10563] = {9'd81,10'd81};
ram[10564] = {9'd84,10'd84};
ram[10565] = {9'd87,10'd87};
ram[10566] = {9'd91,10'd91};
ram[10567] = {9'd94,10'd94};
ram[10568] = {9'd97,10'd97};
ram[10569] = {-9'd100,10'd100};
ram[10570] = {-9'd97,10'd103};
ram[10571] = {-9'd94,10'd106};
ram[10572] = {-9'd91,10'd109};
ram[10573] = {-9'd88,10'd113};
ram[10574] = {-9'd85,10'd116};
ram[10575] = {-9'd81,10'd119};
ram[10576] = {-9'd78,10'd122};
ram[10577] = {-9'd75,10'd125};
ram[10578] = {-9'd72,10'd128};
ram[10579] = {-9'd69,10'd131};
ram[10580] = {-9'd66,10'd135};
ram[10581] = {-9'd63,10'd138};
ram[10582] = {-9'd59,10'd141};
ram[10583] = {-9'd56,10'd144};
ram[10584] = {-9'd53,10'd147};
ram[10585] = {-9'd50,10'd150};
ram[10586] = {-9'd47,10'd153};
ram[10587] = {-9'd44,10'd157};
ram[10588] = {-9'd41,10'd160};
ram[10589] = {-9'd37,10'd163};
ram[10590] = {-9'd34,10'd166};
ram[10591] = {-9'd31,10'd169};
ram[10592] = {-9'd28,10'd172};
ram[10593] = {-9'd25,10'd175};
ram[10594] = {-9'd22,10'd179};
ram[10595] = {-9'd19,10'd182};
ram[10596] = {-9'd15,10'd185};
ram[10597] = {-9'd12,10'd188};
ram[10598] = {-9'd9,10'd191};
ram[10599] = {-9'd6,10'd194};
ram[10600] = {-9'd3,10'd197};
ram[10601] = {9'd0,10'd201};
ram[10602] = {9'd3,10'd204};
ram[10603] = {9'd7,10'd207};
ram[10604] = {9'd10,10'd210};
ram[10605] = {9'd13,10'd213};
ram[10606] = {9'd16,10'd216};
ram[10607] = {9'd19,10'd219};
ram[10608] = {9'd22,10'd223};
ram[10609] = {9'd25,10'd226};
ram[10610] = {9'd29,10'd229};
ram[10611] = {9'd32,10'd232};
ram[10612] = {9'd35,10'd235};
ram[10613] = {9'd38,10'd238};
ram[10614] = {9'd41,10'd241};
ram[10615] = {9'd44,10'd245};
ram[10616] = {9'd47,10'd248};
ram[10617] = {9'd51,10'd251};
ram[10618] = {9'd54,10'd254};
ram[10619] = {9'd57,10'd257};
ram[10620] = {9'd60,10'd260};
ram[10621] = {9'd63,10'd263};
ram[10622] = {9'd66,10'd267};
ram[10623] = {9'd69,10'd270};
ram[10624] = {9'd69,10'd270};
ram[10625] = {9'd73,10'd273};
ram[10626] = {9'd76,10'd276};
ram[10627] = {9'd79,10'd279};
ram[10628] = {9'd82,10'd282};
ram[10629] = {9'd85,10'd285};
ram[10630] = {9'd88,10'd289};
ram[10631] = {9'd91,10'd292};
ram[10632] = {9'd95,10'd295};
ram[10633] = {9'd98,10'd298};
ram[10634] = {-9'd99,10'd301};
ram[10635] = {-9'd96,10'd304};
ram[10636] = {-9'd93,10'd307};
ram[10637] = {-9'd90,10'd311};
ram[10638] = {-9'd87,10'd314};
ram[10639] = {-9'd84,10'd317};
ram[10640] = {-9'd81,10'd320};
ram[10641] = {-9'd77,10'd323};
ram[10642] = {-9'd74,10'd326};
ram[10643] = {-9'd71,10'd329};
ram[10644] = {-9'd68,10'd333};
ram[10645] = {-9'd65,10'd336};
ram[10646] = {-9'd62,10'd339};
ram[10647] = {-9'd59,10'd342};
ram[10648] = {-9'd55,10'd345};
ram[10649] = {-9'd52,10'd348};
ram[10650] = {-9'd49,10'd351};
ram[10651] = {-9'd46,10'd354};
ram[10652] = {-9'd43,10'd358};
ram[10653] = {-9'd40,10'd361};
ram[10654] = {-9'd37,10'd364};
ram[10655] = {-9'd33,10'd367};
ram[10656] = {-9'd30,10'd370};
ram[10657] = {-9'd27,10'd373};
ram[10658] = {-9'd24,10'd376};
ram[10659] = {-9'd21,10'd380};
ram[10660] = {-9'd18,10'd383};
ram[10661] = {-9'd15,10'd386};
ram[10662] = {-9'd11,10'd389};
ram[10663] = {-9'd8,10'd392};
ram[10664] = {-9'd5,10'd395};
ram[10665] = {-9'd2,10'd398};
ram[10666] = {9'd1,-10'd399};
ram[10667] = {9'd4,-10'd396};
ram[10668] = {9'd7,-10'd393};
ram[10669] = {9'd10,-10'd390};
ram[10670] = {9'd14,-10'd387};
ram[10671] = {9'd17,-10'd384};
ram[10672] = {9'd20,-10'd381};
ram[10673] = {9'd23,-10'd377};
ram[10674] = {9'd26,-10'd374};
ram[10675] = {9'd29,-10'd371};
ram[10676] = {9'd32,-10'd368};
ram[10677] = {9'd36,-10'd365};
ram[10678] = {9'd39,-10'd362};
ram[10679] = {9'd42,-10'd359};
ram[10680] = {9'd45,-10'd355};
ram[10681] = {9'd48,-10'd352};
ram[10682] = {9'd51,-10'd349};
ram[10683] = {9'd54,-10'd346};
ram[10684] = {9'd58,-10'd343};
ram[10685] = {9'd61,-10'd340};
ram[10686] = {9'd64,-10'd337};
ram[10687] = {9'd67,-10'd334};
ram[10688] = {9'd70,-10'd330};
ram[10689] = {9'd73,-10'd327};
ram[10690] = {9'd76,-10'd324};
ram[10691] = {9'd80,-10'd321};
ram[10692] = {9'd83,-10'd318};
ram[10693] = {9'd86,-10'd315};
ram[10694] = {9'd89,-10'd312};
ram[10695] = {9'd92,-10'd308};
ram[10696] = {9'd95,-10'd305};
ram[10697] = {9'd98,-10'd302};
ram[10698] = {-9'd99,-10'd299};
ram[10699] = {-9'd96,-10'd296};
ram[10700] = {-9'd92,-10'd293};
ram[10701] = {-9'd89,-10'd290};
ram[10702] = {-9'd86,-10'd286};
ram[10703] = {-9'd83,-10'd283};
ram[10704] = {-9'd80,-10'd280};
ram[10705] = {-9'd77,-10'd277};
ram[10706] = {-9'd74,-10'd274};
ram[10707] = {-9'd70,-10'd271};
ram[10708] = {-9'd67,-10'd268};
ram[10709] = {-9'd64,-10'd264};
ram[10710] = {-9'd61,-10'd261};
ram[10711] = {-9'd58,-10'd258};
ram[10712] = {-9'd55,-10'd255};
ram[10713] = {-9'd52,-10'd252};
ram[10714] = {-9'd48,-10'd249};
ram[10715] = {-9'd45,-10'd246};
ram[10716] = {-9'd42,-10'd242};
ram[10717] = {-9'd39,-10'd239};
ram[10718] = {-9'd36,-10'd236};
ram[10719] = {-9'd33,-10'd233};
ram[10720] = {-9'd30,-10'd230};
ram[10721] = {-9'd26,-10'd227};
ram[10722] = {-9'd23,-10'd224};
ram[10723] = {-9'd20,-10'd220};
ram[10724] = {-9'd17,-10'd217};
ram[10725] = {-9'd14,-10'd214};
ram[10726] = {-9'd11,-10'd211};
ram[10727] = {-9'd8,-10'd208};
ram[10728] = {-9'd4,-10'd205};
ram[10729] = {-9'd1,-10'd202};
ram[10730] = {9'd2,-10'd198};
ram[10731] = {9'd5,-10'd195};
ram[10732] = {9'd8,-10'd192};
ram[10733] = {9'd11,-10'd189};
ram[10734] = {9'd14,-10'd186};
ram[10735] = {9'd18,-10'd183};
ram[10736] = {9'd21,-10'd180};
ram[10737] = {9'd24,-10'd176};
ram[10738] = {9'd27,-10'd173};
ram[10739] = {9'd30,-10'd170};
ram[10740] = {9'd33,-10'd167};
ram[10741] = {9'd36,-10'd164};
ram[10742] = {9'd40,-10'd161};
ram[10743] = {9'd43,-10'd158};
ram[10744] = {9'd46,-10'd154};
ram[10745] = {9'd49,-10'd151};
ram[10746] = {9'd52,-10'd148};
ram[10747] = {9'd55,-10'd145};
ram[10748] = {9'd58,-10'd142};
ram[10749] = {9'd62,-10'd139};
ram[10750] = {9'd65,-10'd136};
ram[10751] = {9'd68,-10'd132};
ram[10752] = {9'd68,-10'd132};
ram[10753] = {9'd71,-10'd129};
ram[10754] = {9'd74,-10'd126};
ram[10755] = {9'd77,-10'd123};
ram[10756] = {9'd80,-10'd120};
ram[10757] = {9'd84,-10'd117};
ram[10758] = {9'd87,-10'd114};
ram[10759] = {9'd90,-10'd110};
ram[10760] = {9'd93,-10'd107};
ram[10761] = {9'd96,-10'd104};
ram[10762] = {9'd99,-10'd101};
ram[10763] = {-9'd98,-10'd98};
ram[10764] = {-9'd95,-10'd95};
ram[10765] = {-9'd92,-10'd92};
ram[10766] = {-9'd88,-10'd88};
ram[10767] = {-9'd85,-10'd85};
ram[10768] = {-9'd82,-10'd82};
ram[10769] = {-9'd79,-10'd79};
ram[10770] = {-9'd76,-10'd76};
ram[10771] = {-9'd73,-10'd73};
ram[10772] = {-9'd70,-10'd70};
ram[10773] = {-9'd66,-10'd66};
ram[10774] = {-9'd63,-10'd63};
ram[10775] = {-9'd60,-10'd60};
ram[10776] = {-9'd57,-10'd57};
ram[10777] = {-9'd54,-10'd54};
ram[10778] = {-9'd51,-10'd51};
ram[10779] = {-9'd48,-10'd48};
ram[10780] = {-9'd44,-10'd44};
ram[10781] = {-9'd41,-10'd41};
ram[10782] = {-9'd38,-10'd38};
ram[10783] = {-9'd35,-10'd35};
ram[10784] = {-9'd32,-10'd32};
ram[10785] = {-9'd29,-10'd29};
ram[10786] = {-9'd26,-10'd26};
ram[10787] = {-9'd22,-10'd22};
ram[10788] = {-9'd19,-10'd19};
ram[10789] = {-9'd16,-10'd16};
ram[10790] = {-9'd13,-10'd13};
ram[10791] = {-9'd10,-10'd10};
ram[10792] = {-9'd7,-10'd7};
ram[10793] = {-9'd4,-10'd4};
ram[10794] = {9'd0,10'd0};
ram[10795] = {9'd3,10'd3};
ram[10796] = {9'd6,10'd6};
ram[10797] = {9'd9,10'd9};
ram[10798] = {9'd12,10'd12};
ram[10799] = {9'd15,10'd15};
ram[10800] = {9'd18,10'd18};
ram[10801] = {9'd21,10'd21};
ram[10802] = {9'd25,10'd25};
ram[10803] = {9'd28,10'd28};
ram[10804] = {9'd31,10'd31};
ram[10805] = {9'd34,10'd34};
ram[10806] = {9'd37,10'd37};
ram[10807] = {9'd40,10'd40};
ram[10808] = {9'd43,10'd43};
ram[10809] = {9'd47,10'd47};
ram[10810] = {9'd50,10'd50};
ram[10811] = {9'd53,10'd53};
ram[10812] = {9'd56,10'd56};
ram[10813] = {9'd59,10'd59};
ram[10814] = {9'd62,10'd62};
ram[10815] = {9'd65,10'd65};
ram[10816] = {9'd69,10'd69};
ram[10817] = {9'd72,10'd72};
ram[10818] = {9'd75,10'd75};
ram[10819] = {9'd78,10'd78};
ram[10820] = {9'd81,10'd81};
ram[10821] = {9'd84,10'd84};
ram[10822] = {9'd87,10'd87};
ram[10823] = {9'd91,10'd91};
ram[10824] = {9'd94,10'd94};
ram[10825] = {9'd97,10'd97};
ram[10826] = {-9'd100,10'd100};
ram[10827] = {-9'd97,10'd103};
ram[10828] = {-9'd94,10'd106};
ram[10829] = {-9'd91,10'd109};
ram[10830] = {-9'd88,10'd113};
ram[10831] = {-9'd85,10'd116};
ram[10832] = {-9'd81,10'd119};
ram[10833] = {-9'd78,10'd122};
ram[10834] = {-9'd75,10'd125};
ram[10835] = {-9'd72,10'd128};
ram[10836] = {-9'd69,10'd131};
ram[10837] = {-9'd66,10'd135};
ram[10838] = {-9'd63,10'd138};
ram[10839] = {-9'd59,10'd141};
ram[10840] = {-9'd56,10'd144};
ram[10841] = {-9'd53,10'd147};
ram[10842] = {-9'd50,10'd150};
ram[10843] = {-9'd47,10'd153};
ram[10844] = {-9'd44,10'd157};
ram[10845] = {-9'd41,10'd160};
ram[10846] = {-9'd37,10'd163};
ram[10847] = {-9'd34,10'd166};
ram[10848] = {-9'd31,10'd169};
ram[10849] = {-9'd28,10'd172};
ram[10850] = {-9'd25,10'd175};
ram[10851] = {-9'd22,10'd179};
ram[10852] = {-9'd19,10'd182};
ram[10853] = {-9'd15,10'd185};
ram[10854] = {-9'd12,10'd188};
ram[10855] = {-9'd9,10'd191};
ram[10856] = {-9'd6,10'd194};
ram[10857] = {-9'd3,10'd197};
ram[10858] = {9'd0,10'd201};
ram[10859] = {9'd3,10'd204};
ram[10860] = {9'd7,10'd207};
ram[10861] = {9'd10,10'd210};
ram[10862] = {9'd13,10'd213};
ram[10863] = {9'd16,10'd216};
ram[10864] = {9'd19,10'd219};
ram[10865] = {9'd22,10'd223};
ram[10866] = {9'd25,10'd226};
ram[10867] = {9'd29,10'd229};
ram[10868] = {9'd32,10'd232};
ram[10869] = {9'd35,10'd235};
ram[10870] = {9'd38,10'd238};
ram[10871] = {9'd41,10'd241};
ram[10872] = {9'd44,10'd245};
ram[10873] = {9'd47,10'd248};
ram[10874] = {9'd51,10'd251};
ram[10875] = {9'd54,10'd254};
ram[10876] = {9'd57,10'd257};
ram[10877] = {9'd60,10'd260};
ram[10878] = {9'd63,10'd263};
ram[10879] = {9'd66,10'd267};
ram[10880] = {9'd66,10'd267};
ram[10881] = {9'd69,10'd270};
ram[10882] = {9'd73,10'd273};
ram[10883] = {9'd76,10'd276};
ram[10884] = {9'd79,10'd279};
ram[10885] = {9'd82,10'd282};
ram[10886] = {9'd85,10'd285};
ram[10887] = {9'd88,10'd289};
ram[10888] = {9'd91,10'd292};
ram[10889] = {9'd95,10'd295};
ram[10890] = {9'd98,10'd298};
ram[10891] = {-9'd99,10'd301};
ram[10892] = {-9'd96,10'd304};
ram[10893] = {-9'd93,10'd307};
ram[10894] = {-9'd90,10'd311};
ram[10895] = {-9'd87,10'd314};
ram[10896] = {-9'd84,10'd317};
ram[10897] = {-9'd81,10'd320};
ram[10898] = {-9'd77,10'd323};
ram[10899] = {-9'd74,10'd326};
ram[10900] = {-9'd71,10'd329};
ram[10901] = {-9'd68,10'd333};
ram[10902] = {-9'd65,10'd336};
ram[10903] = {-9'd62,10'd339};
ram[10904] = {-9'd59,10'd342};
ram[10905] = {-9'd55,10'd345};
ram[10906] = {-9'd52,10'd348};
ram[10907] = {-9'd49,10'd351};
ram[10908] = {-9'd46,10'd354};
ram[10909] = {-9'd43,10'd358};
ram[10910] = {-9'd40,10'd361};
ram[10911] = {-9'd37,10'd364};
ram[10912] = {-9'd33,10'd367};
ram[10913] = {-9'd30,10'd370};
ram[10914] = {-9'd27,10'd373};
ram[10915] = {-9'd24,10'd376};
ram[10916] = {-9'd21,10'd380};
ram[10917] = {-9'd18,10'd383};
ram[10918] = {-9'd15,10'd386};
ram[10919] = {-9'd11,10'd389};
ram[10920] = {-9'd8,10'd392};
ram[10921] = {-9'd5,10'd395};
ram[10922] = {-9'd2,10'd398};
ram[10923] = {9'd1,-10'd399};
ram[10924] = {9'd4,-10'd396};
ram[10925] = {9'd7,-10'd393};
ram[10926] = {9'd10,-10'd390};
ram[10927] = {9'd14,-10'd387};
ram[10928] = {9'd17,-10'd384};
ram[10929] = {9'd20,-10'd381};
ram[10930] = {9'd23,-10'd377};
ram[10931] = {9'd26,-10'd374};
ram[10932] = {9'd29,-10'd371};
ram[10933] = {9'd32,-10'd368};
ram[10934] = {9'd36,-10'd365};
ram[10935] = {9'd39,-10'd362};
ram[10936] = {9'd42,-10'd359};
ram[10937] = {9'd45,-10'd355};
ram[10938] = {9'd48,-10'd352};
ram[10939] = {9'd51,-10'd349};
ram[10940] = {9'd54,-10'd346};
ram[10941] = {9'd58,-10'd343};
ram[10942] = {9'd61,-10'd340};
ram[10943] = {9'd64,-10'd337};
ram[10944] = {9'd67,-10'd334};
ram[10945] = {9'd70,-10'd330};
ram[10946] = {9'd73,-10'd327};
ram[10947] = {9'd76,-10'd324};
ram[10948] = {9'd80,-10'd321};
ram[10949] = {9'd83,-10'd318};
ram[10950] = {9'd86,-10'd315};
ram[10951] = {9'd89,-10'd312};
ram[10952] = {9'd92,-10'd308};
ram[10953] = {9'd95,-10'd305};
ram[10954] = {9'd98,-10'd302};
ram[10955] = {-9'd99,-10'd299};
ram[10956] = {-9'd96,-10'd296};
ram[10957] = {-9'd92,-10'd293};
ram[10958] = {-9'd89,-10'd290};
ram[10959] = {-9'd86,-10'd286};
ram[10960] = {-9'd83,-10'd283};
ram[10961] = {-9'd80,-10'd280};
ram[10962] = {-9'd77,-10'd277};
ram[10963] = {-9'd74,-10'd274};
ram[10964] = {-9'd70,-10'd271};
ram[10965] = {-9'd67,-10'd268};
ram[10966] = {-9'd64,-10'd264};
ram[10967] = {-9'd61,-10'd261};
ram[10968] = {-9'd58,-10'd258};
ram[10969] = {-9'd55,-10'd255};
ram[10970] = {-9'd52,-10'd252};
ram[10971] = {-9'd48,-10'd249};
ram[10972] = {-9'd45,-10'd246};
ram[10973] = {-9'd42,-10'd242};
ram[10974] = {-9'd39,-10'd239};
ram[10975] = {-9'd36,-10'd236};
ram[10976] = {-9'd33,-10'd233};
ram[10977] = {-9'd30,-10'd230};
ram[10978] = {-9'd26,-10'd227};
ram[10979] = {-9'd23,-10'd224};
ram[10980] = {-9'd20,-10'd220};
ram[10981] = {-9'd17,-10'd217};
ram[10982] = {-9'd14,-10'd214};
ram[10983] = {-9'd11,-10'd211};
ram[10984] = {-9'd8,-10'd208};
ram[10985] = {-9'd4,-10'd205};
ram[10986] = {-9'd1,-10'd202};
ram[10987] = {9'd2,-10'd198};
ram[10988] = {9'd5,-10'd195};
ram[10989] = {9'd8,-10'd192};
ram[10990] = {9'd11,-10'd189};
ram[10991] = {9'd14,-10'd186};
ram[10992] = {9'd18,-10'd183};
ram[10993] = {9'd21,-10'd180};
ram[10994] = {9'd24,-10'd176};
ram[10995] = {9'd27,-10'd173};
ram[10996] = {9'd30,-10'd170};
ram[10997] = {9'd33,-10'd167};
ram[10998] = {9'd36,-10'd164};
ram[10999] = {9'd40,-10'd161};
ram[11000] = {9'd43,-10'd158};
ram[11001] = {9'd46,-10'd154};
ram[11002] = {9'd49,-10'd151};
ram[11003] = {9'd52,-10'd148};
ram[11004] = {9'd55,-10'd145};
ram[11005] = {9'd58,-10'd142};
ram[11006] = {9'd62,-10'd139};
ram[11007] = {9'd65,-10'd136};
ram[11008] = {9'd65,-10'd136};
ram[11009] = {9'd68,-10'd132};
ram[11010] = {9'd71,-10'd129};
ram[11011] = {9'd74,-10'd126};
ram[11012] = {9'd77,-10'd123};
ram[11013] = {9'd80,-10'd120};
ram[11014] = {9'd84,-10'd117};
ram[11015] = {9'd87,-10'd114};
ram[11016] = {9'd90,-10'd110};
ram[11017] = {9'd93,-10'd107};
ram[11018] = {9'd96,-10'd104};
ram[11019] = {9'd99,-10'd101};
ram[11020] = {-9'd98,-10'd98};
ram[11021] = {-9'd95,-10'd95};
ram[11022] = {-9'd92,-10'd92};
ram[11023] = {-9'd88,-10'd88};
ram[11024] = {-9'd85,-10'd85};
ram[11025] = {-9'd82,-10'd82};
ram[11026] = {-9'd79,-10'd79};
ram[11027] = {-9'd76,-10'd76};
ram[11028] = {-9'd73,-10'd73};
ram[11029] = {-9'd70,-10'd70};
ram[11030] = {-9'd66,-10'd66};
ram[11031] = {-9'd63,-10'd63};
ram[11032] = {-9'd60,-10'd60};
ram[11033] = {-9'd57,-10'd57};
ram[11034] = {-9'd54,-10'd54};
ram[11035] = {-9'd51,-10'd51};
ram[11036] = {-9'd48,-10'd48};
ram[11037] = {-9'd44,-10'd44};
ram[11038] = {-9'd41,-10'd41};
ram[11039] = {-9'd38,-10'd38};
ram[11040] = {-9'd35,-10'd35};
ram[11041] = {-9'd32,-10'd32};
ram[11042] = {-9'd29,-10'd29};
ram[11043] = {-9'd26,-10'd26};
ram[11044] = {-9'd22,-10'd22};
ram[11045] = {-9'd19,-10'd19};
ram[11046] = {-9'd16,-10'd16};
ram[11047] = {-9'd13,-10'd13};
ram[11048] = {-9'd10,-10'd10};
ram[11049] = {-9'd7,-10'd7};
ram[11050] = {-9'd4,-10'd4};
ram[11051] = {9'd0,10'd0};
ram[11052] = {9'd3,10'd3};
ram[11053] = {9'd6,10'd6};
ram[11054] = {9'd9,10'd9};
ram[11055] = {9'd12,10'd12};
ram[11056] = {9'd15,10'd15};
ram[11057] = {9'd18,10'd18};
ram[11058] = {9'd21,10'd21};
ram[11059] = {9'd25,10'd25};
ram[11060] = {9'd28,10'd28};
ram[11061] = {9'd31,10'd31};
ram[11062] = {9'd34,10'd34};
ram[11063] = {9'd37,10'd37};
ram[11064] = {9'd40,10'd40};
ram[11065] = {9'd43,10'd43};
ram[11066] = {9'd47,10'd47};
ram[11067] = {9'd50,10'd50};
ram[11068] = {9'd53,10'd53};
ram[11069] = {9'd56,10'd56};
ram[11070] = {9'd59,10'd59};
ram[11071] = {9'd62,10'd62};
ram[11072] = {9'd65,10'd65};
ram[11073] = {9'd69,10'd69};
ram[11074] = {9'd72,10'd72};
ram[11075] = {9'd75,10'd75};
ram[11076] = {9'd78,10'd78};
ram[11077] = {9'd81,10'd81};
ram[11078] = {9'd84,10'd84};
ram[11079] = {9'd87,10'd87};
ram[11080] = {9'd91,10'd91};
ram[11081] = {9'd94,10'd94};
ram[11082] = {9'd97,10'd97};
ram[11083] = {-9'd100,10'd100};
ram[11084] = {-9'd97,10'd103};
ram[11085] = {-9'd94,10'd106};
ram[11086] = {-9'd91,10'd109};
ram[11087] = {-9'd88,10'd113};
ram[11088] = {-9'd85,10'd116};
ram[11089] = {-9'd81,10'd119};
ram[11090] = {-9'd78,10'd122};
ram[11091] = {-9'd75,10'd125};
ram[11092] = {-9'd72,10'd128};
ram[11093] = {-9'd69,10'd131};
ram[11094] = {-9'd66,10'd135};
ram[11095] = {-9'd63,10'd138};
ram[11096] = {-9'd59,10'd141};
ram[11097] = {-9'd56,10'd144};
ram[11098] = {-9'd53,10'd147};
ram[11099] = {-9'd50,10'd150};
ram[11100] = {-9'd47,10'd153};
ram[11101] = {-9'd44,10'd157};
ram[11102] = {-9'd41,10'd160};
ram[11103] = {-9'd37,10'd163};
ram[11104] = {-9'd34,10'd166};
ram[11105] = {-9'd31,10'd169};
ram[11106] = {-9'd28,10'd172};
ram[11107] = {-9'd25,10'd175};
ram[11108] = {-9'd22,10'd179};
ram[11109] = {-9'd19,10'd182};
ram[11110] = {-9'd15,10'd185};
ram[11111] = {-9'd12,10'd188};
ram[11112] = {-9'd9,10'd191};
ram[11113] = {-9'd6,10'd194};
ram[11114] = {-9'd3,10'd197};
ram[11115] = {9'd0,10'd201};
ram[11116] = {9'd3,10'd204};
ram[11117] = {9'd7,10'd207};
ram[11118] = {9'd10,10'd210};
ram[11119] = {9'd13,10'd213};
ram[11120] = {9'd16,10'd216};
ram[11121] = {9'd19,10'd219};
ram[11122] = {9'd22,10'd223};
ram[11123] = {9'd25,10'd226};
ram[11124] = {9'd29,10'd229};
ram[11125] = {9'd32,10'd232};
ram[11126] = {9'd35,10'd235};
ram[11127] = {9'd38,10'd238};
ram[11128] = {9'd41,10'd241};
ram[11129] = {9'd44,10'd245};
ram[11130] = {9'd47,10'd248};
ram[11131] = {9'd51,10'd251};
ram[11132] = {9'd54,10'd254};
ram[11133] = {9'd57,10'd257};
ram[11134] = {9'd60,10'd260};
ram[11135] = {9'd63,10'd263};
ram[11136] = {9'd63,10'd263};
ram[11137] = {9'd66,10'd267};
ram[11138] = {9'd69,10'd270};
ram[11139] = {9'd73,10'd273};
ram[11140] = {9'd76,10'd276};
ram[11141] = {9'd79,10'd279};
ram[11142] = {9'd82,10'd282};
ram[11143] = {9'd85,10'd285};
ram[11144] = {9'd88,10'd289};
ram[11145] = {9'd91,10'd292};
ram[11146] = {9'd95,10'd295};
ram[11147] = {9'd98,10'd298};
ram[11148] = {-9'd99,10'd301};
ram[11149] = {-9'd96,10'd304};
ram[11150] = {-9'd93,10'd307};
ram[11151] = {-9'd90,10'd311};
ram[11152] = {-9'd87,10'd314};
ram[11153] = {-9'd84,10'd317};
ram[11154] = {-9'd81,10'd320};
ram[11155] = {-9'd77,10'd323};
ram[11156] = {-9'd74,10'd326};
ram[11157] = {-9'd71,10'd329};
ram[11158] = {-9'd68,10'd333};
ram[11159] = {-9'd65,10'd336};
ram[11160] = {-9'd62,10'd339};
ram[11161] = {-9'd59,10'd342};
ram[11162] = {-9'd55,10'd345};
ram[11163] = {-9'd52,10'd348};
ram[11164] = {-9'd49,10'd351};
ram[11165] = {-9'd46,10'd354};
ram[11166] = {-9'd43,10'd358};
ram[11167] = {-9'd40,10'd361};
ram[11168] = {-9'd37,10'd364};
ram[11169] = {-9'd33,10'd367};
ram[11170] = {-9'd30,10'd370};
ram[11171] = {-9'd27,10'd373};
ram[11172] = {-9'd24,10'd376};
ram[11173] = {-9'd21,10'd380};
ram[11174] = {-9'd18,10'd383};
ram[11175] = {-9'd15,10'd386};
ram[11176] = {-9'd11,10'd389};
ram[11177] = {-9'd8,10'd392};
ram[11178] = {-9'd5,10'd395};
ram[11179] = {-9'd2,10'd398};
ram[11180] = {9'd1,-10'd399};
ram[11181] = {9'd4,-10'd396};
ram[11182] = {9'd7,-10'd393};
ram[11183] = {9'd10,-10'd390};
ram[11184] = {9'd14,-10'd387};
ram[11185] = {9'd17,-10'd384};
ram[11186] = {9'd20,-10'd381};
ram[11187] = {9'd23,-10'd377};
ram[11188] = {9'd26,-10'd374};
ram[11189] = {9'd29,-10'd371};
ram[11190] = {9'd32,-10'd368};
ram[11191] = {9'd36,-10'd365};
ram[11192] = {9'd39,-10'd362};
ram[11193] = {9'd42,-10'd359};
ram[11194] = {9'd45,-10'd355};
ram[11195] = {9'd48,-10'd352};
ram[11196] = {9'd51,-10'd349};
ram[11197] = {9'd54,-10'd346};
ram[11198] = {9'd58,-10'd343};
ram[11199] = {9'd61,-10'd340};
ram[11200] = {9'd64,-10'd337};
ram[11201] = {9'd67,-10'd334};
ram[11202] = {9'd70,-10'd330};
ram[11203] = {9'd73,-10'd327};
ram[11204] = {9'd76,-10'd324};
ram[11205] = {9'd80,-10'd321};
ram[11206] = {9'd83,-10'd318};
ram[11207] = {9'd86,-10'd315};
ram[11208] = {9'd89,-10'd312};
ram[11209] = {9'd92,-10'd308};
ram[11210] = {9'd95,-10'd305};
ram[11211] = {9'd98,-10'd302};
ram[11212] = {-9'd99,-10'd299};
ram[11213] = {-9'd96,-10'd296};
ram[11214] = {-9'd92,-10'd293};
ram[11215] = {-9'd89,-10'd290};
ram[11216] = {-9'd86,-10'd286};
ram[11217] = {-9'd83,-10'd283};
ram[11218] = {-9'd80,-10'd280};
ram[11219] = {-9'd77,-10'd277};
ram[11220] = {-9'd74,-10'd274};
ram[11221] = {-9'd70,-10'd271};
ram[11222] = {-9'd67,-10'd268};
ram[11223] = {-9'd64,-10'd264};
ram[11224] = {-9'd61,-10'd261};
ram[11225] = {-9'd58,-10'd258};
ram[11226] = {-9'd55,-10'd255};
ram[11227] = {-9'd52,-10'd252};
ram[11228] = {-9'd48,-10'd249};
ram[11229] = {-9'd45,-10'd246};
ram[11230] = {-9'd42,-10'd242};
ram[11231] = {-9'd39,-10'd239};
ram[11232] = {-9'd36,-10'd236};
ram[11233] = {-9'd33,-10'd233};
ram[11234] = {-9'd30,-10'd230};
ram[11235] = {-9'd26,-10'd227};
ram[11236] = {-9'd23,-10'd224};
ram[11237] = {-9'd20,-10'd220};
ram[11238] = {-9'd17,-10'd217};
ram[11239] = {-9'd14,-10'd214};
ram[11240] = {-9'd11,-10'd211};
ram[11241] = {-9'd8,-10'd208};
ram[11242] = {-9'd4,-10'd205};
ram[11243] = {-9'd1,-10'd202};
ram[11244] = {9'd2,-10'd198};
ram[11245] = {9'd5,-10'd195};
ram[11246] = {9'd8,-10'd192};
ram[11247] = {9'd11,-10'd189};
ram[11248] = {9'd14,-10'd186};
ram[11249] = {9'd18,-10'd183};
ram[11250] = {9'd21,-10'd180};
ram[11251] = {9'd24,-10'd176};
ram[11252] = {9'd27,-10'd173};
ram[11253] = {9'd30,-10'd170};
ram[11254] = {9'd33,-10'd167};
ram[11255] = {9'd36,-10'd164};
ram[11256] = {9'd40,-10'd161};
ram[11257] = {9'd43,-10'd158};
ram[11258] = {9'd46,-10'd154};
ram[11259] = {9'd49,-10'd151};
ram[11260] = {9'd52,-10'd148};
ram[11261] = {9'd55,-10'd145};
ram[11262] = {9'd58,-10'd142};
ram[11263] = {9'd62,-10'd139};
ram[11264] = {9'd62,-10'd139};
ram[11265] = {9'd65,-10'd136};
ram[11266] = {9'd68,-10'd132};
ram[11267] = {9'd71,-10'd129};
ram[11268] = {9'd74,-10'd126};
ram[11269] = {9'd77,-10'd123};
ram[11270] = {9'd80,-10'd120};
ram[11271] = {9'd84,-10'd117};
ram[11272] = {9'd87,-10'd114};
ram[11273] = {9'd90,-10'd110};
ram[11274] = {9'd93,-10'd107};
ram[11275] = {9'd96,-10'd104};
ram[11276] = {9'd99,-10'd101};
ram[11277] = {-9'd98,-10'd98};
ram[11278] = {-9'd95,-10'd95};
ram[11279] = {-9'd92,-10'd92};
ram[11280] = {-9'd88,-10'd88};
ram[11281] = {-9'd85,-10'd85};
ram[11282] = {-9'd82,-10'd82};
ram[11283] = {-9'd79,-10'd79};
ram[11284] = {-9'd76,-10'd76};
ram[11285] = {-9'd73,-10'd73};
ram[11286] = {-9'd70,-10'd70};
ram[11287] = {-9'd66,-10'd66};
ram[11288] = {-9'd63,-10'd63};
ram[11289] = {-9'd60,-10'd60};
ram[11290] = {-9'd57,-10'd57};
ram[11291] = {-9'd54,-10'd54};
ram[11292] = {-9'd51,-10'd51};
ram[11293] = {-9'd48,-10'd48};
ram[11294] = {-9'd44,-10'd44};
ram[11295] = {-9'd41,-10'd41};
ram[11296] = {-9'd38,-10'd38};
ram[11297] = {-9'd35,-10'd35};
ram[11298] = {-9'd32,-10'd32};
ram[11299] = {-9'd29,-10'd29};
ram[11300] = {-9'd26,-10'd26};
ram[11301] = {-9'd22,-10'd22};
ram[11302] = {-9'd19,-10'd19};
ram[11303] = {-9'd16,-10'd16};
ram[11304] = {-9'd13,-10'd13};
ram[11305] = {-9'd10,-10'd10};
ram[11306] = {-9'd7,-10'd7};
ram[11307] = {-9'd4,-10'd4};
ram[11308] = {9'd0,10'd0};
ram[11309] = {9'd3,10'd3};
ram[11310] = {9'd6,10'd6};
ram[11311] = {9'd9,10'd9};
ram[11312] = {9'd12,10'd12};
ram[11313] = {9'd15,10'd15};
ram[11314] = {9'd18,10'd18};
ram[11315] = {9'd21,10'd21};
ram[11316] = {9'd25,10'd25};
ram[11317] = {9'd28,10'd28};
ram[11318] = {9'd31,10'd31};
ram[11319] = {9'd34,10'd34};
ram[11320] = {9'd37,10'd37};
ram[11321] = {9'd40,10'd40};
ram[11322] = {9'd43,10'd43};
ram[11323] = {9'd47,10'd47};
ram[11324] = {9'd50,10'd50};
ram[11325] = {9'd53,10'd53};
ram[11326] = {9'd56,10'd56};
ram[11327] = {9'd59,10'd59};
ram[11328] = {9'd62,10'd62};
ram[11329] = {9'd65,10'd65};
ram[11330] = {9'd69,10'd69};
ram[11331] = {9'd72,10'd72};
ram[11332] = {9'd75,10'd75};
ram[11333] = {9'd78,10'd78};
ram[11334] = {9'd81,10'd81};
ram[11335] = {9'd84,10'd84};
ram[11336] = {9'd87,10'd87};
ram[11337] = {9'd91,10'd91};
ram[11338] = {9'd94,10'd94};
ram[11339] = {9'd97,10'd97};
ram[11340] = {-9'd100,10'd100};
ram[11341] = {-9'd97,10'd103};
ram[11342] = {-9'd94,10'd106};
ram[11343] = {-9'd91,10'd109};
ram[11344] = {-9'd88,10'd113};
ram[11345] = {-9'd85,10'd116};
ram[11346] = {-9'd81,10'd119};
ram[11347] = {-9'd78,10'd122};
ram[11348] = {-9'd75,10'd125};
ram[11349] = {-9'd72,10'd128};
ram[11350] = {-9'd69,10'd131};
ram[11351] = {-9'd66,10'd135};
ram[11352] = {-9'd63,10'd138};
ram[11353] = {-9'd59,10'd141};
ram[11354] = {-9'd56,10'd144};
ram[11355] = {-9'd53,10'd147};
ram[11356] = {-9'd50,10'd150};
ram[11357] = {-9'd47,10'd153};
ram[11358] = {-9'd44,10'd157};
ram[11359] = {-9'd41,10'd160};
ram[11360] = {-9'd37,10'd163};
ram[11361] = {-9'd34,10'd166};
ram[11362] = {-9'd31,10'd169};
ram[11363] = {-9'd28,10'd172};
ram[11364] = {-9'd25,10'd175};
ram[11365] = {-9'd22,10'd179};
ram[11366] = {-9'd19,10'd182};
ram[11367] = {-9'd15,10'd185};
ram[11368] = {-9'd12,10'd188};
ram[11369] = {-9'd9,10'd191};
ram[11370] = {-9'd6,10'd194};
ram[11371] = {-9'd3,10'd197};
ram[11372] = {9'd0,10'd201};
ram[11373] = {9'd3,10'd204};
ram[11374] = {9'd7,10'd207};
ram[11375] = {9'd10,10'd210};
ram[11376] = {9'd13,10'd213};
ram[11377] = {9'd16,10'd216};
ram[11378] = {9'd19,10'd219};
ram[11379] = {9'd22,10'd223};
ram[11380] = {9'd25,10'd226};
ram[11381] = {9'd29,10'd229};
ram[11382] = {9'd32,10'd232};
ram[11383] = {9'd35,10'd235};
ram[11384] = {9'd38,10'd238};
ram[11385] = {9'd41,10'd241};
ram[11386] = {9'd44,10'd245};
ram[11387] = {9'd47,10'd248};
ram[11388] = {9'd51,10'd251};
ram[11389] = {9'd54,10'd254};
ram[11390] = {9'd57,10'd257};
ram[11391] = {9'd60,10'd260};
ram[11392] = {9'd60,10'd260};
ram[11393] = {9'd63,10'd263};
ram[11394] = {9'd66,10'd267};
ram[11395] = {9'd69,10'd270};
ram[11396] = {9'd73,10'd273};
ram[11397] = {9'd76,10'd276};
ram[11398] = {9'd79,10'd279};
ram[11399] = {9'd82,10'd282};
ram[11400] = {9'd85,10'd285};
ram[11401] = {9'd88,10'd289};
ram[11402] = {9'd91,10'd292};
ram[11403] = {9'd95,10'd295};
ram[11404] = {9'd98,10'd298};
ram[11405] = {-9'd99,10'd301};
ram[11406] = {-9'd96,10'd304};
ram[11407] = {-9'd93,10'd307};
ram[11408] = {-9'd90,10'd311};
ram[11409] = {-9'd87,10'd314};
ram[11410] = {-9'd84,10'd317};
ram[11411] = {-9'd81,10'd320};
ram[11412] = {-9'd77,10'd323};
ram[11413] = {-9'd74,10'd326};
ram[11414] = {-9'd71,10'd329};
ram[11415] = {-9'd68,10'd333};
ram[11416] = {-9'd65,10'd336};
ram[11417] = {-9'd62,10'd339};
ram[11418] = {-9'd59,10'd342};
ram[11419] = {-9'd55,10'd345};
ram[11420] = {-9'd52,10'd348};
ram[11421] = {-9'd49,10'd351};
ram[11422] = {-9'd46,10'd354};
ram[11423] = {-9'd43,10'd358};
ram[11424] = {-9'd40,10'd361};
ram[11425] = {-9'd37,10'd364};
ram[11426] = {-9'd33,10'd367};
ram[11427] = {-9'd30,10'd370};
ram[11428] = {-9'd27,10'd373};
ram[11429] = {-9'd24,10'd376};
ram[11430] = {-9'd21,10'd380};
ram[11431] = {-9'd18,10'd383};
ram[11432] = {-9'd15,10'd386};
ram[11433] = {-9'd11,10'd389};
ram[11434] = {-9'd8,10'd392};
ram[11435] = {-9'd5,10'd395};
ram[11436] = {-9'd2,10'd398};
ram[11437] = {9'd1,-10'd399};
ram[11438] = {9'd4,-10'd396};
ram[11439] = {9'd7,-10'd393};
ram[11440] = {9'd10,-10'd390};
ram[11441] = {9'd14,-10'd387};
ram[11442] = {9'd17,-10'd384};
ram[11443] = {9'd20,-10'd381};
ram[11444] = {9'd23,-10'd377};
ram[11445] = {9'd26,-10'd374};
ram[11446] = {9'd29,-10'd371};
ram[11447] = {9'd32,-10'd368};
ram[11448] = {9'd36,-10'd365};
ram[11449] = {9'd39,-10'd362};
ram[11450] = {9'd42,-10'd359};
ram[11451] = {9'd45,-10'd355};
ram[11452] = {9'd48,-10'd352};
ram[11453] = {9'd51,-10'd349};
ram[11454] = {9'd54,-10'd346};
ram[11455] = {9'd58,-10'd343};
ram[11456] = {9'd61,-10'd340};
ram[11457] = {9'd64,-10'd337};
ram[11458] = {9'd67,-10'd334};
ram[11459] = {9'd70,-10'd330};
ram[11460] = {9'd73,-10'd327};
ram[11461] = {9'd76,-10'd324};
ram[11462] = {9'd80,-10'd321};
ram[11463] = {9'd83,-10'd318};
ram[11464] = {9'd86,-10'd315};
ram[11465] = {9'd89,-10'd312};
ram[11466] = {9'd92,-10'd308};
ram[11467] = {9'd95,-10'd305};
ram[11468] = {9'd98,-10'd302};
ram[11469] = {-9'd99,-10'd299};
ram[11470] = {-9'd96,-10'd296};
ram[11471] = {-9'd92,-10'd293};
ram[11472] = {-9'd89,-10'd290};
ram[11473] = {-9'd86,-10'd286};
ram[11474] = {-9'd83,-10'd283};
ram[11475] = {-9'd80,-10'd280};
ram[11476] = {-9'd77,-10'd277};
ram[11477] = {-9'd74,-10'd274};
ram[11478] = {-9'd70,-10'd271};
ram[11479] = {-9'd67,-10'd268};
ram[11480] = {-9'd64,-10'd264};
ram[11481] = {-9'd61,-10'd261};
ram[11482] = {-9'd58,-10'd258};
ram[11483] = {-9'd55,-10'd255};
ram[11484] = {-9'd52,-10'd252};
ram[11485] = {-9'd48,-10'd249};
ram[11486] = {-9'd45,-10'd246};
ram[11487] = {-9'd42,-10'd242};
ram[11488] = {-9'd39,-10'd239};
ram[11489] = {-9'd36,-10'd236};
ram[11490] = {-9'd33,-10'd233};
ram[11491] = {-9'd30,-10'd230};
ram[11492] = {-9'd26,-10'd227};
ram[11493] = {-9'd23,-10'd224};
ram[11494] = {-9'd20,-10'd220};
ram[11495] = {-9'd17,-10'd217};
ram[11496] = {-9'd14,-10'd214};
ram[11497] = {-9'd11,-10'd211};
ram[11498] = {-9'd8,-10'd208};
ram[11499] = {-9'd4,-10'd205};
ram[11500] = {-9'd1,-10'd202};
ram[11501] = {9'd2,-10'd198};
ram[11502] = {9'd5,-10'd195};
ram[11503] = {9'd8,-10'd192};
ram[11504] = {9'd11,-10'd189};
ram[11505] = {9'd14,-10'd186};
ram[11506] = {9'd18,-10'd183};
ram[11507] = {9'd21,-10'd180};
ram[11508] = {9'd24,-10'd176};
ram[11509] = {9'd27,-10'd173};
ram[11510] = {9'd30,-10'd170};
ram[11511] = {9'd33,-10'd167};
ram[11512] = {9'd36,-10'd164};
ram[11513] = {9'd40,-10'd161};
ram[11514] = {9'd43,-10'd158};
ram[11515] = {9'd46,-10'd154};
ram[11516] = {9'd49,-10'd151};
ram[11517] = {9'd52,-10'd148};
ram[11518] = {9'd55,-10'd145};
ram[11519] = {9'd58,-10'd142};
ram[11520] = {9'd58,-10'd142};
ram[11521] = {9'd62,-10'd139};
ram[11522] = {9'd65,-10'd136};
ram[11523] = {9'd68,-10'd132};
ram[11524] = {9'd71,-10'd129};
ram[11525] = {9'd74,-10'd126};
ram[11526] = {9'd77,-10'd123};
ram[11527] = {9'd80,-10'd120};
ram[11528] = {9'd84,-10'd117};
ram[11529] = {9'd87,-10'd114};
ram[11530] = {9'd90,-10'd110};
ram[11531] = {9'd93,-10'd107};
ram[11532] = {9'd96,-10'd104};
ram[11533] = {9'd99,-10'd101};
ram[11534] = {-9'd98,-10'd98};
ram[11535] = {-9'd95,-10'd95};
ram[11536] = {-9'd92,-10'd92};
ram[11537] = {-9'd88,-10'd88};
ram[11538] = {-9'd85,-10'd85};
ram[11539] = {-9'd82,-10'd82};
ram[11540] = {-9'd79,-10'd79};
ram[11541] = {-9'd76,-10'd76};
ram[11542] = {-9'd73,-10'd73};
ram[11543] = {-9'd70,-10'd70};
ram[11544] = {-9'd66,-10'd66};
ram[11545] = {-9'd63,-10'd63};
ram[11546] = {-9'd60,-10'd60};
ram[11547] = {-9'd57,-10'd57};
ram[11548] = {-9'd54,-10'd54};
ram[11549] = {-9'd51,-10'd51};
ram[11550] = {-9'd48,-10'd48};
ram[11551] = {-9'd44,-10'd44};
ram[11552] = {-9'd41,-10'd41};
ram[11553] = {-9'd38,-10'd38};
ram[11554] = {-9'd35,-10'd35};
ram[11555] = {-9'd32,-10'd32};
ram[11556] = {-9'd29,-10'd29};
ram[11557] = {-9'd26,-10'd26};
ram[11558] = {-9'd22,-10'd22};
ram[11559] = {-9'd19,-10'd19};
ram[11560] = {-9'd16,-10'd16};
ram[11561] = {-9'd13,-10'd13};
ram[11562] = {-9'd10,-10'd10};
ram[11563] = {-9'd7,-10'd7};
ram[11564] = {-9'd4,-10'd4};
ram[11565] = {9'd0,10'd0};
ram[11566] = {9'd3,10'd3};
ram[11567] = {9'd6,10'd6};
ram[11568] = {9'd9,10'd9};
ram[11569] = {9'd12,10'd12};
ram[11570] = {9'd15,10'd15};
ram[11571] = {9'd18,10'd18};
ram[11572] = {9'd21,10'd21};
ram[11573] = {9'd25,10'd25};
ram[11574] = {9'd28,10'd28};
ram[11575] = {9'd31,10'd31};
ram[11576] = {9'd34,10'd34};
ram[11577] = {9'd37,10'd37};
ram[11578] = {9'd40,10'd40};
ram[11579] = {9'd43,10'd43};
ram[11580] = {9'd47,10'd47};
ram[11581] = {9'd50,10'd50};
ram[11582] = {9'd53,10'd53};
ram[11583] = {9'd56,10'd56};
ram[11584] = {9'd59,10'd59};
ram[11585] = {9'd62,10'd62};
ram[11586] = {9'd65,10'd65};
ram[11587] = {9'd69,10'd69};
ram[11588] = {9'd72,10'd72};
ram[11589] = {9'd75,10'd75};
ram[11590] = {9'd78,10'd78};
ram[11591] = {9'd81,10'd81};
ram[11592] = {9'd84,10'd84};
ram[11593] = {9'd87,10'd87};
ram[11594] = {9'd91,10'd91};
ram[11595] = {9'd94,10'd94};
ram[11596] = {9'd97,10'd97};
ram[11597] = {-9'd100,10'd100};
ram[11598] = {-9'd97,10'd103};
ram[11599] = {-9'd94,10'd106};
ram[11600] = {-9'd91,10'd109};
ram[11601] = {-9'd88,10'd113};
ram[11602] = {-9'd85,10'd116};
ram[11603] = {-9'd81,10'd119};
ram[11604] = {-9'd78,10'd122};
ram[11605] = {-9'd75,10'd125};
ram[11606] = {-9'd72,10'd128};
ram[11607] = {-9'd69,10'd131};
ram[11608] = {-9'd66,10'd135};
ram[11609] = {-9'd63,10'd138};
ram[11610] = {-9'd59,10'd141};
ram[11611] = {-9'd56,10'd144};
ram[11612] = {-9'd53,10'd147};
ram[11613] = {-9'd50,10'd150};
ram[11614] = {-9'd47,10'd153};
ram[11615] = {-9'd44,10'd157};
ram[11616] = {-9'd41,10'd160};
ram[11617] = {-9'd37,10'd163};
ram[11618] = {-9'd34,10'd166};
ram[11619] = {-9'd31,10'd169};
ram[11620] = {-9'd28,10'd172};
ram[11621] = {-9'd25,10'd175};
ram[11622] = {-9'd22,10'd179};
ram[11623] = {-9'd19,10'd182};
ram[11624] = {-9'd15,10'd185};
ram[11625] = {-9'd12,10'd188};
ram[11626] = {-9'd9,10'd191};
ram[11627] = {-9'd6,10'd194};
ram[11628] = {-9'd3,10'd197};
ram[11629] = {9'd0,10'd201};
ram[11630] = {9'd3,10'd204};
ram[11631] = {9'd7,10'd207};
ram[11632] = {9'd10,10'd210};
ram[11633] = {9'd13,10'd213};
ram[11634] = {9'd16,10'd216};
ram[11635] = {9'd19,10'd219};
ram[11636] = {9'd22,10'd223};
ram[11637] = {9'd25,10'd226};
ram[11638] = {9'd29,10'd229};
ram[11639] = {9'd32,10'd232};
ram[11640] = {9'd35,10'd235};
ram[11641] = {9'd38,10'd238};
ram[11642] = {9'd41,10'd241};
ram[11643] = {9'd44,10'd245};
ram[11644] = {9'd47,10'd248};
ram[11645] = {9'd51,10'd251};
ram[11646] = {9'd54,10'd254};
ram[11647] = {9'd57,10'd257};
ram[11648] = {9'd57,10'd257};
ram[11649] = {9'd60,10'd260};
ram[11650] = {9'd63,10'd263};
ram[11651] = {9'd66,10'd267};
ram[11652] = {9'd69,10'd270};
ram[11653] = {9'd73,10'd273};
ram[11654] = {9'd76,10'd276};
ram[11655] = {9'd79,10'd279};
ram[11656] = {9'd82,10'd282};
ram[11657] = {9'd85,10'd285};
ram[11658] = {9'd88,10'd289};
ram[11659] = {9'd91,10'd292};
ram[11660] = {9'd95,10'd295};
ram[11661] = {9'd98,10'd298};
ram[11662] = {-9'd99,10'd301};
ram[11663] = {-9'd96,10'd304};
ram[11664] = {-9'd93,10'd307};
ram[11665] = {-9'd90,10'd311};
ram[11666] = {-9'd87,10'd314};
ram[11667] = {-9'd84,10'd317};
ram[11668] = {-9'd81,10'd320};
ram[11669] = {-9'd77,10'd323};
ram[11670] = {-9'd74,10'd326};
ram[11671] = {-9'd71,10'd329};
ram[11672] = {-9'd68,10'd333};
ram[11673] = {-9'd65,10'd336};
ram[11674] = {-9'd62,10'd339};
ram[11675] = {-9'd59,10'd342};
ram[11676] = {-9'd55,10'd345};
ram[11677] = {-9'd52,10'd348};
ram[11678] = {-9'd49,10'd351};
ram[11679] = {-9'd46,10'd354};
ram[11680] = {-9'd43,10'd358};
ram[11681] = {-9'd40,10'd361};
ram[11682] = {-9'd37,10'd364};
ram[11683] = {-9'd33,10'd367};
ram[11684] = {-9'd30,10'd370};
ram[11685] = {-9'd27,10'd373};
ram[11686] = {-9'd24,10'd376};
ram[11687] = {-9'd21,10'd380};
ram[11688] = {-9'd18,10'd383};
ram[11689] = {-9'd15,10'd386};
ram[11690] = {-9'd11,10'd389};
ram[11691] = {-9'd8,10'd392};
ram[11692] = {-9'd5,10'd395};
ram[11693] = {-9'd2,10'd398};
ram[11694] = {9'd1,-10'd399};
ram[11695] = {9'd4,-10'd396};
ram[11696] = {9'd7,-10'd393};
ram[11697] = {9'd10,-10'd390};
ram[11698] = {9'd14,-10'd387};
ram[11699] = {9'd17,-10'd384};
ram[11700] = {9'd20,-10'd381};
ram[11701] = {9'd23,-10'd377};
ram[11702] = {9'd26,-10'd374};
ram[11703] = {9'd29,-10'd371};
ram[11704] = {9'd32,-10'd368};
ram[11705] = {9'd36,-10'd365};
ram[11706] = {9'd39,-10'd362};
ram[11707] = {9'd42,-10'd359};
ram[11708] = {9'd45,-10'd355};
ram[11709] = {9'd48,-10'd352};
ram[11710] = {9'd51,-10'd349};
ram[11711] = {9'd54,-10'd346};
ram[11712] = {9'd58,-10'd343};
ram[11713] = {9'd61,-10'd340};
ram[11714] = {9'd64,-10'd337};
ram[11715] = {9'd67,-10'd334};
ram[11716] = {9'd70,-10'd330};
ram[11717] = {9'd73,-10'd327};
ram[11718] = {9'd76,-10'd324};
ram[11719] = {9'd80,-10'd321};
ram[11720] = {9'd83,-10'd318};
ram[11721] = {9'd86,-10'd315};
ram[11722] = {9'd89,-10'd312};
ram[11723] = {9'd92,-10'd308};
ram[11724] = {9'd95,-10'd305};
ram[11725] = {9'd98,-10'd302};
ram[11726] = {-9'd99,-10'd299};
ram[11727] = {-9'd96,-10'd296};
ram[11728] = {-9'd92,-10'd293};
ram[11729] = {-9'd89,-10'd290};
ram[11730] = {-9'd86,-10'd286};
ram[11731] = {-9'd83,-10'd283};
ram[11732] = {-9'd80,-10'd280};
ram[11733] = {-9'd77,-10'd277};
ram[11734] = {-9'd74,-10'd274};
ram[11735] = {-9'd70,-10'd271};
ram[11736] = {-9'd67,-10'd268};
ram[11737] = {-9'd64,-10'd264};
ram[11738] = {-9'd61,-10'd261};
ram[11739] = {-9'd58,-10'd258};
ram[11740] = {-9'd55,-10'd255};
ram[11741] = {-9'd52,-10'd252};
ram[11742] = {-9'd48,-10'd249};
ram[11743] = {-9'd45,-10'd246};
ram[11744] = {-9'd42,-10'd242};
ram[11745] = {-9'd39,-10'd239};
ram[11746] = {-9'd36,-10'd236};
ram[11747] = {-9'd33,-10'd233};
ram[11748] = {-9'd30,-10'd230};
ram[11749] = {-9'd26,-10'd227};
ram[11750] = {-9'd23,-10'd224};
ram[11751] = {-9'd20,-10'd220};
ram[11752] = {-9'd17,-10'd217};
ram[11753] = {-9'd14,-10'd214};
ram[11754] = {-9'd11,-10'd211};
ram[11755] = {-9'd8,-10'd208};
ram[11756] = {-9'd4,-10'd205};
ram[11757] = {-9'd1,-10'd202};
ram[11758] = {9'd2,-10'd198};
ram[11759] = {9'd5,-10'd195};
ram[11760] = {9'd8,-10'd192};
ram[11761] = {9'd11,-10'd189};
ram[11762] = {9'd14,-10'd186};
ram[11763] = {9'd18,-10'd183};
ram[11764] = {9'd21,-10'd180};
ram[11765] = {9'd24,-10'd176};
ram[11766] = {9'd27,-10'd173};
ram[11767] = {9'd30,-10'd170};
ram[11768] = {9'd33,-10'd167};
ram[11769] = {9'd36,-10'd164};
ram[11770] = {9'd40,-10'd161};
ram[11771] = {9'd43,-10'd158};
ram[11772] = {9'd46,-10'd154};
ram[11773] = {9'd49,-10'd151};
ram[11774] = {9'd52,-10'd148};
ram[11775] = {9'd55,-10'd145};
ram[11776] = {9'd55,-10'd145};
ram[11777] = {9'd58,-10'd142};
ram[11778] = {9'd62,-10'd139};
ram[11779] = {9'd65,-10'd136};
ram[11780] = {9'd68,-10'd132};
ram[11781] = {9'd71,-10'd129};
ram[11782] = {9'd74,-10'd126};
ram[11783] = {9'd77,-10'd123};
ram[11784] = {9'd80,-10'd120};
ram[11785] = {9'd84,-10'd117};
ram[11786] = {9'd87,-10'd114};
ram[11787] = {9'd90,-10'd110};
ram[11788] = {9'd93,-10'd107};
ram[11789] = {9'd96,-10'd104};
ram[11790] = {9'd99,-10'd101};
ram[11791] = {-9'd98,-10'd98};
ram[11792] = {-9'd95,-10'd95};
ram[11793] = {-9'd92,-10'd92};
ram[11794] = {-9'd88,-10'd88};
ram[11795] = {-9'd85,-10'd85};
ram[11796] = {-9'd82,-10'd82};
ram[11797] = {-9'd79,-10'd79};
ram[11798] = {-9'd76,-10'd76};
ram[11799] = {-9'd73,-10'd73};
ram[11800] = {-9'd70,-10'd70};
ram[11801] = {-9'd66,-10'd66};
ram[11802] = {-9'd63,-10'd63};
ram[11803] = {-9'd60,-10'd60};
ram[11804] = {-9'd57,-10'd57};
ram[11805] = {-9'd54,-10'd54};
ram[11806] = {-9'd51,-10'd51};
ram[11807] = {-9'd48,-10'd48};
ram[11808] = {-9'd44,-10'd44};
ram[11809] = {-9'd41,-10'd41};
ram[11810] = {-9'd38,-10'd38};
ram[11811] = {-9'd35,-10'd35};
ram[11812] = {-9'd32,-10'd32};
ram[11813] = {-9'd29,-10'd29};
ram[11814] = {-9'd26,-10'd26};
ram[11815] = {-9'd22,-10'd22};
ram[11816] = {-9'd19,-10'd19};
ram[11817] = {-9'd16,-10'd16};
ram[11818] = {-9'd13,-10'd13};
ram[11819] = {-9'd10,-10'd10};
ram[11820] = {-9'd7,-10'd7};
ram[11821] = {-9'd4,-10'd4};
ram[11822] = {9'd0,10'd0};
ram[11823] = {9'd3,10'd3};
ram[11824] = {9'd6,10'd6};
ram[11825] = {9'd9,10'd9};
ram[11826] = {9'd12,10'd12};
ram[11827] = {9'd15,10'd15};
ram[11828] = {9'd18,10'd18};
ram[11829] = {9'd21,10'd21};
ram[11830] = {9'd25,10'd25};
ram[11831] = {9'd28,10'd28};
ram[11832] = {9'd31,10'd31};
ram[11833] = {9'd34,10'd34};
ram[11834] = {9'd37,10'd37};
ram[11835] = {9'd40,10'd40};
ram[11836] = {9'd43,10'd43};
ram[11837] = {9'd47,10'd47};
ram[11838] = {9'd50,10'd50};
ram[11839] = {9'd53,10'd53};
ram[11840] = {9'd56,10'd56};
ram[11841] = {9'd59,10'd59};
ram[11842] = {9'd62,10'd62};
ram[11843] = {9'd65,10'd65};
ram[11844] = {9'd69,10'd69};
ram[11845] = {9'd72,10'd72};
ram[11846] = {9'd75,10'd75};
ram[11847] = {9'd78,10'd78};
ram[11848] = {9'd81,10'd81};
ram[11849] = {9'd84,10'd84};
ram[11850] = {9'd87,10'd87};
ram[11851] = {9'd91,10'd91};
ram[11852] = {9'd94,10'd94};
ram[11853] = {9'd97,10'd97};
ram[11854] = {-9'd100,10'd100};
ram[11855] = {-9'd97,10'd103};
ram[11856] = {-9'd94,10'd106};
ram[11857] = {-9'd91,10'd109};
ram[11858] = {-9'd88,10'd113};
ram[11859] = {-9'd85,10'd116};
ram[11860] = {-9'd81,10'd119};
ram[11861] = {-9'd78,10'd122};
ram[11862] = {-9'd75,10'd125};
ram[11863] = {-9'd72,10'd128};
ram[11864] = {-9'd69,10'd131};
ram[11865] = {-9'd66,10'd135};
ram[11866] = {-9'd63,10'd138};
ram[11867] = {-9'd59,10'd141};
ram[11868] = {-9'd56,10'd144};
ram[11869] = {-9'd53,10'd147};
ram[11870] = {-9'd50,10'd150};
ram[11871] = {-9'd47,10'd153};
ram[11872] = {-9'd44,10'd157};
ram[11873] = {-9'd41,10'd160};
ram[11874] = {-9'd37,10'd163};
ram[11875] = {-9'd34,10'd166};
ram[11876] = {-9'd31,10'd169};
ram[11877] = {-9'd28,10'd172};
ram[11878] = {-9'd25,10'd175};
ram[11879] = {-9'd22,10'd179};
ram[11880] = {-9'd19,10'd182};
ram[11881] = {-9'd15,10'd185};
ram[11882] = {-9'd12,10'd188};
ram[11883] = {-9'd9,10'd191};
ram[11884] = {-9'd6,10'd194};
ram[11885] = {-9'd3,10'd197};
ram[11886] = {9'd0,10'd201};
ram[11887] = {9'd3,10'd204};
ram[11888] = {9'd7,10'd207};
ram[11889] = {9'd10,10'd210};
ram[11890] = {9'd13,10'd213};
ram[11891] = {9'd16,10'd216};
ram[11892] = {9'd19,10'd219};
ram[11893] = {9'd22,10'd223};
ram[11894] = {9'd25,10'd226};
ram[11895] = {9'd29,10'd229};
ram[11896] = {9'd32,10'd232};
ram[11897] = {9'd35,10'd235};
ram[11898] = {9'd38,10'd238};
ram[11899] = {9'd41,10'd241};
ram[11900] = {9'd44,10'd245};
ram[11901] = {9'd47,10'd248};
ram[11902] = {9'd51,10'd251};
ram[11903] = {9'd54,10'd254};
ram[11904] = {9'd54,10'd254};
ram[11905] = {9'd57,10'd257};
ram[11906] = {9'd60,10'd260};
ram[11907] = {9'd63,10'd263};
ram[11908] = {9'd66,10'd267};
ram[11909] = {9'd69,10'd270};
ram[11910] = {9'd73,10'd273};
ram[11911] = {9'd76,10'd276};
ram[11912] = {9'd79,10'd279};
ram[11913] = {9'd82,10'd282};
ram[11914] = {9'd85,10'd285};
ram[11915] = {9'd88,10'd289};
ram[11916] = {9'd91,10'd292};
ram[11917] = {9'd95,10'd295};
ram[11918] = {9'd98,10'd298};
ram[11919] = {-9'd99,10'd301};
ram[11920] = {-9'd96,10'd304};
ram[11921] = {-9'd93,10'd307};
ram[11922] = {-9'd90,10'd311};
ram[11923] = {-9'd87,10'd314};
ram[11924] = {-9'd84,10'd317};
ram[11925] = {-9'd81,10'd320};
ram[11926] = {-9'd77,10'd323};
ram[11927] = {-9'd74,10'd326};
ram[11928] = {-9'd71,10'd329};
ram[11929] = {-9'd68,10'd333};
ram[11930] = {-9'd65,10'd336};
ram[11931] = {-9'd62,10'd339};
ram[11932] = {-9'd59,10'd342};
ram[11933] = {-9'd55,10'd345};
ram[11934] = {-9'd52,10'd348};
ram[11935] = {-9'd49,10'd351};
ram[11936] = {-9'd46,10'd354};
ram[11937] = {-9'd43,10'd358};
ram[11938] = {-9'd40,10'd361};
ram[11939] = {-9'd37,10'd364};
ram[11940] = {-9'd33,10'd367};
ram[11941] = {-9'd30,10'd370};
ram[11942] = {-9'd27,10'd373};
ram[11943] = {-9'd24,10'd376};
ram[11944] = {-9'd21,10'd380};
ram[11945] = {-9'd18,10'd383};
ram[11946] = {-9'd15,10'd386};
ram[11947] = {-9'd11,10'd389};
ram[11948] = {-9'd8,10'd392};
ram[11949] = {-9'd5,10'd395};
ram[11950] = {-9'd2,10'd398};
ram[11951] = {9'd1,-10'd399};
ram[11952] = {9'd4,-10'd396};
ram[11953] = {9'd7,-10'd393};
ram[11954] = {9'd10,-10'd390};
ram[11955] = {9'd14,-10'd387};
ram[11956] = {9'd17,-10'd384};
ram[11957] = {9'd20,-10'd381};
ram[11958] = {9'd23,-10'd377};
ram[11959] = {9'd26,-10'd374};
ram[11960] = {9'd29,-10'd371};
ram[11961] = {9'd32,-10'd368};
ram[11962] = {9'd36,-10'd365};
ram[11963] = {9'd39,-10'd362};
ram[11964] = {9'd42,-10'd359};
ram[11965] = {9'd45,-10'd355};
ram[11966] = {9'd48,-10'd352};
ram[11967] = {9'd51,-10'd349};
ram[11968] = {9'd54,-10'd346};
ram[11969] = {9'd58,-10'd343};
ram[11970] = {9'd61,-10'd340};
ram[11971] = {9'd64,-10'd337};
ram[11972] = {9'd67,-10'd334};
ram[11973] = {9'd70,-10'd330};
ram[11974] = {9'd73,-10'd327};
ram[11975] = {9'd76,-10'd324};
ram[11976] = {9'd80,-10'd321};
ram[11977] = {9'd83,-10'd318};
ram[11978] = {9'd86,-10'd315};
ram[11979] = {9'd89,-10'd312};
ram[11980] = {9'd92,-10'd308};
ram[11981] = {9'd95,-10'd305};
ram[11982] = {9'd98,-10'd302};
ram[11983] = {-9'd99,-10'd299};
ram[11984] = {-9'd96,-10'd296};
ram[11985] = {-9'd92,-10'd293};
ram[11986] = {-9'd89,-10'd290};
ram[11987] = {-9'd86,-10'd286};
ram[11988] = {-9'd83,-10'd283};
ram[11989] = {-9'd80,-10'd280};
ram[11990] = {-9'd77,-10'd277};
ram[11991] = {-9'd74,-10'd274};
ram[11992] = {-9'd70,-10'd271};
ram[11993] = {-9'd67,-10'd268};
ram[11994] = {-9'd64,-10'd264};
ram[11995] = {-9'd61,-10'd261};
ram[11996] = {-9'd58,-10'd258};
ram[11997] = {-9'd55,-10'd255};
ram[11998] = {-9'd52,-10'd252};
ram[11999] = {-9'd48,-10'd249};
ram[12000] = {-9'd45,-10'd246};
ram[12001] = {-9'd42,-10'd242};
ram[12002] = {-9'd39,-10'd239};
ram[12003] = {-9'd36,-10'd236};
ram[12004] = {-9'd33,-10'd233};
ram[12005] = {-9'd30,-10'd230};
ram[12006] = {-9'd26,-10'd227};
ram[12007] = {-9'd23,-10'd224};
ram[12008] = {-9'd20,-10'd220};
ram[12009] = {-9'd17,-10'd217};
ram[12010] = {-9'd14,-10'd214};
ram[12011] = {-9'd11,-10'd211};
ram[12012] = {-9'd8,-10'd208};
ram[12013] = {-9'd4,-10'd205};
ram[12014] = {-9'd1,-10'd202};
ram[12015] = {9'd2,-10'd198};
ram[12016] = {9'd5,-10'd195};
ram[12017] = {9'd8,-10'd192};
ram[12018] = {9'd11,-10'd189};
ram[12019] = {9'd14,-10'd186};
ram[12020] = {9'd18,-10'd183};
ram[12021] = {9'd21,-10'd180};
ram[12022] = {9'd24,-10'd176};
ram[12023] = {9'd27,-10'd173};
ram[12024] = {9'd30,-10'd170};
ram[12025] = {9'd33,-10'd167};
ram[12026] = {9'd36,-10'd164};
ram[12027] = {9'd40,-10'd161};
ram[12028] = {9'd43,-10'd158};
ram[12029] = {9'd46,-10'd154};
ram[12030] = {9'd49,-10'd151};
ram[12031] = {9'd52,-10'd148};
ram[12032] = {9'd52,-10'd148};
ram[12033] = {9'd55,-10'd145};
ram[12034] = {9'd58,-10'd142};
ram[12035] = {9'd62,-10'd139};
ram[12036] = {9'd65,-10'd136};
ram[12037] = {9'd68,-10'd132};
ram[12038] = {9'd71,-10'd129};
ram[12039] = {9'd74,-10'd126};
ram[12040] = {9'd77,-10'd123};
ram[12041] = {9'd80,-10'd120};
ram[12042] = {9'd84,-10'd117};
ram[12043] = {9'd87,-10'd114};
ram[12044] = {9'd90,-10'd110};
ram[12045] = {9'd93,-10'd107};
ram[12046] = {9'd96,-10'd104};
ram[12047] = {9'd99,-10'd101};
ram[12048] = {-9'd98,-10'd98};
ram[12049] = {-9'd95,-10'd95};
ram[12050] = {-9'd92,-10'd92};
ram[12051] = {-9'd88,-10'd88};
ram[12052] = {-9'd85,-10'd85};
ram[12053] = {-9'd82,-10'd82};
ram[12054] = {-9'd79,-10'd79};
ram[12055] = {-9'd76,-10'd76};
ram[12056] = {-9'd73,-10'd73};
ram[12057] = {-9'd70,-10'd70};
ram[12058] = {-9'd66,-10'd66};
ram[12059] = {-9'd63,-10'd63};
ram[12060] = {-9'd60,-10'd60};
ram[12061] = {-9'd57,-10'd57};
ram[12062] = {-9'd54,-10'd54};
ram[12063] = {-9'd51,-10'd51};
ram[12064] = {-9'd48,-10'd48};
ram[12065] = {-9'd44,-10'd44};
ram[12066] = {-9'd41,-10'd41};
ram[12067] = {-9'd38,-10'd38};
ram[12068] = {-9'd35,-10'd35};
ram[12069] = {-9'd32,-10'd32};
ram[12070] = {-9'd29,-10'd29};
ram[12071] = {-9'd26,-10'd26};
ram[12072] = {-9'd22,-10'd22};
ram[12073] = {-9'd19,-10'd19};
ram[12074] = {-9'd16,-10'd16};
ram[12075] = {-9'd13,-10'd13};
ram[12076] = {-9'd10,-10'd10};
ram[12077] = {-9'd7,-10'd7};
ram[12078] = {-9'd4,-10'd4};
ram[12079] = {9'd0,10'd0};
ram[12080] = {9'd3,10'd3};
ram[12081] = {9'd6,10'd6};
ram[12082] = {9'd9,10'd9};
ram[12083] = {9'd12,10'd12};
ram[12084] = {9'd15,10'd15};
ram[12085] = {9'd18,10'd18};
ram[12086] = {9'd21,10'd21};
ram[12087] = {9'd25,10'd25};
ram[12088] = {9'd28,10'd28};
ram[12089] = {9'd31,10'd31};
ram[12090] = {9'd34,10'd34};
ram[12091] = {9'd37,10'd37};
ram[12092] = {9'd40,10'd40};
ram[12093] = {9'd43,10'd43};
ram[12094] = {9'd47,10'd47};
ram[12095] = {9'd50,10'd50};
ram[12096] = {9'd53,10'd53};
ram[12097] = {9'd56,10'd56};
ram[12098] = {9'd59,10'd59};
ram[12099] = {9'd62,10'd62};
ram[12100] = {9'd65,10'd65};
ram[12101] = {9'd69,10'd69};
ram[12102] = {9'd72,10'd72};
ram[12103] = {9'd75,10'd75};
ram[12104] = {9'd78,10'd78};
ram[12105] = {9'd81,10'd81};
ram[12106] = {9'd84,10'd84};
ram[12107] = {9'd87,10'd87};
ram[12108] = {9'd91,10'd91};
ram[12109] = {9'd94,10'd94};
ram[12110] = {9'd97,10'd97};
ram[12111] = {-9'd100,10'd100};
ram[12112] = {-9'd97,10'd103};
ram[12113] = {-9'd94,10'd106};
ram[12114] = {-9'd91,10'd109};
ram[12115] = {-9'd88,10'd113};
ram[12116] = {-9'd85,10'd116};
ram[12117] = {-9'd81,10'd119};
ram[12118] = {-9'd78,10'd122};
ram[12119] = {-9'd75,10'd125};
ram[12120] = {-9'd72,10'd128};
ram[12121] = {-9'd69,10'd131};
ram[12122] = {-9'd66,10'd135};
ram[12123] = {-9'd63,10'd138};
ram[12124] = {-9'd59,10'd141};
ram[12125] = {-9'd56,10'd144};
ram[12126] = {-9'd53,10'd147};
ram[12127] = {-9'd50,10'd150};
ram[12128] = {-9'd47,10'd153};
ram[12129] = {-9'd44,10'd157};
ram[12130] = {-9'd41,10'd160};
ram[12131] = {-9'd37,10'd163};
ram[12132] = {-9'd34,10'd166};
ram[12133] = {-9'd31,10'd169};
ram[12134] = {-9'd28,10'd172};
ram[12135] = {-9'd25,10'd175};
ram[12136] = {-9'd22,10'd179};
ram[12137] = {-9'd19,10'd182};
ram[12138] = {-9'd15,10'd185};
ram[12139] = {-9'd12,10'd188};
ram[12140] = {-9'd9,10'd191};
ram[12141] = {-9'd6,10'd194};
ram[12142] = {-9'd3,10'd197};
ram[12143] = {9'd0,10'd201};
ram[12144] = {9'd3,10'd204};
ram[12145] = {9'd7,10'd207};
ram[12146] = {9'd10,10'd210};
ram[12147] = {9'd13,10'd213};
ram[12148] = {9'd16,10'd216};
ram[12149] = {9'd19,10'd219};
ram[12150] = {9'd22,10'd223};
ram[12151] = {9'd25,10'd226};
ram[12152] = {9'd29,10'd229};
ram[12153] = {9'd32,10'd232};
ram[12154] = {9'd35,10'd235};
ram[12155] = {9'd38,10'd238};
ram[12156] = {9'd41,10'd241};
ram[12157] = {9'd44,10'd245};
ram[12158] = {9'd47,10'd248};
ram[12159] = {9'd51,10'd251};
ram[12160] = {9'd51,10'd251};
ram[12161] = {9'd54,10'd254};
ram[12162] = {9'd57,10'd257};
ram[12163] = {9'd60,10'd260};
ram[12164] = {9'd63,10'd263};
ram[12165] = {9'd66,10'd267};
ram[12166] = {9'd69,10'd270};
ram[12167] = {9'd73,10'd273};
ram[12168] = {9'd76,10'd276};
ram[12169] = {9'd79,10'd279};
ram[12170] = {9'd82,10'd282};
ram[12171] = {9'd85,10'd285};
ram[12172] = {9'd88,10'd289};
ram[12173] = {9'd91,10'd292};
ram[12174] = {9'd95,10'd295};
ram[12175] = {9'd98,10'd298};
ram[12176] = {-9'd99,10'd301};
ram[12177] = {-9'd96,10'd304};
ram[12178] = {-9'd93,10'd307};
ram[12179] = {-9'd90,10'd311};
ram[12180] = {-9'd87,10'd314};
ram[12181] = {-9'd84,10'd317};
ram[12182] = {-9'd81,10'd320};
ram[12183] = {-9'd77,10'd323};
ram[12184] = {-9'd74,10'd326};
ram[12185] = {-9'd71,10'd329};
ram[12186] = {-9'd68,10'd333};
ram[12187] = {-9'd65,10'd336};
ram[12188] = {-9'd62,10'd339};
ram[12189] = {-9'd59,10'd342};
ram[12190] = {-9'd55,10'd345};
ram[12191] = {-9'd52,10'd348};
ram[12192] = {-9'd49,10'd351};
ram[12193] = {-9'd46,10'd354};
ram[12194] = {-9'd43,10'd358};
ram[12195] = {-9'd40,10'd361};
ram[12196] = {-9'd37,10'd364};
ram[12197] = {-9'd33,10'd367};
ram[12198] = {-9'd30,10'd370};
ram[12199] = {-9'd27,10'd373};
ram[12200] = {-9'd24,10'd376};
ram[12201] = {-9'd21,10'd380};
ram[12202] = {-9'd18,10'd383};
ram[12203] = {-9'd15,10'd386};
ram[12204] = {-9'd11,10'd389};
ram[12205] = {-9'd8,10'd392};
ram[12206] = {-9'd5,10'd395};
ram[12207] = {-9'd2,10'd398};
ram[12208] = {9'd1,-10'd399};
ram[12209] = {9'd4,-10'd396};
ram[12210] = {9'd7,-10'd393};
ram[12211] = {9'd10,-10'd390};
ram[12212] = {9'd14,-10'd387};
ram[12213] = {9'd17,-10'd384};
ram[12214] = {9'd20,-10'd381};
ram[12215] = {9'd23,-10'd377};
ram[12216] = {9'd26,-10'd374};
ram[12217] = {9'd29,-10'd371};
ram[12218] = {9'd32,-10'd368};
ram[12219] = {9'd36,-10'd365};
ram[12220] = {9'd39,-10'd362};
ram[12221] = {9'd42,-10'd359};
ram[12222] = {9'd45,-10'd355};
ram[12223] = {9'd48,-10'd352};
ram[12224] = {9'd51,-10'd349};
ram[12225] = {9'd54,-10'd346};
ram[12226] = {9'd58,-10'd343};
ram[12227] = {9'd61,-10'd340};
ram[12228] = {9'd64,-10'd337};
ram[12229] = {9'd67,-10'd334};
ram[12230] = {9'd70,-10'd330};
ram[12231] = {9'd73,-10'd327};
ram[12232] = {9'd76,-10'd324};
ram[12233] = {9'd80,-10'd321};
ram[12234] = {9'd83,-10'd318};
ram[12235] = {9'd86,-10'd315};
ram[12236] = {9'd89,-10'd312};
ram[12237] = {9'd92,-10'd308};
ram[12238] = {9'd95,-10'd305};
ram[12239] = {9'd98,-10'd302};
ram[12240] = {-9'd99,-10'd299};
ram[12241] = {-9'd96,-10'd296};
ram[12242] = {-9'd92,-10'd293};
ram[12243] = {-9'd89,-10'd290};
ram[12244] = {-9'd86,-10'd286};
ram[12245] = {-9'd83,-10'd283};
ram[12246] = {-9'd80,-10'd280};
ram[12247] = {-9'd77,-10'd277};
ram[12248] = {-9'd74,-10'd274};
ram[12249] = {-9'd70,-10'd271};
ram[12250] = {-9'd67,-10'd268};
ram[12251] = {-9'd64,-10'd264};
ram[12252] = {-9'd61,-10'd261};
ram[12253] = {-9'd58,-10'd258};
ram[12254] = {-9'd55,-10'd255};
ram[12255] = {-9'd52,-10'd252};
ram[12256] = {-9'd48,-10'd249};
ram[12257] = {-9'd45,-10'd246};
ram[12258] = {-9'd42,-10'd242};
ram[12259] = {-9'd39,-10'd239};
ram[12260] = {-9'd36,-10'd236};
ram[12261] = {-9'd33,-10'd233};
ram[12262] = {-9'd30,-10'd230};
ram[12263] = {-9'd26,-10'd227};
ram[12264] = {-9'd23,-10'd224};
ram[12265] = {-9'd20,-10'd220};
ram[12266] = {-9'd17,-10'd217};
ram[12267] = {-9'd14,-10'd214};
ram[12268] = {-9'd11,-10'd211};
ram[12269] = {-9'd8,-10'd208};
ram[12270] = {-9'd4,-10'd205};
ram[12271] = {-9'd1,-10'd202};
ram[12272] = {9'd2,-10'd198};
ram[12273] = {9'd5,-10'd195};
ram[12274] = {9'd8,-10'd192};
ram[12275] = {9'd11,-10'd189};
ram[12276] = {9'd14,-10'd186};
ram[12277] = {9'd18,-10'd183};
ram[12278] = {9'd21,-10'd180};
ram[12279] = {9'd24,-10'd176};
ram[12280] = {9'd27,-10'd173};
ram[12281] = {9'd30,-10'd170};
ram[12282] = {9'd33,-10'd167};
ram[12283] = {9'd36,-10'd164};
ram[12284] = {9'd40,-10'd161};
ram[12285] = {9'd43,-10'd158};
ram[12286] = {9'd46,-10'd154};
ram[12287] = {9'd49,-10'd151};
ram[12288] = {9'd49,-10'd151};
ram[12289] = {9'd52,-10'd148};
ram[12290] = {9'd55,-10'd145};
ram[12291] = {9'd58,-10'd142};
ram[12292] = {9'd62,-10'd139};
ram[12293] = {9'd65,-10'd136};
ram[12294] = {9'd68,-10'd132};
ram[12295] = {9'd71,-10'd129};
ram[12296] = {9'd74,-10'd126};
ram[12297] = {9'd77,-10'd123};
ram[12298] = {9'd80,-10'd120};
ram[12299] = {9'd84,-10'd117};
ram[12300] = {9'd87,-10'd114};
ram[12301] = {9'd90,-10'd110};
ram[12302] = {9'd93,-10'd107};
ram[12303] = {9'd96,-10'd104};
ram[12304] = {9'd99,-10'd101};
ram[12305] = {-9'd98,-10'd98};
ram[12306] = {-9'd95,-10'd95};
ram[12307] = {-9'd92,-10'd92};
ram[12308] = {-9'd88,-10'd88};
ram[12309] = {-9'd85,-10'd85};
ram[12310] = {-9'd82,-10'd82};
ram[12311] = {-9'd79,-10'd79};
ram[12312] = {-9'd76,-10'd76};
ram[12313] = {-9'd73,-10'd73};
ram[12314] = {-9'd70,-10'd70};
ram[12315] = {-9'd66,-10'd66};
ram[12316] = {-9'd63,-10'd63};
ram[12317] = {-9'd60,-10'd60};
ram[12318] = {-9'd57,-10'd57};
ram[12319] = {-9'd54,-10'd54};
ram[12320] = {-9'd51,-10'd51};
ram[12321] = {-9'd48,-10'd48};
ram[12322] = {-9'd44,-10'd44};
ram[12323] = {-9'd41,-10'd41};
ram[12324] = {-9'd38,-10'd38};
ram[12325] = {-9'd35,-10'd35};
ram[12326] = {-9'd32,-10'd32};
ram[12327] = {-9'd29,-10'd29};
ram[12328] = {-9'd26,-10'd26};
ram[12329] = {-9'd22,-10'd22};
ram[12330] = {-9'd19,-10'd19};
ram[12331] = {-9'd16,-10'd16};
ram[12332] = {-9'd13,-10'd13};
ram[12333] = {-9'd10,-10'd10};
ram[12334] = {-9'd7,-10'd7};
ram[12335] = {-9'd4,-10'd4};
ram[12336] = {9'd0,10'd0};
ram[12337] = {9'd3,10'd3};
ram[12338] = {9'd6,10'd6};
ram[12339] = {9'd9,10'd9};
ram[12340] = {9'd12,10'd12};
ram[12341] = {9'd15,10'd15};
ram[12342] = {9'd18,10'd18};
ram[12343] = {9'd21,10'd21};
ram[12344] = {9'd25,10'd25};
ram[12345] = {9'd28,10'd28};
ram[12346] = {9'd31,10'd31};
ram[12347] = {9'd34,10'd34};
ram[12348] = {9'd37,10'd37};
ram[12349] = {9'd40,10'd40};
ram[12350] = {9'd43,10'd43};
ram[12351] = {9'd47,10'd47};
ram[12352] = {9'd50,10'd50};
ram[12353] = {9'd53,10'd53};
ram[12354] = {9'd56,10'd56};
ram[12355] = {9'd59,10'd59};
ram[12356] = {9'd62,10'd62};
ram[12357] = {9'd65,10'd65};
ram[12358] = {9'd69,10'd69};
ram[12359] = {9'd72,10'd72};
ram[12360] = {9'd75,10'd75};
ram[12361] = {9'd78,10'd78};
ram[12362] = {9'd81,10'd81};
ram[12363] = {9'd84,10'd84};
ram[12364] = {9'd87,10'd87};
ram[12365] = {9'd91,10'd91};
ram[12366] = {9'd94,10'd94};
ram[12367] = {9'd97,10'd97};
ram[12368] = {-9'd100,10'd100};
ram[12369] = {-9'd97,10'd103};
ram[12370] = {-9'd94,10'd106};
ram[12371] = {-9'd91,10'd109};
ram[12372] = {-9'd88,10'd113};
ram[12373] = {-9'd85,10'd116};
ram[12374] = {-9'd81,10'd119};
ram[12375] = {-9'd78,10'd122};
ram[12376] = {-9'd75,10'd125};
ram[12377] = {-9'd72,10'd128};
ram[12378] = {-9'd69,10'd131};
ram[12379] = {-9'd66,10'd135};
ram[12380] = {-9'd63,10'd138};
ram[12381] = {-9'd59,10'd141};
ram[12382] = {-9'd56,10'd144};
ram[12383] = {-9'd53,10'd147};
ram[12384] = {-9'd50,10'd150};
ram[12385] = {-9'd47,10'd153};
ram[12386] = {-9'd44,10'd157};
ram[12387] = {-9'd41,10'd160};
ram[12388] = {-9'd37,10'd163};
ram[12389] = {-9'd34,10'd166};
ram[12390] = {-9'd31,10'd169};
ram[12391] = {-9'd28,10'd172};
ram[12392] = {-9'd25,10'd175};
ram[12393] = {-9'd22,10'd179};
ram[12394] = {-9'd19,10'd182};
ram[12395] = {-9'd15,10'd185};
ram[12396] = {-9'd12,10'd188};
ram[12397] = {-9'd9,10'd191};
ram[12398] = {-9'd6,10'd194};
ram[12399] = {-9'd3,10'd197};
ram[12400] = {9'd0,10'd201};
ram[12401] = {9'd3,10'd204};
ram[12402] = {9'd7,10'd207};
ram[12403] = {9'd10,10'd210};
ram[12404] = {9'd13,10'd213};
ram[12405] = {9'd16,10'd216};
ram[12406] = {9'd19,10'd219};
ram[12407] = {9'd22,10'd223};
ram[12408] = {9'd25,10'd226};
ram[12409] = {9'd29,10'd229};
ram[12410] = {9'd32,10'd232};
ram[12411] = {9'd35,10'd235};
ram[12412] = {9'd38,10'd238};
ram[12413] = {9'd41,10'd241};
ram[12414] = {9'd44,10'd245};
ram[12415] = {9'd47,10'd248};
ram[12416] = {9'd47,10'd248};
ram[12417] = {9'd51,10'd251};
ram[12418] = {9'd54,10'd254};
ram[12419] = {9'd57,10'd257};
ram[12420] = {9'd60,10'd260};
ram[12421] = {9'd63,10'd263};
ram[12422] = {9'd66,10'd267};
ram[12423] = {9'd69,10'd270};
ram[12424] = {9'd73,10'd273};
ram[12425] = {9'd76,10'd276};
ram[12426] = {9'd79,10'd279};
ram[12427] = {9'd82,10'd282};
ram[12428] = {9'd85,10'd285};
ram[12429] = {9'd88,10'd289};
ram[12430] = {9'd91,10'd292};
ram[12431] = {9'd95,10'd295};
ram[12432] = {9'd98,10'd298};
ram[12433] = {-9'd99,10'd301};
ram[12434] = {-9'd96,10'd304};
ram[12435] = {-9'd93,10'd307};
ram[12436] = {-9'd90,10'd311};
ram[12437] = {-9'd87,10'd314};
ram[12438] = {-9'd84,10'd317};
ram[12439] = {-9'd81,10'd320};
ram[12440] = {-9'd77,10'd323};
ram[12441] = {-9'd74,10'd326};
ram[12442] = {-9'd71,10'd329};
ram[12443] = {-9'd68,10'd333};
ram[12444] = {-9'd65,10'd336};
ram[12445] = {-9'd62,10'd339};
ram[12446] = {-9'd59,10'd342};
ram[12447] = {-9'd55,10'd345};
ram[12448] = {-9'd52,10'd348};
ram[12449] = {-9'd49,10'd351};
ram[12450] = {-9'd46,10'd354};
ram[12451] = {-9'd43,10'd358};
ram[12452] = {-9'd40,10'd361};
ram[12453] = {-9'd37,10'd364};
ram[12454] = {-9'd33,10'd367};
ram[12455] = {-9'd30,10'd370};
ram[12456] = {-9'd27,10'd373};
ram[12457] = {-9'd24,10'd376};
ram[12458] = {-9'd21,10'd380};
ram[12459] = {-9'd18,10'd383};
ram[12460] = {-9'd15,10'd386};
ram[12461] = {-9'd11,10'd389};
ram[12462] = {-9'd8,10'd392};
ram[12463] = {-9'd5,10'd395};
ram[12464] = {-9'd2,10'd398};
ram[12465] = {9'd1,-10'd399};
ram[12466] = {9'd4,-10'd396};
ram[12467] = {9'd7,-10'd393};
ram[12468] = {9'd10,-10'd390};
ram[12469] = {9'd14,-10'd387};
ram[12470] = {9'd17,-10'd384};
ram[12471] = {9'd20,-10'd381};
ram[12472] = {9'd23,-10'd377};
ram[12473] = {9'd26,-10'd374};
ram[12474] = {9'd29,-10'd371};
ram[12475] = {9'd32,-10'd368};
ram[12476] = {9'd36,-10'd365};
ram[12477] = {9'd39,-10'd362};
ram[12478] = {9'd42,-10'd359};
ram[12479] = {9'd45,-10'd355};
ram[12480] = {9'd48,-10'd352};
ram[12481] = {9'd51,-10'd349};
ram[12482] = {9'd54,-10'd346};
ram[12483] = {9'd58,-10'd343};
ram[12484] = {9'd61,-10'd340};
ram[12485] = {9'd64,-10'd337};
ram[12486] = {9'd67,-10'd334};
ram[12487] = {9'd70,-10'd330};
ram[12488] = {9'd73,-10'd327};
ram[12489] = {9'd76,-10'd324};
ram[12490] = {9'd80,-10'd321};
ram[12491] = {9'd83,-10'd318};
ram[12492] = {9'd86,-10'd315};
ram[12493] = {9'd89,-10'd312};
ram[12494] = {9'd92,-10'd308};
ram[12495] = {9'd95,-10'd305};
ram[12496] = {9'd98,-10'd302};
ram[12497] = {-9'd99,-10'd299};
ram[12498] = {-9'd96,-10'd296};
ram[12499] = {-9'd92,-10'd293};
ram[12500] = {-9'd89,-10'd290};
ram[12501] = {-9'd86,-10'd286};
ram[12502] = {-9'd83,-10'd283};
ram[12503] = {-9'd80,-10'd280};
ram[12504] = {-9'd77,-10'd277};
ram[12505] = {-9'd74,-10'd274};
ram[12506] = {-9'd70,-10'd271};
ram[12507] = {-9'd67,-10'd268};
ram[12508] = {-9'd64,-10'd264};
ram[12509] = {-9'd61,-10'd261};
ram[12510] = {-9'd58,-10'd258};
ram[12511] = {-9'd55,-10'd255};
ram[12512] = {-9'd52,-10'd252};
ram[12513] = {-9'd48,-10'd249};
ram[12514] = {-9'd45,-10'd246};
ram[12515] = {-9'd42,-10'd242};
ram[12516] = {-9'd39,-10'd239};
ram[12517] = {-9'd36,-10'd236};
ram[12518] = {-9'd33,-10'd233};
ram[12519] = {-9'd30,-10'd230};
ram[12520] = {-9'd26,-10'd227};
ram[12521] = {-9'd23,-10'd224};
ram[12522] = {-9'd20,-10'd220};
ram[12523] = {-9'd17,-10'd217};
ram[12524] = {-9'd14,-10'd214};
ram[12525] = {-9'd11,-10'd211};
ram[12526] = {-9'd8,-10'd208};
ram[12527] = {-9'd4,-10'd205};
ram[12528] = {-9'd1,-10'd202};
ram[12529] = {9'd2,-10'd198};
ram[12530] = {9'd5,-10'd195};
ram[12531] = {9'd8,-10'd192};
ram[12532] = {9'd11,-10'd189};
ram[12533] = {9'd14,-10'd186};
ram[12534] = {9'd18,-10'd183};
ram[12535] = {9'd21,-10'd180};
ram[12536] = {9'd24,-10'd176};
ram[12537] = {9'd27,-10'd173};
ram[12538] = {9'd30,-10'd170};
ram[12539] = {9'd33,-10'd167};
ram[12540] = {9'd36,-10'd164};
ram[12541] = {9'd40,-10'd161};
ram[12542] = {9'd43,-10'd158};
ram[12543] = {9'd46,-10'd154};
ram[12544] = {9'd46,-10'd154};
ram[12545] = {9'd49,-10'd151};
ram[12546] = {9'd52,-10'd148};
ram[12547] = {9'd55,-10'd145};
ram[12548] = {9'd58,-10'd142};
ram[12549] = {9'd62,-10'd139};
ram[12550] = {9'd65,-10'd136};
ram[12551] = {9'd68,-10'd132};
ram[12552] = {9'd71,-10'd129};
ram[12553] = {9'd74,-10'd126};
ram[12554] = {9'd77,-10'd123};
ram[12555] = {9'd80,-10'd120};
ram[12556] = {9'd84,-10'd117};
ram[12557] = {9'd87,-10'd114};
ram[12558] = {9'd90,-10'd110};
ram[12559] = {9'd93,-10'd107};
ram[12560] = {9'd96,-10'd104};
ram[12561] = {9'd99,-10'd101};
ram[12562] = {-9'd98,-10'd98};
ram[12563] = {-9'd95,-10'd95};
ram[12564] = {-9'd92,-10'd92};
ram[12565] = {-9'd88,-10'd88};
ram[12566] = {-9'd85,-10'd85};
ram[12567] = {-9'd82,-10'd82};
ram[12568] = {-9'd79,-10'd79};
ram[12569] = {-9'd76,-10'd76};
ram[12570] = {-9'd73,-10'd73};
ram[12571] = {-9'd70,-10'd70};
ram[12572] = {-9'd66,-10'd66};
ram[12573] = {-9'd63,-10'd63};
ram[12574] = {-9'd60,-10'd60};
ram[12575] = {-9'd57,-10'd57};
ram[12576] = {-9'd54,-10'd54};
ram[12577] = {-9'd51,-10'd51};
ram[12578] = {-9'd48,-10'd48};
ram[12579] = {-9'd44,-10'd44};
ram[12580] = {-9'd41,-10'd41};
ram[12581] = {-9'd38,-10'd38};
ram[12582] = {-9'd35,-10'd35};
ram[12583] = {-9'd32,-10'd32};
ram[12584] = {-9'd29,-10'd29};
ram[12585] = {-9'd26,-10'd26};
ram[12586] = {-9'd22,-10'd22};
ram[12587] = {-9'd19,-10'd19};
ram[12588] = {-9'd16,-10'd16};
ram[12589] = {-9'd13,-10'd13};
ram[12590] = {-9'd10,-10'd10};
ram[12591] = {-9'd7,-10'd7};
ram[12592] = {-9'd4,-10'd4};
ram[12593] = {9'd0,10'd0};
ram[12594] = {9'd3,10'd3};
ram[12595] = {9'd6,10'd6};
ram[12596] = {9'd9,10'd9};
ram[12597] = {9'd12,10'd12};
ram[12598] = {9'd15,10'd15};
ram[12599] = {9'd18,10'd18};
ram[12600] = {9'd21,10'd21};
ram[12601] = {9'd25,10'd25};
ram[12602] = {9'd28,10'd28};
ram[12603] = {9'd31,10'd31};
ram[12604] = {9'd34,10'd34};
ram[12605] = {9'd37,10'd37};
ram[12606] = {9'd40,10'd40};
ram[12607] = {9'd43,10'd43};
ram[12608] = {9'd47,10'd47};
ram[12609] = {9'd50,10'd50};
ram[12610] = {9'd53,10'd53};
ram[12611] = {9'd56,10'd56};
ram[12612] = {9'd59,10'd59};
ram[12613] = {9'd62,10'd62};
ram[12614] = {9'd65,10'd65};
ram[12615] = {9'd69,10'd69};
ram[12616] = {9'd72,10'd72};
ram[12617] = {9'd75,10'd75};
ram[12618] = {9'd78,10'd78};
ram[12619] = {9'd81,10'd81};
ram[12620] = {9'd84,10'd84};
ram[12621] = {9'd87,10'd87};
ram[12622] = {9'd91,10'd91};
ram[12623] = {9'd94,10'd94};
ram[12624] = {9'd97,10'd97};
ram[12625] = {-9'd100,10'd100};
ram[12626] = {-9'd97,10'd103};
ram[12627] = {-9'd94,10'd106};
ram[12628] = {-9'd91,10'd109};
ram[12629] = {-9'd88,10'd113};
ram[12630] = {-9'd85,10'd116};
ram[12631] = {-9'd81,10'd119};
ram[12632] = {-9'd78,10'd122};
ram[12633] = {-9'd75,10'd125};
ram[12634] = {-9'd72,10'd128};
ram[12635] = {-9'd69,10'd131};
ram[12636] = {-9'd66,10'd135};
ram[12637] = {-9'd63,10'd138};
ram[12638] = {-9'd59,10'd141};
ram[12639] = {-9'd56,10'd144};
ram[12640] = {-9'd53,10'd147};
ram[12641] = {-9'd50,10'd150};
ram[12642] = {-9'd47,10'd153};
ram[12643] = {-9'd44,10'd157};
ram[12644] = {-9'd41,10'd160};
ram[12645] = {-9'd37,10'd163};
ram[12646] = {-9'd34,10'd166};
ram[12647] = {-9'd31,10'd169};
ram[12648] = {-9'd28,10'd172};
ram[12649] = {-9'd25,10'd175};
ram[12650] = {-9'd22,10'd179};
ram[12651] = {-9'd19,10'd182};
ram[12652] = {-9'd15,10'd185};
ram[12653] = {-9'd12,10'd188};
ram[12654] = {-9'd9,10'd191};
ram[12655] = {-9'd6,10'd194};
ram[12656] = {-9'd3,10'd197};
ram[12657] = {9'd0,10'd201};
ram[12658] = {9'd3,10'd204};
ram[12659] = {9'd7,10'd207};
ram[12660] = {9'd10,10'd210};
ram[12661] = {9'd13,10'd213};
ram[12662] = {9'd16,10'd216};
ram[12663] = {9'd19,10'd219};
ram[12664] = {9'd22,10'd223};
ram[12665] = {9'd25,10'd226};
ram[12666] = {9'd29,10'd229};
ram[12667] = {9'd32,10'd232};
ram[12668] = {9'd35,10'd235};
ram[12669] = {9'd38,10'd238};
ram[12670] = {9'd41,10'd241};
ram[12671] = {9'd44,10'd245};
ram[12672] = {9'd44,10'd245};
ram[12673] = {9'd47,10'd248};
ram[12674] = {9'd51,10'd251};
ram[12675] = {9'd54,10'd254};
ram[12676] = {9'd57,10'd257};
ram[12677] = {9'd60,10'd260};
ram[12678] = {9'd63,10'd263};
ram[12679] = {9'd66,10'd267};
ram[12680] = {9'd69,10'd270};
ram[12681] = {9'd73,10'd273};
ram[12682] = {9'd76,10'd276};
ram[12683] = {9'd79,10'd279};
ram[12684] = {9'd82,10'd282};
ram[12685] = {9'd85,10'd285};
ram[12686] = {9'd88,10'd289};
ram[12687] = {9'd91,10'd292};
ram[12688] = {9'd95,10'd295};
ram[12689] = {9'd98,10'd298};
ram[12690] = {-9'd99,10'd301};
ram[12691] = {-9'd96,10'd304};
ram[12692] = {-9'd93,10'd307};
ram[12693] = {-9'd90,10'd311};
ram[12694] = {-9'd87,10'd314};
ram[12695] = {-9'd84,10'd317};
ram[12696] = {-9'd81,10'd320};
ram[12697] = {-9'd77,10'd323};
ram[12698] = {-9'd74,10'd326};
ram[12699] = {-9'd71,10'd329};
ram[12700] = {-9'd68,10'd333};
ram[12701] = {-9'd65,10'd336};
ram[12702] = {-9'd62,10'd339};
ram[12703] = {-9'd59,10'd342};
ram[12704] = {-9'd55,10'd345};
ram[12705] = {-9'd52,10'd348};
ram[12706] = {-9'd49,10'd351};
ram[12707] = {-9'd46,10'd354};
ram[12708] = {-9'd43,10'd358};
ram[12709] = {-9'd40,10'd361};
ram[12710] = {-9'd37,10'd364};
ram[12711] = {-9'd33,10'd367};
ram[12712] = {-9'd30,10'd370};
ram[12713] = {-9'd27,10'd373};
ram[12714] = {-9'd24,10'd376};
ram[12715] = {-9'd21,10'd380};
ram[12716] = {-9'd18,10'd383};
ram[12717] = {-9'd15,10'd386};
ram[12718] = {-9'd11,10'd389};
ram[12719] = {-9'd8,10'd392};
ram[12720] = {-9'd5,10'd395};
ram[12721] = {-9'd2,10'd398};
ram[12722] = {9'd1,-10'd399};
ram[12723] = {9'd4,-10'd396};
ram[12724] = {9'd7,-10'd393};
ram[12725] = {9'd10,-10'd390};
ram[12726] = {9'd14,-10'd387};
ram[12727] = {9'd17,-10'd384};
ram[12728] = {9'd20,-10'd381};
ram[12729] = {9'd23,-10'd377};
ram[12730] = {9'd26,-10'd374};
ram[12731] = {9'd29,-10'd371};
ram[12732] = {9'd32,-10'd368};
ram[12733] = {9'd36,-10'd365};
ram[12734] = {9'd39,-10'd362};
ram[12735] = {9'd42,-10'd359};
ram[12736] = {9'd45,-10'd355};
ram[12737] = {9'd48,-10'd352};
ram[12738] = {9'd51,-10'd349};
ram[12739] = {9'd54,-10'd346};
ram[12740] = {9'd58,-10'd343};
ram[12741] = {9'd61,-10'd340};
ram[12742] = {9'd64,-10'd337};
ram[12743] = {9'd67,-10'd334};
ram[12744] = {9'd70,-10'd330};
ram[12745] = {9'd73,-10'd327};
ram[12746] = {9'd76,-10'd324};
ram[12747] = {9'd80,-10'd321};
ram[12748] = {9'd83,-10'd318};
ram[12749] = {9'd86,-10'd315};
ram[12750] = {9'd89,-10'd312};
ram[12751] = {9'd92,-10'd308};
ram[12752] = {9'd95,-10'd305};
ram[12753] = {9'd98,-10'd302};
ram[12754] = {-9'd99,-10'd299};
ram[12755] = {-9'd96,-10'd296};
ram[12756] = {-9'd92,-10'd293};
ram[12757] = {-9'd89,-10'd290};
ram[12758] = {-9'd86,-10'd286};
ram[12759] = {-9'd83,-10'd283};
ram[12760] = {-9'd80,-10'd280};
ram[12761] = {-9'd77,-10'd277};
ram[12762] = {-9'd74,-10'd274};
ram[12763] = {-9'd70,-10'd271};
ram[12764] = {-9'd67,-10'd268};
ram[12765] = {-9'd64,-10'd264};
ram[12766] = {-9'd61,-10'd261};
ram[12767] = {-9'd58,-10'd258};
ram[12768] = {-9'd55,-10'd255};
ram[12769] = {-9'd52,-10'd252};
ram[12770] = {-9'd48,-10'd249};
ram[12771] = {-9'd45,-10'd246};
ram[12772] = {-9'd42,-10'd242};
ram[12773] = {-9'd39,-10'd239};
ram[12774] = {-9'd36,-10'd236};
ram[12775] = {-9'd33,-10'd233};
ram[12776] = {-9'd30,-10'd230};
ram[12777] = {-9'd26,-10'd227};
ram[12778] = {-9'd23,-10'd224};
ram[12779] = {-9'd20,-10'd220};
ram[12780] = {-9'd17,-10'd217};
ram[12781] = {-9'd14,-10'd214};
ram[12782] = {-9'd11,-10'd211};
ram[12783] = {-9'd8,-10'd208};
ram[12784] = {-9'd4,-10'd205};
ram[12785] = {-9'd1,-10'd202};
ram[12786] = {9'd2,-10'd198};
ram[12787] = {9'd5,-10'd195};
ram[12788] = {9'd8,-10'd192};
ram[12789] = {9'd11,-10'd189};
ram[12790] = {9'd14,-10'd186};
ram[12791] = {9'd18,-10'd183};
ram[12792] = {9'd21,-10'd180};
ram[12793] = {9'd24,-10'd176};
ram[12794] = {9'd27,-10'd173};
ram[12795] = {9'd30,-10'd170};
ram[12796] = {9'd33,-10'd167};
ram[12797] = {9'd36,-10'd164};
ram[12798] = {9'd40,-10'd161};
ram[12799] = {9'd43,-10'd158};
ram[12800] = {9'd43,-10'd158};
ram[12801] = {9'd46,-10'd154};
ram[12802] = {9'd49,-10'd151};
ram[12803] = {9'd52,-10'd148};
ram[12804] = {9'd55,-10'd145};
ram[12805] = {9'd58,-10'd142};
ram[12806] = {9'd62,-10'd139};
ram[12807] = {9'd65,-10'd136};
ram[12808] = {9'd68,-10'd132};
ram[12809] = {9'd71,-10'd129};
ram[12810] = {9'd74,-10'd126};
ram[12811] = {9'd77,-10'd123};
ram[12812] = {9'd80,-10'd120};
ram[12813] = {9'd84,-10'd117};
ram[12814] = {9'd87,-10'd114};
ram[12815] = {9'd90,-10'd110};
ram[12816] = {9'd93,-10'd107};
ram[12817] = {9'd96,-10'd104};
ram[12818] = {9'd99,-10'd101};
ram[12819] = {-9'd98,-10'd98};
ram[12820] = {-9'd95,-10'd95};
ram[12821] = {-9'd92,-10'd92};
ram[12822] = {-9'd88,-10'd88};
ram[12823] = {-9'd85,-10'd85};
ram[12824] = {-9'd82,-10'd82};
ram[12825] = {-9'd79,-10'd79};
ram[12826] = {-9'd76,-10'd76};
ram[12827] = {-9'd73,-10'd73};
ram[12828] = {-9'd70,-10'd70};
ram[12829] = {-9'd66,-10'd66};
ram[12830] = {-9'd63,-10'd63};
ram[12831] = {-9'd60,-10'd60};
ram[12832] = {-9'd57,-10'd57};
ram[12833] = {-9'd54,-10'd54};
ram[12834] = {-9'd51,-10'd51};
ram[12835] = {-9'd48,-10'd48};
ram[12836] = {-9'd44,-10'd44};
ram[12837] = {-9'd41,-10'd41};
ram[12838] = {-9'd38,-10'd38};
ram[12839] = {-9'd35,-10'd35};
ram[12840] = {-9'd32,-10'd32};
ram[12841] = {-9'd29,-10'd29};
ram[12842] = {-9'd26,-10'd26};
ram[12843] = {-9'd22,-10'd22};
ram[12844] = {-9'd19,-10'd19};
ram[12845] = {-9'd16,-10'd16};
ram[12846] = {-9'd13,-10'd13};
ram[12847] = {-9'd10,-10'd10};
ram[12848] = {-9'd7,-10'd7};
ram[12849] = {-9'd4,-10'd4};
ram[12850] = {9'd0,10'd0};
ram[12851] = {9'd3,10'd3};
ram[12852] = {9'd6,10'd6};
ram[12853] = {9'd9,10'd9};
ram[12854] = {9'd12,10'd12};
ram[12855] = {9'd15,10'd15};
ram[12856] = {9'd18,10'd18};
ram[12857] = {9'd21,10'd21};
ram[12858] = {9'd25,10'd25};
ram[12859] = {9'd28,10'd28};
ram[12860] = {9'd31,10'd31};
ram[12861] = {9'd34,10'd34};
ram[12862] = {9'd37,10'd37};
ram[12863] = {9'd40,10'd40};
ram[12864] = {9'd43,10'd43};
ram[12865] = {9'd47,10'd47};
ram[12866] = {9'd50,10'd50};
ram[12867] = {9'd53,10'd53};
ram[12868] = {9'd56,10'd56};
ram[12869] = {9'd59,10'd59};
ram[12870] = {9'd62,10'd62};
ram[12871] = {9'd65,10'd65};
ram[12872] = {9'd69,10'd69};
ram[12873] = {9'd72,10'd72};
ram[12874] = {9'd75,10'd75};
ram[12875] = {9'd78,10'd78};
ram[12876] = {9'd81,10'd81};
ram[12877] = {9'd84,10'd84};
ram[12878] = {9'd87,10'd87};
ram[12879] = {9'd91,10'd91};
ram[12880] = {9'd94,10'd94};
ram[12881] = {9'd97,10'd97};
ram[12882] = {-9'd100,10'd100};
ram[12883] = {-9'd97,10'd103};
ram[12884] = {-9'd94,10'd106};
ram[12885] = {-9'd91,10'd109};
ram[12886] = {-9'd88,10'd113};
ram[12887] = {-9'd85,10'd116};
ram[12888] = {-9'd81,10'd119};
ram[12889] = {-9'd78,10'd122};
ram[12890] = {-9'd75,10'd125};
ram[12891] = {-9'd72,10'd128};
ram[12892] = {-9'd69,10'd131};
ram[12893] = {-9'd66,10'd135};
ram[12894] = {-9'd63,10'd138};
ram[12895] = {-9'd59,10'd141};
ram[12896] = {-9'd56,10'd144};
ram[12897] = {-9'd53,10'd147};
ram[12898] = {-9'd50,10'd150};
ram[12899] = {-9'd47,10'd153};
ram[12900] = {-9'd44,10'd157};
ram[12901] = {-9'd41,10'd160};
ram[12902] = {-9'd37,10'd163};
ram[12903] = {-9'd34,10'd166};
ram[12904] = {-9'd31,10'd169};
ram[12905] = {-9'd28,10'd172};
ram[12906] = {-9'd25,10'd175};
ram[12907] = {-9'd22,10'd179};
ram[12908] = {-9'd19,10'd182};
ram[12909] = {-9'd15,10'd185};
ram[12910] = {-9'd12,10'd188};
ram[12911] = {-9'd9,10'd191};
ram[12912] = {-9'd6,10'd194};
ram[12913] = {-9'd3,10'd197};
ram[12914] = {9'd0,10'd201};
ram[12915] = {9'd3,10'd204};
ram[12916] = {9'd7,10'd207};
ram[12917] = {9'd10,10'd210};
ram[12918] = {9'd13,10'd213};
ram[12919] = {9'd16,10'd216};
ram[12920] = {9'd19,10'd219};
ram[12921] = {9'd22,10'd223};
ram[12922] = {9'd25,10'd226};
ram[12923] = {9'd29,10'd229};
ram[12924] = {9'd32,10'd232};
ram[12925] = {9'd35,10'd235};
ram[12926] = {9'd38,10'd238};
ram[12927] = {9'd41,10'd241};
ram[12928] = {9'd41,10'd241};
ram[12929] = {9'd44,10'd245};
ram[12930] = {9'd47,10'd248};
ram[12931] = {9'd51,10'd251};
ram[12932] = {9'd54,10'd254};
ram[12933] = {9'd57,10'd257};
ram[12934] = {9'd60,10'd260};
ram[12935] = {9'd63,10'd263};
ram[12936] = {9'd66,10'd267};
ram[12937] = {9'd69,10'd270};
ram[12938] = {9'd73,10'd273};
ram[12939] = {9'd76,10'd276};
ram[12940] = {9'd79,10'd279};
ram[12941] = {9'd82,10'd282};
ram[12942] = {9'd85,10'd285};
ram[12943] = {9'd88,10'd289};
ram[12944] = {9'd91,10'd292};
ram[12945] = {9'd95,10'd295};
ram[12946] = {9'd98,10'd298};
ram[12947] = {-9'd99,10'd301};
ram[12948] = {-9'd96,10'd304};
ram[12949] = {-9'd93,10'd307};
ram[12950] = {-9'd90,10'd311};
ram[12951] = {-9'd87,10'd314};
ram[12952] = {-9'd84,10'd317};
ram[12953] = {-9'd81,10'd320};
ram[12954] = {-9'd77,10'd323};
ram[12955] = {-9'd74,10'd326};
ram[12956] = {-9'd71,10'd329};
ram[12957] = {-9'd68,10'd333};
ram[12958] = {-9'd65,10'd336};
ram[12959] = {-9'd62,10'd339};
ram[12960] = {-9'd59,10'd342};
ram[12961] = {-9'd55,10'd345};
ram[12962] = {-9'd52,10'd348};
ram[12963] = {-9'd49,10'd351};
ram[12964] = {-9'd46,10'd354};
ram[12965] = {-9'd43,10'd358};
ram[12966] = {-9'd40,10'd361};
ram[12967] = {-9'd37,10'd364};
ram[12968] = {-9'd33,10'd367};
ram[12969] = {-9'd30,10'd370};
ram[12970] = {-9'd27,10'd373};
ram[12971] = {-9'd24,10'd376};
ram[12972] = {-9'd21,10'd380};
ram[12973] = {-9'd18,10'd383};
ram[12974] = {-9'd15,10'd386};
ram[12975] = {-9'd11,10'd389};
ram[12976] = {-9'd8,10'd392};
ram[12977] = {-9'd5,10'd395};
ram[12978] = {-9'd2,10'd398};
ram[12979] = {9'd1,-10'd399};
ram[12980] = {9'd4,-10'd396};
ram[12981] = {9'd7,-10'd393};
ram[12982] = {9'd10,-10'd390};
ram[12983] = {9'd14,-10'd387};
ram[12984] = {9'd17,-10'd384};
ram[12985] = {9'd20,-10'd381};
ram[12986] = {9'd23,-10'd377};
ram[12987] = {9'd26,-10'd374};
ram[12988] = {9'd29,-10'd371};
ram[12989] = {9'd32,-10'd368};
ram[12990] = {9'd36,-10'd365};
ram[12991] = {9'd39,-10'd362};
ram[12992] = {9'd42,-10'd359};
ram[12993] = {9'd45,-10'd355};
ram[12994] = {9'd48,-10'd352};
ram[12995] = {9'd51,-10'd349};
ram[12996] = {9'd54,-10'd346};
ram[12997] = {9'd58,-10'd343};
ram[12998] = {9'd61,-10'd340};
ram[12999] = {9'd64,-10'd337};
ram[13000] = {9'd67,-10'd334};
ram[13001] = {9'd70,-10'd330};
ram[13002] = {9'd73,-10'd327};
ram[13003] = {9'd76,-10'd324};
ram[13004] = {9'd80,-10'd321};
ram[13005] = {9'd83,-10'd318};
ram[13006] = {9'd86,-10'd315};
ram[13007] = {9'd89,-10'd312};
ram[13008] = {9'd92,-10'd308};
ram[13009] = {9'd95,-10'd305};
ram[13010] = {9'd98,-10'd302};
ram[13011] = {-9'd99,-10'd299};
ram[13012] = {-9'd96,-10'd296};
ram[13013] = {-9'd92,-10'd293};
ram[13014] = {-9'd89,-10'd290};
ram[13015] = {-9'd86,-10'd286};
ram[13016] = {-9'd83,-10'd283};
ram[13017] = {-9'd80,-10'd280};
ram[13018] = {-9'd77,-10'd277};
ram[13019] = {-9'd74,-10'd274};
ram[13020] = {-9'd70,-10'd271};
ram[13021] = {-9'd67,-10'd268};
ram[13022] = {-9'd64,-10'd264};
ram[13023] = {-9'd61,-10'd261};
ram[13024] = {-9'd58,-10'd258};
ram[13025] = {-9'd55,-10'd255};
ram[13026] = {-9'd52,-10'd252};
ram[13027] = {-9'd48,-10'd249};
ram[13028] = {-9'd45,-10'd246};
ram[13029] = {-9'd42,-10'd242};
ram[13030] = {-9'd39,-10'd239};
ram[13031] = {-9'd36,-10'd236};
ram[13032] = {-9'd33,-10'd233};
ram[13033] = {-9'd30,-10'd230};
ram[13034] = {-9'd26,-10'd227};
ram[13035] = {-9'd23,-10'd224};
ram[13036] = {-9'd20,-10'd220};
ram[13037] = {-9'd17,-10'd217};
ram[13038] = {-9'd14,-10'd214};
ram[13039] = {-9'd11,-10'd211};
ram[13040] = {-9'd8,-10'd208};
ram[13041] = {-9'd4,-10'd205};
ram[13042] = {-9'd1,-10'd202};
ram[13043] = {9'd2,-10'd198};
ram[13044] = {9'd5,-10'd195};
ram[13045] = {9'd8,-10'd192};
ram[13046] = {9'd11,-10'd189};
ram[13047] = {9'd14,-10'd186};
ram[13048] = {9'd18,-10'd183};
ram[13049] = {9'd21,-10'd180};
ram[13050] = {9'd24,-10'd176};
ram[13051] = {9'd27,-10'd173};
ram[13052] = {9'd30,-10'd170};
ram[13053] = {9'd33,-10'd167};
ram[13054] = {9'd36,-10'd164};
ram[13055] = {9'd40,-10'd161};
ram[13056] = {9'd40,-10'd161};
ram[13057] = {9'd43,-10'd158};
ram[13058] = {9'd46,-10'd154};
ram[13059] = {9'd49,-10'd151};
ram[13060] = {9'd52,-10'd148};
ram[13061] = {9'd55,-10'd145};
ram[13062] = {9'd58,-10'd142};
ram[13063] = {9'd62,-10'd139};
ram[13064] = {9'd65,-10'd136};
ram[13065] = {9'd68,-10'd132};
ram[13066] = {9'd71,-10'd129};
ram[13067] = {9'd74,-10'd126};
ram[13068] = {9'd77,-10'd123};
ram[13069] = {9'd80,-10'd120};
ram[13070] = {9'd84,-10'd117};
ram[13071] = {9'd87,-10'd114};
ram[13072] = {9'd90,-10'd110};
ram[13073] = {9'd93,-10'd107};
ram[13074] = {9'd96,-10'd104};
ram[13075] = {9'd99,-10'd101};
ram[13076] = {-9'd98,-10'd98};
ram[13077] = {-9'd95,-10'd95};
ram[13078] = {-9'd92,-10'd92};
ram[13079] = {-9'd88,-10'd88};
ram[13080] = {-9'd85,-10'd85};
ram[13081] = {-9'd82,-10'd82};
ram[13082] = {-9'd79,-10'd79};
ram[13083] = {-9'd76,-10'd76};
ram[13084] = {-9'd73,-10'd73};
ram[13085] = {-9'd70,-10'd70};
ram[13086] = {-9'd66,-10'd66};
ram[13087] = {-9'd63,-10'd63};
ram[13088] = {-9'd60,-10'd60};
ram[13089] = {-9'd57,-10'd57};
ram[13090] = {-9'd54,-10'd54};
ram[13091] = {-9'd51,-10'd51};
ram[13092] = {-9'd48,-10'd48};
ram[13093] = {-9'd44,-10'd44};
ram[13094] = {-9'd41,-10'd41};
ram[13095] = {-9'd38,-10'd38};
ram[13096] = {-9'd35,-10'd35};
ram[13097] = {-9'd32,-10'd32};
ram[13098] = {-9'd29,-10'd29};
ram[13099] = {-9'd26,-10'd26};
ram[13100] = {-9'd22,-10'd22};
ram[13101] = {-9'd19,-10'd19};
ram[13102] = {-9'd16,-10'd16};
ram[13103] = {-9'd13,-10'd13};
ram[13104] = {-9'd10,-10'd10};
ram[13105] = {-9'd7,-10'd7};
ram[13106] = {-9'd4,-10'd4};
ram[13107] = {9'd0,10'd0};
ram[13108] = {9'd3,10'd3};
ram[13109] = {9'd6,10'd6};
ram[13110] = {9'd9,10'd9};
ram[13111] = {9'd12,10'd12};
ram[13112] = {9'd15,10'd15};
ram[13113] = {9'd18,10'd18};
ram[13114] = {9'd21,10'd21};
ram[13115] = {9'd25,10'd25};
ram[13116] = {9'd28,10'd28};
ram[13117] = {9'd31,10'd31};
ram[13118] = {9'd34,10'd34};
ram[13119] = {9'd37,10'd37};
ram[13120] = {9'd40,10'd40};
ram[13121] = {9'd43,10'd43};
ram[13122] = {9'd47,10'd47};
ram[13123] = {9'd50,10'd50};
ram[13124] = {9'd53,10'd53};
ram[13125] = {9'd56,10'd56};
ram[13126] = {9'd59,10'd59};
ram[13127] = {9'd62,10'd62};
ram[13128] = {9'd65,10'd65};
ram[13129] = {9'd69,10'd69};
ram[13130] = {9'd72,10'd72};
ram[13131] = {9'd75,10'd75};
ram[13132] = {9'd78,10'd78};
ram[13133] = {9'd81,10'd81};
ram[13134] = {9'd84,10'd84};
ram[13135] = {9'd87,10'd87};
ram[13136] = {9'd91,10'd91};
ram[13137] = {9'd94,10'd94};
ram[13138] = {9'd97,10'd97};
ram[13139] = {-9'd100,10'd100};
ram[13140] = {-9'd97,10'd103};
ram[13141] = {-9'd94,10'd106};
ram[13142] = {-9'd91,10'd109};
ram[13143] = {-9'd88,10'd113};
ram[13144] = {-9'd85,10'd116};
ram[13145] = {-9'd81,10'd119};
ram[13146] = {-9'd78,10'd122};
ram[13147] = {-9'd75,10'd125};
ram[13148] = {-9'd72,10'd128};
ram[13149] = {-9'd69,10'd131};
ram[13150] = {-9'd66,10'd135};
ram[13151] = {-9'd63,10'd138};
ram[13152] = {-9'd59,10'd141};
ram[13153] = {-9'd56,10'd144};
ram[13154] = {-9'd53,10'd147};
ram[13155] = {-9'd50,10'd150};
ram[13156] = {-9'd47,10'd153};
ram[13157] = {-9'd44,10'd157};
ram[13158] = {-9'd41,10'd160};
ram[13159] = {-9'd37,10'd163};
ram[13160] = {-9'd34,10'd166};
ram[13161] = {-9'd31,10'd169};
ram[13162] = {-9'd28,10'd172};
ram[13163] = {-9'd25,10'd175};
ram[13164] = {-9'd22,10'd179};
ram[13165] = {-9'd19,10'd182};
ram[13166] = {-9'd15,10'd185};
ram[13167] = {-9'd12,10'd188};
ram[13168] = {-9'd9,10'd191};
ram[13169] = {-9'd6,10'd194};
ram[13170] = {-9'd3,10'd197};
ram[13171] = {9'd0,10'd201};
ram[13172] = {9'd3,10'd204};
ram[13173] = {9'd7,10'd207};
ram[13174] = {9'd10,10'd210};
ram[13175] = {9'd13,10'd213};
ram[13176] = {9'd16,10'd216};
ram[13177] = {9'd19,10'd219};
ram[13178] = {9'd22,10'd223};
ram[13179] = {9'd25,10'd226};
ram[13180] = {9'd29,10'd229};
ram[13181] = {9'd32,10'd232};
ram[13182] = {9'd35,10'd235};
ram[13183] = {9'd38,10'd238};
ram[13184] = {9'd38,10'd238};
ram[13185] = {9'd41,10'd241};
ram[13186] = {9'd44,10'd245};
ram[13187] = {9'd47,10'd248};
ram[13188] = {9'd51,10'd251};
ram[13189] = {9'd54,10'd254};
ram[13190] = {9'd57,10'd257};
ram[13191] = {9'd60,10'd260};
ram[13192] = {9'd63,10'd263};
ram[13193] = {9'd66,10'd267};
ram[13194] = {9'd69,10'd270};
ram[13195] = {9'd73,10'd273};
ram[13196] = {9'd76,10'd276};
ram[13197] = {9'd79,10'd279};
ram[13198] = {9'd82,10'd282};
ram[13199] = {9'd85,10'd285};
ram[13200] = {9'd88,10'd289};
ram[13201] = {9'd91,10'd292};
ram[13202] = {9'd95,10'd295};
ram[13203] = {9'd98,10'd298};
ram[13204] = {-9'd99,10'd301};
ram[13205] = {-9'd96,10'd304};
ram[13206] = {-9'd93,10'd307};
ram[13207] = {-9'd90,10'd311};
ram[13208] = {-9'd87,10'd314};
ram[13209] = {-9'd84,10'd317};
ram[13210] = {-9'd81,10'd320};
ram[13211] = {-9'd77,10'd323};
ram[13212] = {-9'd74,10'd326};
ram[13213] = {-9'd71,10'd329};
ram[13214] = {-9'd68,10'd333};
ram[13215] = {-9'd65,10'd336};
ram[13216] = {-9'd62,10'd339};
ram[13217] = {-9'd59,10'd342};
ram[13218] = {-9'd55,10'd345};
ram[13219] = {-9'd52,10'd348};
ram[13220] = {-9'd49,10'd351};
ram[13221] = {-9'd46,10'd354};
ram[13222] = {-9'd43,10'd358};
ram[13223] = {-9'd40,10'd361};
ram[13224] = {-9'd37,10'd364};
ram[13225] = {-9'd33,10'd367};
ram[13226] = {-9'd30,10'd370};
ram[13227] = {-9'd27,10'd373};
ram[13228] = {-9'd24,10'd376};
ram[13229] = {-9'd21,10'd380};
ram[13230] = {-9'd18,10'd383};
ram[13231] = {-9'd15,10'd386};
ram[13232] = {-9'd11,10'd389};
ram[13233] = {-9'd8,10'd392};
ram[13234] = {-9'd5,10'd395};
ram[13235] = {-9'd2,10'd398};
ram[13236] = {9'd1,-10'd399};
ram[13237] = {9'd4,-10'd396};
ram[13238] = {9'd7,-10'd393};
ram[13239] = {9'd10,-10'd390};
ram[13240] = {9'd14,-10'd387};
ram[13241] = {9'd17,-10'd384};
ram[13242] = {9'd20,-10'd381};
ram[13243] = {9'd23,-10'd377};
ram[13244] = {9'd26,-10'd374};
ram[13245] = {9'd29,-10'd371};
ram[13246] = {9'd32,-10'd368};
ram[13247] = {9'd36,-10'd365};
ram[13248] = {9'd39,-10'd362};
ram[13249] = {9'd42,-10'd359};
ram[13250] = {9'd45,-10'd355};
ram[13251] = {9'd48,-10'd352};
ram[13252] = {9'd51,-10'd349};
ram[13253] = {9'd54,-10'd346};
ram[13254] = {9'd58,-10'd343};
ram[13255] = {9'd61,-10'd340};
ram[13256] = {9'd64,-10'd337};
ram[13257] = {9'd67,-10'd334};
ram[13258] = {9'd70,-10'd330};
ram[13259] = {9'd73,-10'd327};
ram[13260] = {9'd76,-10'd324};
ram[13261] = {9'd80,-10'd321};
ram[13262] = {9'd83,-10'd318};
ram[13263] = {9'd86,-10'd315};
ram[13264] = {9'd89,-10'd312};
ram[13265] = {9'd92,-10'd308};
ram[13266] = {9'd95,-10'd305};
ram[13267] = {9'd98,-10'd302};
ram[13268] = {-9'd99,-10'd299};
ram[13269] = {-9'd96,-10'd296};
ram[13270] = {-9'd92,-10'd293};
ram[13271] = {-9'd89,-10'd290};
ram[13272] = {-9'd86,-10'd286};
ram[13273] = {-9'd83,-10'd283};
ram[13274] = {-9'd80,-10'd280};
ram[13275] = {-9'd77,-10'd277};
ram[13276] = {-9'd74,-10'd274};
ram[13277] = {-9'd70,-10'd271};
ram[13278] = {-9'd67,-10'd268};
ram[13279] = {-9'd64,-10'd264};
ram[13280] = {-9'd61,-10'd261};
ram[13281] = {-9'd58,-10'd258};
ram[13282] = {-9'd55,-10'd255};
ram[13283] = {-9'd52,-10'd252};
ram[13284] = {-9'd48,-10'd249};
ram[13285] = {-9'd45,-10'd246};
ram[13286] = {-9'd42,-10'd242};
ram[13287] = {-9'd39,-10'd239};
ram[13288] = {-9'd36,-10'd236};
ram[13289] = {-9'd33,-10'd233};
ram[13290] = {-9'd30,-10'd230};
ram[13291] = {-9'd26,-10'd227};
ram[13292] = {-9'd23,-10'd224};
ram[13293] = {-9'd20,-10'd220};
ram[13294] = {-9'd17,-10'd217};
ram[13295] = {-9'd14,-10'd214};
ram[13296] = {-9'd11,-10'd211};
ram[13297] = {-9'd8,-10'd208};
ram[13298] = {-9'd4,-10'd205};
ram[13299] = {-9'd1,-10'd202};
ram[13300] = {9'd2,-10'd198};
ram[13301] = {9'd5,-10'd195};
ram[13302] = {9'd8,-10'd192};
ram[13303] = {9'd11,-10'd189};
ram[13304] = {9'd14,-10'd186};
ram[13305] = {9'd18,-10'd183};
ram[13306] = {9'd21,-10'd180};
ram[13307] = {9'd24,-10'd176};
ram[13308] = {9'd27,-10'd173};
ram[13309] = {9'd30,-10'd170};
ram[13310] = {9'd33,-10'd167};
ram[13311] = {9'd36,-10'd164};
ram[13312] = {9'd36,-10'd164};
ram[13313] = {9'd40,-10'd161};
ram[13314] = {9'd43,-10'd158};
ram[13315] = {9'd46,-10'd154};
ram[13316] = {9'd49,-10'd151};
ram[13317] = {9'd52,-10'd148};
ram[13318] = {9'd55,-10'd145};
ram[13319] = {9'd58,-10'd142};
ram[13320] = {9'd62,-10'd139};
ram[13321] = {9'd65,-10'd136};
ram[13322] = {9'd68,-10'd132};
ram[13323] = {9'd71,-10'd129};
ram[13324] = {9'd74,-10'd126};
ram[13325] = {9'd77,-10'd123};
ram[13326] = {9'd80,-10'd120};
ram[13327] = {9'd84,-10'd117};
ram[13328] = {9'd87,-10'd114};
ram[13329] = {9'd90,-10'd110};
ram[13330] = {9'd93,-10'd107};
ram[13331] = {9'd96,-10'd104};
ram[13332] = {9'd99,-10'd101};
ram[13333] = {-9'd98,-10'd98};
ram[13334] = {-9'd95,-10'd95};
ram[13335] = {-9'd92,-10'd92};
ram[13336] = {-9'd88,-10'd88};
ram[13337] = {-9'd85,-10'd85};
ram[13338] = {-9'd82,-10'd82};
ram[13339] = {-9'd79,-10'd79};
ram[13340] = {-9'd76,-10'd76};
ram[13341] = {-9'd73,-10'd73};
ram[13342] = {-9'd70,-10'd70};
ram[13343] = {-9'd66,-10'd66};
ram[13344] = {-9'd63,-10'd63};
ram[13345] = {-9'd60,-10'd60};
ram[13346] = {-9'd57,-10'd57};
ram[13347] = {-9'd54,-10'd54};
ram[13348] = {-9'd51,-10'd51};
ram[13349] = {-9'd48,-10'd48};
ram[13350] = {-9'd44,-10'd44};
ram[13351] = {-9'd41,-10'd41};
ram[13352] = {-9'd38,-10'd38};
ram[13353] = {-9'd35,-10'd35};
ram[13354] = {-9'd32,-10'd32};
ram[13355] = {-9'd29,-10'd29};
ram[13356] = {-9'd26,-10'd26};
ram[13357] = {-9'd22,-10'd22};
ram[13358] = {-9'd19,-10'd19};
ram[13359] = {-9'd16,-10'd16};
ram[13360] = {-9'd13,-10'd13};
ram[13361] = {-9'd10,-10'd10};
ram[13362] = {-9'd7,-10'd7};
ram[13363] = {-9'd4,-10'd4};
ram[13364] = {9'd0,10'd0};
ram[13365] = {9'd3,10'd3};
ram[13366] = {9'd6,10'd6};
ram[13367] = {9'd9,10'd9};
ram[13368] = {9'd12,10'd12};
ram[13369] = {9'd15,10'd15};
ram[13370] = {9'd18,10'd18};
ram[13371] = {9'd21,10'd21};
ram[13372] = {9'd25,10'd25};
ram[13373] = {9'd28,10'd28};
ram[13374] = {9'd31,10'd31};
ram[13375] = {9'd34,10'd34};
ram[13376] = {9'd37,10'd37};
ram[13377] = {9'd40,10'd40};
ram[13378] = {9'd43,10'd43};
ram[13379] = {9'd47,10'd47};
ram[13380] = {9'd50,10'd50};
ram[13381] = {9'd53,10'd53};
ram[13382] = {9'd56,10'd56};
ram[13383] = {9'd59,10'd59};
ram[13384] = {9'd62,10'd62};
ram[13385] = {9'd65,10'd65};
ram[13386] = {9'd69,10'd69};
ram[13387] = {9'd72,10'd72};
ram[13388] = {9'd75,10'd75};
ram[13389] = {9'd78,10'd78};
ram[13390] = {9'd81,10'd81};
ram[13391] = {9'd84,10'd84};
ram[13392] = {9'd87,10'd87};
ram[13393] = {9'd91,10'd91};
ram[13394] = {9'd94,10'd94};
ram[13395] = {9'd97,10'd97};
ram[13396] = {-9'd100,10'd100};
ram[13397] = {-9'd97,10'd103};
ram[13398] = {-9'd94,10'd106};
ram[13399] = {-9'd91,10'd109};
ram[13400] = {-9'd88,10'd113};
ram[13401] = {-9'd85,10'd116};
ram[13402] = {-9'd81,10'd119};
ram[13403] = {-9'd78,10'd122};
ram[13404] = {-9'd75,10'd125};
ram[13405] = {-9'd72,10'd128};
ram[13406] = {-9'd69,10'd131};
ram[13407] = {-9'd66,10'd135};
ram[13408] = {-9'd63,10'd138};
ram[13409] = {-9'd59,10'd141};
ram[13410] = {-9'd56,10'd144};
ram[13411] = {-9'd53,10'd147};
ram[13412] = {-9'd50,10'd150};
ram[13413] = {-9'd47,10'd153};
ram[13414] = {-9'd44,10'd157};
ram[13415] = {-9'd41,10'd160};
ram[13416] = {-9'd37,10'd163};
ram[13417] = {-9'd34,10'd166};
ram[13418] = {-9'd31,10'd169};
ram[13419] = {-9'd28,10'd172};
ram[13420] = {-9'd25,10'd175};
ram[13421] = {-9'd22,10'd179};
ram[13422] = {-9'd19,10'd182};
ram[13423] = {-9'd15,10'd185};
ram[13424] = {-9'd12,10'd188};
ram[13425] = {-9'd9,10'd191};
ram[13426] = {-9'd6,10'd194};
ram[13427] = {-9'd3,10'd197};
ram[13428] = {9'd0,10'd201};
ram[13429] = {9'd3,10'd204};
ram[13430] = {9'd7,10'd207};
ram[13431] = {9'd10,10'd210};
ram[13432] = {9'd13,10'd213};
ram[13433] = {9'd16,10'd216};
ram[13434] = {9'd19,10'd219};
ram[13435] = {9'd22,10'd223};
ram[13436] = {9'd25,10'd226};
ram[13437] = {9'd29,10'd229};
ram[13438] = {9'd32,10'd232};
ram[13439] = {9'd35,10'd235};
ram[13440] = {9'd35,10'd235};
ram[13441] = {9'd38,10'd238};
ram[13442] = {9'd41,10'd241};
ram[13443] = {9'd44,10'd245};
ram[13444] = {9'd47,10'd248};
ram[13445] = {9'd51,10'd251};
ram[13446] = {9'd54,10'd254};
ram[13447] = {9'd57,10'd257};
ram[13448] = {9'd60,10'd260};
ram[13449] = {9'd63,10'd263};
ram[13450] = {9'd66,10'd267};
ram[13451] = {9'd69,10'd270};
ram[13452] = {9'd73,10'd273};
ram[13453] = {9'd76,10'd276};
ram[13454] = {9'd79,10'd279};
ram[13455] = {9'd82,10'd282};
ram[13456] = {9'd85,10'd285};
ram[13457] = {9'd88,10'd289};
ram[13458] = {9'd91,10'd292};
ram[13459] = {9'd95,10'd295};
ram[13460] = {9'd98,10'd298};
ram[13461] = {-9'd99,10'd301};
ram[13462] = {-9'd96,10'd304};
ram[13463] = {-9'd93,10'd307};
ram[13464] = {-9'd90,10'd311};
ram[13465] = {-9'd87,10'd314};
ram[13466] = {-9'd84,10'd317};
ram[13467] = {-9'd81,10'd320};
ram[13468] = {-9'd77,10'd323};
ram[13469] = {-9'd74,10'd326};
ram[13470] = {-9'd71,10'd329};
ram[13471] = {-9'd68,10'd333};
ram[13472] = {-9'd65,10'd336};
ram[13473] = {-9'd62,10'd339};
ram[13474] = {-9'd59,10'd342};
ram[13475] = {-9'd55,10'd345};
ram[13476] = {-9'd52,10'd348};
ram[13477] = {-9'd49,10'd351};
ram[13478] = {-9'd46,10'd354};
ram[13479] = {-9'd43,10'd358};
ram[13480] = {-9'd40,10'd361};
ram[13481] = {-9'd37,10'd364};
ram[13482] = {-9'd33,10'd367};
ram[13483] = {-9'd30,10'd370};
ram[13484] = {-9'd27,10'd373};
ram[13485] = {-9'd24,10'd376};
ram[13486] = {-9'd21,10'd380};
ram[13487] = {-9'd18,10'd383};
ram[13488] = {-9'd15,10'd386};
ram[13489] = {-9'd11,10'd389};
ram[13490] = {-9'd8,10'd392};
ram[13491] = {-9'd5,10'd395};
ram[13492] = {-9'd2,10'd398};
ram[13493] = {9'd1,-10'd399};
ram[13494] = {9'd4,-10'd396};
ram[13495] = {9'd7,-10'd393};
ram[13496] = {9'd10,-10'd390};
ram[13497] = {9'd14,-10'd387};
ram[13498] = {9'd17,-10'd384};
ram[13499] = {9'd20,-10'd381};
ram[13500] = {9'd23,-10'd377};
ram[13501] = {9'd26,-10'd374};
ram[13502] = {9'd29,-10'd371};
ram[13503] = {9'd32,-10'd368};
ram[13504] = {9'd36,-10'd365};
ram[13505] = {9'd39,-10'd362};
ram[13506] = {9'd42,-10'd359};
ram[13507] = {9'd45,-10'd355};
ram[13508] = {9'd48,-10'd352};
ram[13509] = {9'd51,-10'd349};
ram[13510] = {9'd54,-10'd346};
ram[13511] = {9'd58,-10'd343};
ram[13512] = {9'd61,-10'd340};
ram[13513] = {9'd64,-10'd337};
ram[13514] = {9'd67,-10'd334};
ram[13515] = {9'd70,-10'd330};
ram[13516] = {9'd73,-10'd327};
ram[13517] = {9'd76,-10'd324};
ram[13518] = {9'd80,-10'd321};
ram[13519] = {9'd83,-10'd318};
ram[13520] = {9'd86,-10'd315};
ram[13521] = {9'd89,-10'd312};
ram[13522] = {9'd92,-10'd308};
ram[13523] = {9'd95,-10'd305};
ram[13524] = {9'd98,-10'd302};
ram[13525] = {-9'd99,-10'd299};
ram[13526] = {-9'd96,-10'd296};
ram[13527] = {-9'd92,-10'd293};
ram[13528] = {-9'd89,-10'd290};
ram[13529] = {-9'd86,-10'd286};
ram[13530] = {-9'd83,-10'd283};
ram[13531] = {-9'd80,-10'd280};
ram[13532] = {-9'd77,-10'd277};
ram[13533] = {-9'd74,-10'd274};
ram[13534] = {-9'd70,-10'd271};
ram[13535] = {-9'd67,-10'd268};
ram[13536] = {-9'd64,-10'd264};
ram[13537] = {-9'd61,-10'd261};
ram[13538] = {-9'd58,-10'd258};
ram[13539] = {-9'd55,-10'd255};
ram[13540] = {-9'd52,-10'd252};
ram[13541] = {-9'd48,-10'd249};
ram[13542] = {-9'd45,-10'd246};
ram[13543] = {-9'd42,-10'd242};
ram[13544] = {-9'd39,-10'd239};
ram[13545] = {-9'd36,-10'd236};
ram[13546] = {-9'd33,-10'd233};
ram[13547] = {-9'd30,-10'd230};
ram[13548] = {-9'd26,-10'd227};
ram[13549] = {-9'd23,-10'd224};
ram[13550] = {-9'd20,-10'd220};
ram[13551] = {-9'd17,-10'd217};
ram[13552] = {-9'd14,-10'd214};
ram[13553] = {-9'd11,-10'd211};
ram[13554] = {-9'd8,-10'd208};
ram[13555] = {-9'd4,-10'd205};
ram[13556] = {-9'd1,-10'd202};
ram[13557] = {9'd2,-10'd198};
ram[13558] = {9'd5,-10'd195};
ram[13559] = {9'd8,-10'd192};
ram[13560] = {9'd11,-10'd189};
ram[13561] = {9'd14,-10'd186};
ram[13562] = {9'd18,-10'd183};
ram[13563] = {9'd21,-10'd180};
ram[13564] = {9'd24,-10'd176};
ram[13565] = {9'd27,-10'd173};
ram[13566] = {9'd30,-10'd170};
ram[13567] = {9'd33,-10'd167};
ram[13568] = {9'd33,-10'd167};
ram[13569] = {9'd36,-10'd164};
ram[13570] = {9'd40,-10'd161};
ram[13571] = {9'd43,-10'd158};
ram[13572] = {9'd46,-10'd154};
ram[13573] = {9'd49,-10'd151};
ram[13574] = {9'd52,-10'd148};
ram[13575] = {9'd55,-10'd145};
ram[13576] = {9'd58,-10'd142};
ram[13577] = {9'd62,-10'd139};
ram[13578] = {9'd65,-10'd136};
ram[13579] = {9'd68,-10'd132};
ram[13580] = {9'd71,-10'd129};
ram[13581] = {9'd74,-10'd126};
ram[13582] = {9'd77,-10'd123};
ram[13583] = {9'd80,-10'd120};
ram[13584] = {9'd84,-10'd117};
ram[13585] = {9'd87,-10'd114};
ram[13586] = {9'd90,-10'd110};
ram[13587] = {9'd93,-10'd107};
ram[13588] = {9'd96,-10'd104};
ram[13589] = {9'd99,-10'd101};
ram[13590] = {-9'd98,-10'd98};
ram[13591] = {-9'd95,-10'd95};
ram[13592] = {-9'd92,-10'd92};
ram[13593] = {-9'd88,-10'd88};
ram[13594] = {-9'd85,-10'd85};
ram[13595] = {-9'd82,-10'd82};
ram[13596] = {-9'd79,-10'd79};
ram[13597] = {-9'd76,-10'd76};
ram[13598] = {-9'd73,-10'd73};
ram[13599] = {-9'd70,-10'd70};
ram[13600] = {-9'd66,-10'd66};
ram[13601] = {-9'd63,-10'd63};
ram[13602] = {-9'd60,-10'd60};
ram[13603] = {-9'd57,-10'd57};
ram[13604] = {-9'd54,-10'd54};
ram[13605] = {-9'd51,-10'd51};
ram[13606] = {-9'd48,-10'd48};
ram[13607] = {-9'd44,-10'd44};
ram[13608] = {-9'd41,-10'd41};
ram[13609] = {-9'd38,-10'd38};
ram[13610] = {-9'd35,-10'd35};
ram[13611] = {-9'd32,-10'd32};
ram[13612] = {-9'd29,-10'd29};
ram[13613] = {-9'd26,-10'd26};
ram[13614] = {-9'd22,-10'd22};
ram[13615] = {-9'd19,-10'd19};
ram[13616] = {-9'd16,-10'd16};
ram[13617] = {-9'd13,-10'd13};
ram[13618] = {-9'd10,-10'd10};
ram[13619] = {-9'd7,-10'd7};
ram[13620] = {-9'd4,-10'd4};
ram[13621] = {9'd0,10'd0};
ram[13622] = {9'd3,10'd3};
ram[13623] = {9'd6,10'd6};
ram[13624] = {9'd9,10'd9};
ram[13625] = {9'd12,10'd12};
ram[13626] = {9'd15,10'd15};
ram[13627] = {9'd18,10'd18};
ram[13628] = {9'd21,10'd21};
ram[13629] = {9'd25,10'd25};
ram[13630] = {9'd28,10'd28};
ram[13631] = {9'd31,10'd31};
ram[13632] = {9'd34,10'd34};
ram[13633] = {9'd37,10'd37};
ram[13634] = {9'd40,10'd40};
ram[13635] = {9'd43,10'd43};
ram[13636] = {9'd47,10'd47};
ram[13637] = {9'd50,10'd50};
ram[13638] = {9'd53,10'd53};
ram[13639] = {9'd56,10'd56};
ram[13640] = {9'd59,10'd59};
ram[13641] = {9'd62,10'd62};
ram[13642] = {9'd65,10'd65};
ram[13643] = {9'd69,10'd69};
ram[13644] = {9'd72,10'd72};
ram[13645] = {9'd75,10'd75};
ram[13646] = {9'd78,10'd78};
ram[13647] = {9'd81,10'd81};
ram[13648] = {9'd84,10'd84};
ram[13649] = {9'd87,10'd87};
ram[13650] = {9'd91,10'd91};
ram[13651] = {9'd94,10'd94};
ram[13652] = {9'd97,10'd97};
ram[13653] = {-9'd100,10'd100};
ram[13654] = {-9'd97,10'd103};
ram[13655] = {-9'd94,10'd106};
ram[13656] = {-9'd91,10'd109};
ram[13657] = {-9'd88,10'd113};
ram[13658] = {-9'd85,10'd116};
ram[13659] = {-9'd81,10'd119};
ram[13660] = {-9'd78,10'd122};
ram[13661] = {-9'd75,10'd125};
ram[13662] = {-9'd72,10'd128};
ram[13663] = {-9'd69,10'd131};
ram[13664] = {-9'd66,10'd135};
ram[13665] = {-9'd63,10'd138};
ram[13666] = {-9'd59,10'd141};
ram[13667] = {-9'd56,10'd144};
ram[13668] = {-9'd53,10'd147};
ram[13669] = {-9'd50,10'd150};
ram[13670] = {-9'd47,10'd153};
ram[13671] = {-9'd44,10'd157};
ram[13672] = {-9'd41,10'd160};
ram[13673] = {-9'd37,10'd163};
ram[13674] = {-9'd34,10'd166};
ram[13675] = {-9'd31,10'd169};
ram[13676] = {-9'd28,10'd172};
ram[13677] = {-9'd25,10'd175};
ram[13678] = {-9'd22,10'd179};
ram[13679] = {-9'd19,10'd182};
ram[13680] = {-9'd15,10'd185};
ram[13681] = {-9'd12,10'd188};
ram[13682] = {-9'd9,10'd191};
ram[13683] = {-9'd6,10'd194};
ram[13684] = {-9'd3,10'd197};
ram[13685] = {9'd0,10'd201};
ram[13686] = {9'd3,10'd204};
ram[13687] = {9'd7,10'd207};
ram[13688] = {9'd10,10'd210};
ram[13689] = {9'd13,10'd213};
ram[13690] = {9'd16,10'd216};
ram[13691] = {9'd19,10'd219};
ram[13692] = {9'd22,10'd223};
ram[13693] = {9'd25,10'd226};
ram[13694] = {9'd29,10'd229};
ram[13695] = {9'd32,10'd232};
ram[13696] = {9'd32,10'd232};
ram[13697] = {9'd35,10'd235};
ram[13698] = {9'd38,10'd238};
ram[13699] = {9'd41,10'd241};
ram[13700] = {9'd44,10'd245};
ram[13701] = {9'd47,10'd248};
ram[13702] = {9'd51,10'd251};
ram[13703] = {9'd54,10'd254};
ram[13704] = {9'd57,10'd257};
ram[13705] = {9'd60,10'd260};
ram[13706] = {9'd63,10'd263};
ram[13707] = {9'd66,10'd267};
ram[13708] = {9'd69,10'd270};
ram[13709] = {9'd73,10'd273};
ram[13710] = {9'd76,10'd276};
ram[13711] = {9'd79,10'd279};
ram[13712] = {9'd82,10'd282};
ram[13713] = {9'd85,10'd285};
ram[13714] = {9'd88,10'd289};
ram[13715] = {9'd91,10'd292};
ram[13716] = {9'd95,10'd295};
ram[13717] = {9'd98,10'd298};
ram[13718] = {-9'd99,10'd301};
ram[13719] = {-9'd96,10'd304};
ram[13720] = {-9'd93,10'd307};
ram[13721] = {-9'd90,10'd311};
ram[13722] = {-9'd87,10'd314};
ram[13723] = {-9'd84,10'd317};
ram[13724] = {-9'd81,10'd320};
ram[13725] = {-9'd77,10'd323};
ram[13726] = {-9'd74,10'd326};
ram[13727] = {-9'd71,10'd329};
ram[13728] = {-9'd68,10'd333};
ram[13729] = {-9'd65,10'd336};
ram[13730] = {-9'd62,10'd339};
ram[13731] = {-9'd59,10'd342};
ram[13732] = {-9'd55,10'd345};
ram[13733] = {-9'd52,10'd348};
ram[13734] = {-9'd49,10'd351};
ram[13735] = {-9'd46,10'd354};
ram[13736] = {-9'd43,10'd358};
ram[13737] = {-9'd40,10'd361};
ram[13738] = {-9'd37,10'd364};
ram[13739] = {-9'd33,10'd367};
ram[13740] = {-9'd30,10'd370};
ram[13741] = {-9'd27,10'd373};
ram[13742] = {-9'd24,10'd376};
ram[13743] = {-9'd21,10'd380};
ram[13744] = {-9'd18,10'd383};
ram[13745] = {-9'd15,10'd386};
ram[13746] = {-9'd11,10'd389};
ram[13747] = {-9'd8,10'd392};
ram[13748] = {-9'd5,10'd395};
ram[13749] = {-9'd2,10'd398};
ram[13750] = {9'd1,-10'd399};
ram[13751] = {9'd4,-10'd396};
ram[13752] = {9'd7,-10'd393};
ram[13753] = {9'd10,-10'd390};
ram[13754] = {9'd14,-10'd387};
ram[13755] = {9'd17,-10'd384};
ram[13756] = {9'd20,-10'd381};
ram[13757] = {9'd23,-10'd377};
ram[13758] = {9'd26,-10'd374};
ram[13759] = {9'd29,-10'd371};
ram[13760] = {9'd32,-10'd368};
ram[13761] = {9'd36,-10'd365};
ram[13762] = {9'd39,-10'd362};
ram[13763] = {9'd42,-10'd359};
ram[13764] = {9'd45,-10'd355};
ram[13765] = {9'd48,-10'd352};
ram[13766] = {9'd51,-10'd349};
ram[13767] = {9'd54,-10'd346};
ram[13768] = {9'd58,-10'd343};
ram[13769] = {9'd61,-10'd340};
ram[13770] = {9'd64,-10'd337};
ram[13771] = {9'd67,-10'd334};
ram[13772] = {9'd70,-10'd330};
ram[13773] = {9'd73,-10'd327};
ram[13774] = {9'd76,-10'd324};
ram[13775] = {9'd80,-10'd321};
ram[13776] = {9'd83,-10'd318};
ram[13777] = {9'd86,-10'd315};
ram[13778] = {9'd89,-10'd312};
ram[13779] = {9'd92,-10'd308};
ram[13780] = {9'd95,-10'd305};
ram[13781] = {9'd98,-10'd302};
ram[13782] = {-9'd99,-10'd299};
ram[13783] = {-9'd96,-10'd296};
ram[13784] = {-9'd92,-10'd293};
ram[13785] = {-9'd89,-10'd290};
ram[13786] = {-9'd86,-10'd286};
ram[13787] = {-9'd83,-10'd283};
ram[13788] = {-9'd80,-10'd280};
ram[13789] = {-9'd77,-10'd277};
ram[13790] = {-9'd74,-10'd274};
ram[13791] = {-9'd70,-10'd271};
ram[13792] = {-9'd67,-10'd268};
ram[13793] = {-9'd64,-10'd264};
ram[13794] = {-9'd61,-10'd261};
ram[13795] = {-9'd58,-10'd258};
ram[13796] = {-9'd55,-10'd255};
ram[13797] = {-9'd52,-10'd252};
ram[13798] = {-9'd48,-10'd249};
ram[13799] = {-9'd45,-10'd246};
ram[13800] = {-9'd42,-10'd242};
ram[13801] = {-9'd39,-10'd239};
ram[13802] = {-9'd36,-10'd236};
ram[13803] = {-9'd33,-10'd233};
ram[13804] = {-9'd30,-10'd230};
ram[13805] = {-9'd26,-10'd227};
ram[13806] = {-9'd23,-10'd224};
ram[13807] = {-9'd20,-10'd220};
ram[13808] = {-9'd17,-10'd217};
ram[13809] = {-9'd14,-10'd214};
ram[13810] = {-9'd11,-10'd211};
ram[13811] = {-9'd8,-10'd208};
ram[13812] = {-9'd4,-10'd205};
ram[13813] = {-9'd1,-10'd202};
ram[13814] = {9'd2,-10'd198};
ram[13815] = {9'd5,-10'd195};
ram[13816] = {9'd8,-10'd192};
ram[13817] = {9'd11,-10'd189};
ram[13818] = {9'd14,-10'd186};
ram[13819] = {9'd18,-10'd183};
ram[13820] = {9'd21,-10'd180};
ram[13821] = {9'd24,-10'd176};
ram[13822] = {9'd27,-10'd173};
ram[13823] = {9'd30,-10'd170};
ram[13824] = {9'd30,-10'd170};
ram[13825] = {9'd33,-10'd167};
ram[13826] = {9'd36,-10'd164};
ram[13827] = {9'd40,-10'd161};
ram[13828] = {9'd43,-10'd158};
ram[13829] = {9'd46,-10'd154};
ram[13830] = {9'd49,-10'd151};
ram[13831] = {9'd52,-10'd148};
ram[13832] = {9'd55,-10'd145};
ram[13833] = {9'd58,-10'd142};
ram[13834] = {9'd62,-10'd139};
ram[13835] = {9'd65,-10'd136};
ram[13836] = {9'd68,-10'd132};
ram[13837] = {9'd71,-10'd129};
ram[13838] = {9'd74,-10'd126};
ram[13839] = {9'd77,-10'd123};
ram[13840] = {9'd80,-10'd120};
ram[13841] = {9'd84,-10'd117};
ram[13842] = {9'd87,-10'd114};
ram[13843] = {9'd90,-10'd110};
ram[13844] = {9'd93,-10'd107};
ram[13845] = {9'd96,-10'd104};
ram[13846] = {9'd99,-10'd101};
ram[13847] = {-9'd98,-10'd98};
ram[13848] = {-9'd95,-10'd95};
ram[13849] = {-9'd92,-10'd92};
ram[13850] = {-9'd88,-10'd88};
ram[13851] = {-9'd85,-10'd85};
ram[13852] = {-9'd82,-10'd82};
ram[13853] = {-9'd79,-10'd79};
ram[13854] = {-9'd76,-10'd76};
ram[13855] = {-9'd73,-10'd73};
ram[13856] = {-9'd70,-10'd70};
ram[13857] = {-9'd66,-10'd66};
ram[13858] = {-9'd63,-10'd63};
ram[13859] = {-9'd60,-10'd60};
ram[13860] = {-9'd57,-10'd57};
ram[13861] = {-9'd54,-10'd54};
ram[13862] = {-9'd51,-10'd51};
ram[13863] = {-9'd48,-10'd48};
ram[13864] = {-9'd44,-10'd44};
ram[13865] = {-9'd41,-10'd41};
ram[13866] = {-9'd38,-10'd38};
ram[13867] = {-9'd35,-10'd35};
ram[13868] = {-9'd32,-10'd32};
ram[13869] = {-9'd29,-10'd29};
ram[13870] = {-9'd26,-10'd26};
ram[13871] = {-9'd22,-10'd22};
ram[13872] = {-9'd19,-10'd19};
ram[13873] = {-9'd16,-10'd16};
ram[13874] = {-9'd13,-10'd13};
ram[13875] = {-9'd10,-10'd10};
ram[13876] = {-9'd7,-10'd7};
ram[13877] = {-9'd4,-10'd4};
ram[13878] = {9'd0,10'd0};
ram[13879] = {9'd3,10'd3};
ram[13880] = {9'd6,10'd6};
ram[13881] = {9'd9,10'd9};
ram[13882] = {9'd12,10'd12};
ram[13883] = {9'd15,10'd15};
ram[13884] = {9'd18,10'd18};
ram[13885] = {9'd21,10'd21};
ram[13886] = {9'd25,10'd25};
ram[13887] = {9'd28,10'd28};
ram[13888] = {9'd31,10'd31};
ram[13889] = {9'd34,10'd34};
ram[13890] = {9'd37,10'd37};
ram[13891] = {9'd40,10'd40};
ram[13892] = {9'd43,10'd43};
ram[13893] = {9'd47,10'd47};
ram[13894] = {9'd50,10'd50};
ram[13895] = {9'd53,10'd53};
ram[13896] = {9'd56,10'd56};
ram[13897] = {9'd59,10'd59};
ram[13898] = {9'd62,10'd62};
ram[13899] = {9'd65,10'd65};
ram[13900] = {9'd69,10'd69};
ram[13901] = {9'd72,10'd72};
ram[13902] = {9'd75,10'd75};
ram[13903] = {9'd78,10'd78};
ram[13904] = {9'd81,10'd81};
ram[13905] = {9'd84,10'd84};
ram[13906] = {9'd87,10'd87};
ram[13907] = {9'd91,10'd91};
ram[13908] = {9'd94,10'd94};
ram[13909] = {9'd97,10'd97};
ram[13910] = {-9'd100,10'd100};
ram[13911] = {-9'd97,10'd103};
ram[13912] = {-9'd94,10'd106};
ram[13913] = {-9'd91,10'd109};
ram[13914] = {-9'd88,10'd113};
ram[13915] = {-9'd85,10'd116};
ram[13916] = {-9'd81,10'd119};
ram[13917] = {-9'd78,10'd122};
ram[13918] = {-9'd75,10'd125};
ram[13919] = {-9'd72,10'd128};
ram[13920] = {-9'd69,10'd131};
ram[13921] = {-9'd66,10'd135};
ram[13922] = {-9'd63,10'd138};
ram[13923] = {-9'd59,10'd141};
ram[13924] = {-9'd56,10'd144};
ram[13925] = {-9'd53,10'd147};
ram[13926] = {-9'd50,10'd150};
ram[13927] = {-9'd47,10'd153};
ram[13928] = {-9'd44,10'd157};
ram[13929] = {-9'd41,10'd160};
ram[13930] = {-9'd37,10'd163};
ram[13931] = {-9'd34,10'd166};
ram[13932] = {-9'd31,10'd169};
ram[13933] = {-9'd28,10'd172};
ram[13934] = {-9'd25,10'd175};
ram[13935] = {-9'd22,10'd179};
ram[13936] = {-9'd19,10'd182};
ram[13937] = {-9'd15,10'd185};
ram[13938] = {-9'd12,10'd188};
ram[13939] = {-9'd9,10'd191};
ram[13940] = {-9'd6,10'd194};
ram[13941] = {-9'd3,10'd197};
ram[13942] = {9'd0,10'd201};
ram[13943] = {9'd3,10'd204};
ram[13944] = {9'd7,10'd207};
ram[13945] = {9'd10,10'd210};
ram[13946] = {9'd13,10'd213};
ram[13947] = {9'd16,10'd216};
ram[13948] = {9'd19,10'd219};
ram[13949] = {9'd22,10'd223};
ram[13950] = {9'd25,10'd226};
ram[13951] = {9'd29,10'd229};
ram[13952] = {9'd29,10'd229};
ram[13953] = {9'd32,10'd232};
ram[13954] = {9'd35,10'd235};
ram[13955] = {9'd38,10'd238};
ram[13956] = {9'd41,10'd241};
ram[13957] = {9'd44,10'd245};
ram[13958] = {9'd47,10'd248};
ram[13959] = {9'd51,10'd251};
ram[13960] = {9'd54,10'd254};
ram[13961] = {9'd57,10'd257};
ram[13962] = {9'd60,10'd260};
ram[13963] = {9'd63,10'd263};
ram[13964] = {9'd66,10'd267};
ram[13965] = {9'd69,10'd270};
ram[13966] = {9'd73,10'd273};
ram[13967] = {9'd76,10'd276};
ram[13968] = {9'd79,10'd279};
ram[13969] = {9'd82,10'd282};
ram[13970] = {9'd85,10'd285};
ram[13971] = {9'd88,10'd289};
ram[13972] = {9'd91,10'd292};
ram[13973] = {9'd95,10'd295};
ram[13974] = {9'd98,10'd298};
ram[13975] = {-9'd99,10'd301};
ram[13976] = {-9'd96,10'd304};
ram[13977] = {-9'd93,10'd307};
ram[13978] = {-9'd90,10'd311};
ram[13979] = {-9'd87,10'd314};
ram[13980] = {-9'd84,10'd317};
ram[13981] = {-9'd81,10'd320};
ram[13982] = {-9'd77,10'd323};
ram[13983] = {-9'd74,10'd326};
ram[13984] = {-9'd71,10'd329};
ram[13985] = {-9'd68,10'd333};
ram[13986] = {-9'd65,10'd336};
ram[13987] = {-9'd62,10'd339};
ram[13988] = {-9'd59,10'd342};
ram[13989] = {-9'd55,10'd345};
ram[13990] = {-9'd52,10'd348};
ram[13991] = {-9'd49,10'd351};
ram[13992] = {-9'd46,10'd354};
ram[13993] = {-9'd43,10'd358};
ram[13994] = {-9'd40,10'd361};
ram[13995] = {-9'd37,10'd364};
ram[13996] = {-9'd33,10'd367};
ram[13997] = {-9'd30,10'd370};
ram[13998] = {-9'd27,10'd373};
ram[13999] = {-9'd24,10'd376};
ram[14000] = {-9'd21,10'd380};
ram[14001] = {-9'd18,10'd383};
ram[14002] = {-9'd15,10'd386};
ram[14003] = {-9'd11,10'd389};
ram[14004] = {-9'd8,10'd392};
ram[14005] = {-9'd5,10'd395};
ram[14006] = {-9'd2,10'd398};
ram[14007] = {9'd1,-10'd399};
ram[14008] = {9'd4,-10'd396};
ram[14009] = {9'd7,-10'd393};
ram[14010] = {9'd10,-10'd390};
ram[14011] = {9'd14,-10'd387};
ram[14012] = {9'd17,-10'd384};
ram[14013] = {9'd20,-10'd381};
ram[14014] = {9'd23,-10'd377};
ram[14015] = {9'd26,-10'd374};
ram[14016] = {9'd29,-10'd371};
ram[14017] = {9'd32,-10'd368};
ram[14018] = {9'd36,-10'd365};
ram[14019] = {9'd39,-10'd362};
ram[14020] = {9'd42,-10'd359};
ram[14021] = {9'd45,-10'd355};
ram[14022] = {9'd48,-10'd352};
ram[14023] = {9'd51,-10'd349};
ram[14024] = {9'd54,-10'd346};
ram[14025] = {9'd58,-10'd343};
ram[14026] = {9'd61,-10'd340};
ram[14027] = {9'd64,-10'd337};
ram[14028] = {9'd67,-10'd334};
ram[14029] = {9'd70,-10'd330};
ram[14030] = {9'd73,-10'd327};
ram[14031] = {9'd76,-10'd324};
ram[14032] = {9'd80,-10'd321};
ram[14033] = {9'd83,-10'd318};
ram[14034] = {9'd86,-10'd315};
ram[14035] = {9'd89,-10'd312};
ram[14036] = {9'd92,-10'd308};
ram[14037] = {9'd95,-10'd305};
ram[14038] = {9'd98,-10'd302};
ram[14039] = {-9'd99,-10'd299};
ram[14040] = {-9'd96,-10'd296};
ram[14041] = {-9'd92,-10'd293};
ram[14042] = {-9'd89,-10'd290};
ram[14043] = {-9'd86,-10'd286};
ram[14044] = {-9'd83,-10'd283};
ram[14045] = {-9'd80,-10'd280};
ram[14046] = {-9'd77,-10'd277};
ram[14047] = {-9'd74,-10'd274};
ram[14048] = {-9'd70,-10'd271};
ram[14049] = {-9'd67,-10'd268};
ram[14050] = {-9'd64,-10'd264};
ram[14051] = {-9'd61,-10'd261};
ram[14052] = {-9'd58,-10'd258};
ram[14053] = {-9'd55,-10'd255};
ram[14054] = {-9'd52,-10'd252};
ram[14055] = {-9'd48,-10'd249};
ram[14056] = {-9'd45,-10'd246};
ram[14057] = {-9'd42,-10'd242};
ram[14058] = {-9'd39,-10'd239};
ram[14059] = {-9'd36,-10'd236};
ram[14060] = {-9'd33,-10'd233};
ram[14061] = {-9'd30,-10'd230};
ram[14062] = {-9'd26,-10'd227};
ram[14063] = {-9'd23,-10'd224};
ram[14064] = {-9'd20,-10'd220};
ram[14065] = {-9'd17,-10'd217};
ram[14066] = {-9'd14,-10'd214};
ram[14067] = {-9'd11,-10'd211};
ram[14068] = {-9'd8,-10'd208};
ram[14069] = {-9'd4,-10'd205};
ram[14070] = {-9'd1,-10'd202};
ram[14071] = {9'd2,-10'd198};
ram[14072] = {9'd5,-10'd195};
ram[14073] = {9'd8,-10'd192};
ram[14074] = {9'd11,-10'd189};
ram[14075] = {9'd14,-10'd186};
ram[14076] = {9'd18,-10'd183};
ram[14077] = {9'd21,-10'd180};
ram[14078] = {9'd24,-10'd176};
ram[14079] = {9'd27,-10'd173};
ram[14080] = {9'd27,-10'd173};
ram[14081] = {9'd30,-10'd170};
ram[14082] = {9'd33,-10'd167};
ram[14083] = {9'd36,-10'd164};
ram[14084] = {9'd40,-10'd161};
ram[14085] = {9'd43,-10'd158};
ram[14086] = {9'd46,-10'd154};
ram[14087] = {9'd49,-10'd151};
ram[14088] = {9'd52,-10'd148};
ram[14089] = {9'd55,-10'd145};
ram[14090] = {9'd58,-10'd142};
ram[14091] = {9'd62,-10'd139};
ram[14092] = {9'd65,-10'd136};
ram[14093] = {9'd68,-10'd132};
ram[14094] = {9'd71,-10'd129};
ram[14095] = {9'd74,-10'd126};
ram[14096] = {9'd77,-10'd123};
ram[14097] = {9'd80,-10'd120};
ram[14098] = {9'd84,-10'd117};
ram[14099] = {9'd87,-10'd114};
ram[14100] = {9'd90,-10'd110};
ram[14101] = {9'd93,-10'd107};
ram[14102] = {9'd96,-10'd104};
ram[14103] = {9'd99,-10'd101};
ram[14104] = {-9'd98,-10'd98};
ram[14105] = {-9'd95,-10'd95};
ram[14106] = {-9'd92,-10'd92};
ram[14107] = {-9'd88,-10'd88};
ram[14108] = {-9'd85,-10'd85};
ram[14109] = {-9'd82,-10'd82};
ram[14110] = {-9'd79,-10'd79};
ram[14111] = {-9'd76,-10'd76};
ram[14112] = {-9'd73,-10'd73};
ram[14113] = {-9'd70,-10'd70};
ram[14114] = {-9'd66,-10'd66};
ram[14115] = {-9'd63,-10'd63};
ram[14116] = {-9'd60,-10'd60};
ram[14117] = {-9'd57,-10'd57};
ram[14118] = {-9'd54,-10'd54};
ram[14119] = {-9'd51,-10'd51};
ram[14120] = {-9'd48,-10'd48};
ram[14121] = {-9'd44,-10'd44};
ram[14122] = {-9'd41,-10'd41};
ram[14123] = {-9'd38,-10'd38};
ram[14124] = {-9'd35,-10'd35};
ram[14125] = {-9'd32,-10'd32};
ram[14126] = {-9'd29,-10'd29};
ram[14127] = {-9'd26,-10'd26};
ram[14128] = {-9'd22,-10'd22};
ram[14129] = {-9'd19,-10'd19};
ram[14130] = {-9'd16,-10'd16};
ram[14131] = {-9'd13,-10'd13};
ram[14132] = {-9'd10,-10'd10};
ram[14133] = {-9'd7,-10'd7};
ram[14134] = {-9'd4,-10'd4};
ram[14135] = {9'd0,10'd0};
ram[14136] = {9'd3,10'd3};
ram[14137] = {9'd6,10'd6};
ram[14138] = {9'd9,10'd9};
ram[14139] = {9'd12,10'd12};
ram[14140] = {9'd15,10'd15};
ram[14141] = {9'd18,10'd18};
ram[14142] = {9'd21,10'd21};
ram[14143] = {9'd25,10'd25};
ram[14144] = {9'd28,10'd28};
ram[14145] = {9'd31,10'd31};
ram[14146] = {9'd34,10'd34};
ram[14147] = {9'd37,10'd37};
ram[14148] = {9'd40,10'd40};
ram[14149] = {9'd43,10'd43};
ram[14150] = {9'd47,10'd47};
ram[14151] = {9'd50,10'd50};
ram[14152] = {9'd53,10'd53};
ram[14153] = {9'd56,10'd56};
ram[14154] = {9'd59,10'd59};
ram[14155] = {9'd62,10'd62};
ram[14156] = {9'd65,10'd65};
ram[14157] = {9'd69,10'd69};
ram[14158] = {9'd72,10'd72};
ram[14159] = {9'd75,10'd75};
ram[14160] = {9'd78,10'd78};
ram[14161] = {9'd81,10'd81};
ram[14162] = {9'd84,10'd84};
ram[14163] = {9'd87,10'd87};
ram[14164] = {9'd91,10'd91};
ram[14165] = {9'd94,10'd94};
ram[14166] = {9'd97,10'd97};
ram[14167] = {-9'd100,10'd100};
ram[14168] = {-9'd97,10'd103};
ram[14169] = {-9'd94,10'd106};
ram[14170] = {-9'd91,10'd109};
ram[14171] = {-9'd88,10'd113};
ram[14172] = {-9'd85,10'd116};
ram[14173] = {-9'd81,10'd119};
ram[14174] = {-9'd78,10'd122};
ram[14175] = {-9'd75,10'd125};
ram[14176] = {-9'd72,10'd128};
ram[14177] = {-9'd69,10'd131};
ram[14178] = {-9'd66,10'd135};
ram[14179] = {-9'd63,10'd138};
ram[14180] = {-9'd59,10'd141};
ram[14181] = {-9'd56,10'd144};
ram[14182] = {-9'd53,10'd147};
ram[14183] = {-9'd50,10'd150};
ram[14184] = {-9'd47,10'd153};
ram[14185] = {-9'd44,10'd157};
ram[14186] = {-9'd41,10'd160};
ram[14187] = {-9'd37,10'd163};
ram[14188] = {-9'd34,10'd166};
ram[14189] = {-9'd31,10'd169};
ram[14190] = {-9'd28,10'd172};
ram[14191] = {-9'd25,10'd175};
ram[14192] = {-9'd22,10'd179};
ram[14193] = {-9'd19,10'd182};
ram[14194] = {-9'd15,10'd185};
ram[14195] = {-9'd12,10'd188};
ram[14196] = {-9'd9,10'd191};
ram[14197] = {-9'd6,10'd194};
ram[14198] = {-9'd3,10'd197};
ram[14199] = {9'd0,10'd201};
ram[14200] = {9'd3,10'd204};
ram[14201] = {9'd7,10'd207};
ram[14202] = {9'd10,10'd210};
ram[14203] = {9'd13,10'd213};
ram[14204] = {9'd16,10'd216};
ram[14205] = {9'd19,10'd219};
ram[14206] = {9'd22,10'd223};
ram[14207] = {9'd25,10'd226};
ram[14208] = {9'd25,10'd226};
ram[14209] = {9'd29,10'd229};
ram[14210] = {9'd32,10'd232};
ram[14211] = {9'd35,10'd235};
ram[14212] = {9'd38,10'd238};
ram[14213] = {9'd41,10'd241};
ram[14214] = {9'd44,10'd245};
ram[14215] = {9'd47,10'd248};
ram[14216] = {9'd51,10'd251};
ram[14217] = {9'd54,10'd254};
ram[14218] = {9'd57,10'd257};
ram[14219] = {9'd60,10'd260};
ram[14220] = {9'd63,10'd263};
ram[14221] = {9'd66,10'd267};
ram[14222] = {9'd69,10'd270};
ram[14223] = {9'd73,10'd273};
ram[14224] = {9'd76,10'd276};
ram[14225] = {9'd79,10'd279};
ram[14226] = {9'd82,10'd282};
ram[14227] = {9'd85,10'd285};
ram[14228] = {9'd88,10'd289};
ram[14229] = {9'd91,10'd292};
ram[14230] = {9'd95,10'd295};
ram[14231] = {9'd98,10'd298};
ram[14232] = {-9'd99,10'd301};
ram[14233] = {-9'd96,10'd304};
ram[14234] = {-9'd93,10'd307};
ram[14235] = {-9'd90,10'd311};
ram[14236] = {-9'd87,10'd314};
ram[14237] = {-9'd84,10'd317};
ram[14238] = {-9'd81,10'd320};
ram[14239] = {-9'd77,10'd323};
ram[14240] = {-9'd74,10'd326};
ram[14241] = {-9'd71,10'd329};
ram[14242] = {-9'd68,10'd333};
ram[14243] = {-9'd65,10'd336};
ram[14244] = {-9'd62,10'd339};
ram[14245] = {-9'd59,10'd342};
ram[14246] = {-9'd55,10'd345};
ram[14247] = {-9'd52,10'd348};
ram[14248] = {-9'd49,10'd351};
ram[14249] = {-9'd46,10'd354};
ram[14250] = {-9'd43,10'd358};
ram[14251] = {-9'd40,10'd361};
ram[14252] = {-9'd37,10'd364};
ram[14253] = {-9'd33,10'd367};
ram[14254] = {-9'd30,10'd370};
ram[14255] = {-9'd27,10'd373};
ram[14256] = {-9'd24,10'd376};
ram[14257] = {-9'd21,10'd380};
ram[14258] = {-9'd18,10'd383};
ram[14259] = {-9'd15,10'd386};
ram[14260] = {-9'd11,10'd389};
ram[14261] = {-9'd8,10'd392};
ram[14262] = {-9'd5,10'd395};
ram[14263] = {-9'd2,10'd398};
ram[14264] = {9'd1,-10'd399};
ram[14265] = {9'd4,-10'd396};
ram[14266] = {9'd7,-10'd393};
ram[14267] = {9'd10,-10'd390};
ram[14268] = {9'd14,-10'd387};
ram[14269] = {9'd17,-10'd384};
ram[14270] = {9'd20,-10'd381};
ram[14271] = {9'd23,-10'd377};
ram[14272] = {9'd26,-10'd374};
ram[14273] = {9'd29,-10'd371};
ram[14274] = {9'd32,-10'd368};
ram[14275] = {9'd36,-10'd365};
ram[14276] = {9'd39,-10'd362};
ram[14277] = {9'd42,-10'd359};
ram[14278] = {9'd45,-10'd355};
ram[14279] = {9'd48,-10'd352};
ram[14280] = {9'd51,-10'd349};
ram[14281] = {9'd54,-10'd346};
ram[14282] = {9'd58,-10'd343};
ram[14283] = {9'd61,-10'd340};
ram[14284] = {9'd64,-10'd337};
ram[14285] = {9'd67,-10'd334};
ram[14286] = {9'd70,-10'd330};
ram[14287] = {9'd73,-10'd327};
ram[14288] = {9'd76,-10'd324};
ram[14289] = {9'd80,-10'd321};
ram[14290] = {9'd83,-10'd318};
ram[14291] = {9'd86,-10'd315};
ram[14292] = {9'd89,-10'd312};
ram[14293] = {9'd92,-10'd308};
ram[14294] = {9'd95,-10'd305};
ram[14295] = {9'd98,-10'd302};
ram[14296] = {-9'd99,-10'd299};
ram[14297] = {-9'd96,-10'd296};
ram[14298] = {-9'd92,-10'd293};
ram[14299] = {-9'd89,-10'd290};
ram[14300] = {-9'd86,-10'd286};
ram[14301] = {-9'd83,-10'd283};
ram[14302] = {-9'd80,-10'd280};
ram[14303] = {-9'd77,-10'd277};
ram[14304] = {-9'd74,-10'd274};
ram[14305] = {-9'd70,-10'd271};
ram[14306] = {-9'd67,-10'd268};
ram[14307] = {-9'd64,-10'd264};
ram[14308] = {-9'd61,-10'd261};
ram[14309] = {-9'd58,-10'd258};
ram[14310] = {-9'd55,-10'd255};
ram[14311] = {-9'd52,-10'd252};
ram[14312] = {-9'd48,-10'd249};
ram[14313] = {-9'd45,-10'd246};
ram[14314] = {-9'd42,-10'd242};
ram[14315] = {-9'd39,-10'd239};
ram[14316] = {-9'd36,-10'd236};
ram[14317] = {-9'd33,-10'd233};
ram[14318] = {-9'd30,-10'd230};
ram[14319] = {-9'd26,-10'd227};
ram[14320] = {-9'd23,-10'd224};
ram[14321] = {-9'd20,-10'd220};
ram[14322] = {-9'd17,-10'd217};
ram[14323] = {-9'd14,-10'd214};
ram[14324] = {-9'd11,-10'd211};
ram[14325] = {-9'd8,-10'd208};
ram[14326] = {-9'd4,-10'd205};
ram[14327] = {-9'd1,-10'd202};
ram[14328] = {9'd2,-10'd198};
ram[14329] = {9'd5,-10'd195};
ram[14330] = {9'd8,-10'd192};
ram[14331] = {9'd11,-10'd189};
ram[14332] = {9'd14,-10'd186};
ram[14333] = {9'd18,-10'd183};
ram[14334] = {9'd21,-10'd180};
ram[14335] = {9'd24,-10'd176};
ram[14336] = {9'd24,-10'd176};
ram[14337] = {9'd27,-10'd173};
ram[14338] = {9'd30,-10'd170};
ram[14339] = {9'd33,-10'd167};
ram[14340] = {9'd36,-10'd164};
ram[14341] = {9'd40,-10'd161};
ram[14342] = {9'd43,-10'd158};
ram[14343] = {9'd46,-10'd154};
ram[14344] = {9'd49,-10'd151};
ram[14345] = {9'd52,-10'd148};
ram[14346] = {9'd55,-10'd145};
ram[14347] = {9'd58,-10'd142};
ram[14348] = {9'd62,-10'd139};
ram[14349] = {9'd65,-10'd136};
ram[14350] = {9'd68,-10'd132};
ram[14351] = {9'd71,-10'd129};
ram[14352] = {9'd74,-10'd126};
ram[14353] = {9'd77,-10'd123};
ram[14354] = {9'd80,-10'd120};
ram[14355] = {9'd84,-10'd117};
ram[14356] = {9'd87,-10'd114};
ram[14357] = {9'd90,-10'd110};
ram[14358] = {9'd93,-10'd107};
ram[14359] = {9'd96,-10'd104};
ram[14360] = {9'd99,-10'd101};
ram[14361] = {-9'd98,-10'd98};
ram[14362] = {-9'd95,-10'd95};
ram[14363] = {-9'd92,-10'd92};
ram[14364] = {-9'd88,-10'd88};
ram[14365] = {-9'd85,-10'd85};
ram[14366] = {-9'd82,-10'd82};
ram[14367] = {-9'd79,-10'd79};
ram[14368] = {-9'd76,-10'd76};
ram[14369] = {-9'd73,-10'd73};
ram[14370] = {-9'd70,-10'd70};
ram[14371] = {-9'd66,-10'd66};
ram[14372] = {-9'd63,-10'd63};
ram[14373] = {-9'd60,-10'd60};
ram[14374] = {-9'd57,-10'd57};
ram[14375] = {-9'd54,-10'd54};
ram[14376] = {-9'd51,-10'd51};
ram[14377] = {-9'd48,-10'd48};
ram[14378] = {-9'd44,-10'd44};
ram[14379] = {-9'd41,-10'd41};
ram[14380] = {-9'd38,-10'd38};
ram[14381] = {-9'd35,-10'd35};
ram[14382] = {-9'd32,-10'd32};
ram[14383] = {-9'd29,-10'd29};
ram[14384] = {-9'd26,-10'd26};
ram[14385] = {-9'd22,-10'd22};
ram[14386] = {-9'd19,-10'd19};
ram[14387] = {-9'd16,-10'd16};
ram[14388] = {-9'd13,-10'd13};
ram[14389] = {-9'd10,-10'd10};
ram[14390] = {-9'd7,-10'd7};
ram[14391] = {-9'd4,-10'd4};
ram[14392] = {9'd0,10'd0};
ram[14393] = {9'd3,10'd3};
ram[14394] = {9'd6,10'd6};
ram[14395] = {9'd9,10'd9};
ram[14396] = {9'd12,10'd12};
ram[14397] = {9'd15,10'd15};
ram[14398] = {9'd18,10'd18};
ram[14399] = {9'd21,10'd21};
ram[14400] = {9'd25,10'd25};
ram[14401] = {9'd28,10'd28};
ram[14402] = {9'd31,10'd31};
ram[14403] = {9'd34,10'd34};
ram[14404] = {9'd37,10'd37};
ram[14405] = {9'd40,10'd40};
ram[14406] = {9'd43,10'd43};
ram[14407] = {9'd47,10'd47};
ram[14408] = {9'd50,10'd50};
ram[14409] = {9'd53,10'd53};
ram[14410] = {9'd56,10'd56};
ram[14411] = {9'd59,10'd59};
ram[14412] = {9'd62,10'd62};
ram[14413] = {9'd65,10'd65};
ram[14414] = {9'd69,10'd69};
ram[14415] = {9'd72,10'd72};
ram[14416] = {9'd75,10'd75};
ram[14417] = {9'd78,10'd78};
ram[14418] = {9'd81,10'd81};
ram[14419] = {9'd84,10'd84};
ram[14420] = {9'd87,10'd87};
ram[14421] = {9'd91,10'd91};
ram[14422] = {9'd94,10'd94};
ram[14423] = {9'd97,10'd97};
ram[14424] = {-9'd100,10'd100};
ram[14425] = {-9'd97,10'd103};
ram[14426] = {-9'd94,10'd106};
ram[14427] = {-9'd91,10'd109};
ram[14428] = {-9'd88,10'd113};
ram[14429] = {-9'd85,10'd116};
ram[14430] = {-9'd81,10'd119};
ram[14431] = {-9'd78,10'd122};
ram[14432] = {-9'd75,10'd125};
ram[14433] = {-9'd72,10'd128};
ram[14434] = {-9'd69,10'd131};
ram[14435] = {-9'd66,10'd135};
ram[14436] = {-9'd63,10'd138};
ram[14437] = {-9'd59,10'd141};
ram[14438] = {-9'd56,10'd144};
ram[14439] = {-9'd53,10'd147};
ram[14440] = {-9'd50,10'd150};
ram[14441] = {-9'd47,10'd153};
ram[14442] = {-9'd44,10'd157};
ram[14443] = {-9'd41,10'd160};
ram[14444] = {-9'd37,10'd163};
ram[14445] = {-9'd34,10'd166};
ram[14446] = {-9'd31,10'd169};
ram[14447] = {-9'd28,10'd172};
ram[14448] = {-9'd25,10'd175};
ram[14449] = {-9'd22,10'd179};
ram[14450] = {-9'd19,10'd182};
ram[14451] = {-9'd15,10'd185};
ram[14452] = {-9'd12,10'd188};
ram[14453] = {-9'd9,10'd191};
ram[14454] = {-9'd6,10'd194};
ram[14455] = {-9'd3,10'd197};
ram[14456] = {9'd0,10'd201};
ram[14457] = {9'd3,10'd204};
ram[14458] = {9'd7,10'd207};
ram[14459] = {9'd10,10'd210};
ram[14460] = {9'd13,10'd213};
ram[14461] = {9'd16,10'd216};
ram[14462] = {9'd19,10'd219};
ram[14463] = {9'd22,10'd223};
ram[14464] = {9'd22,10'd223};
ram[14465] = {9'd25,10'd226};
ram[14466] = {9'd29,10'd229};
ram[14467] = {9'd32,10'd232};
ram[14468] = {9'd35,10'd235};
ram[14469] = {9'd38,10'd238};
ram[14470] = {9'd41,10'd241};
ram[14471] = {9'd44,10'd245};
ram[14472] = {9'd47,10'd248};
ram[14473] = {9'd51,10'd251};
ram[14474] = {9'd54,10'd254};
ram[14475] = {9'd57,10'd257};
ram[14476] = {9'd60,10'd260};
ram[14477] = {9'd63,10'd263};
ram[14478] = {9'd66,10'd267};
ram[14479] = {9'd69,10'd270};
ram[14480] = {9'd73,10'd273};
ram[14481] = {9'd76,10'd276};
ram[14482] = {9'd79,10'd279};
ram[14483] = {9'd82,10'd282};
ram[14484] = {9'd85,10'd285};
ram[14485] = {9'd88,10'd289};
ram[14486] = {9'd91,10'd292};
ram[14487] = {9'd95,10'd295};
ram[14488] = {9'd98,10'd298};
ram[14489] = {-9'd99,10'd301};
ram[14490] = {-9'd96,10'd304};
ram[14491] = {-9'd93,10'd307};
ram[14492] = {-9'd90,10'd311};
ram[14493] = {-9'd87,10'd314};
ram[14494] = {-9'd84,10'd317};
ram[14495] = {-9'd81,10'd320};
ram[14496] = {-9'd77,10'd323};
ram[14497] = {-9'd74,10'd326};
ram[14498] = {-9'd71,10'd329};
ram[14499] = {-9'd68,10'd333};
ram[14500] = {-9'd65,10'd336};
ram[14501] = {-9'd62,10'd339};
ram[14502] = {-9'd59,10'd342};
ram[14503] = {-9'd55,10'd345};
ram[14504] = {-9'd52,10'd348};
ram[14505] = {-9'd49,10'd351};
ram[14506] = {-9'd46,10'd354};
ram[14507] = {-9'd43,10'd358};
ram[14508] = {-9'd40,10'd361};
ram[14509] = {-9'd37,10'd364};
ram[14510] = {-9'd33,10'd367};
ram[14511] = {-9'd30,10'd370};
ram[14512] = {-9'd27,10'd373};
ram[14513] = {-9'd24,10'd376};
ram[14514] = {-9'd21,10'd380};
ram[14515] = {-9'd18,10'd383};
ram[14516] = {-9'd15,10'd386};
ram[14517] = {-9'd11,10'd389};
ram[14518] = {-9'd8,10'd392};
ram[14519] = {-9'd5,10'd395};
ram[14520] = {-9'd2,10'd398};
ram[14521] = {9'd1,-10'd399};
ram[14522] = {9'd4,-10'd396};
ram[14523] = {9'd7,-10'd393};
ram[14524] = {9'd10,-10'd390};
ram[14525] = {9'd14,-10'd387};
ram[14526] = {9'd17,-10'd384};
ram[14527] = {9'd20,-10'd381};
ram[14528] = {9'd23,-10'd377};
ram[14529] = {9'd26,-10'd374};
ram[14530] = {9'd29,-10'd371};
ram[14531] = {9'd32,-10'd368};
ram[14532] = {9'd36,-10'd365};
ram[14533] = {9'd39,-10'd362};
ram[14534] = {9'd42,-10'd359};
ram[14535] = {9'd45,-10'd355};
ram[14536] = {9'd48,-10'd352};
ram[14537] = {9'd51,-10'd349};
ram[14538] = {9'd54,-10'd346};
ram[14539] = {9'd58,-10'd343};
ram[14540] = {9'd61,-10'd340};
ram[14541] = {9'd64,-10'd337};
ram[14542] = {9'd67,-10'd334};
ram[14543] = {9'd70,-10'd330};
ram[14544] = {9'd73,-10'd327};
ram[14545] = {9'd76,-10'd324};
ram[14546] = {9'd80,-10'd321};
ram[14547] = {9'd83,-10'd318};
ram[14548] = {9'd86,-10'd315};
ram[14549] = {9'd89,-10'd312};
ram[14550] = {9'd92,-10'd308};
ram[14551] = {9'd95,-10'd305};
ram[14552] = {9'd98,-10'd302};
ram[14553] = {-9'd99,-10'd299};
ram[14554] = {-9'd96,-10'd296};
ram[14555] = {-9'd92,-10'd293};
ram[14556] = {-9'd89,-10'd290};
ram[14557] = {-9'd86,-10'd286};
ram[14558] = {-9'd83,-10'd283};
ram[14559] = {-9'd80,-10'd280};
ram[14560] = {-9'd77,-10'd277};
ram[14561] = {-9'd74,-10'd274};
ram[14562] = {-9'd70,-10'd271};
ram[14563] = {-9'd67,-10'd268};
ram[14564] = {-9'd64,-10'd264};
ram[14565] = {-9'd61,-10'd261};
ram[14566] = {-9'd58,-10'd258};
ram[14567] = {-9'd55,-10'd255};
ram[14568] = {-9'd52,-10'd252};
ram[14569] = {-9'd48,-10'd249};
ram[14570] = {-9'd45,-10'd246};
ram[14571] = {-9'd42,-10'd242};
ram[14572] = {-9'd39,-10'd239};
ram[14573] = {-9'd36,-10'd236};
ram[14574] = {-9'd33,-10'd233};
ram[14575] = {-9'd30,-10'd230};
ram[14576] = {-9'd26,-10'd227};
ram[14577] = {-9'd23,-10'd224};
ram[14578] = {-9'd20,-10'd220};
ram[14579] = {-9'd17,-10'd217};
ram[14580] = {-9'd14,-10'd214};
ram[14581] = {-9'd11,-10'd211};
ram[14582] = {-9'd8,-10'd208};
ram[14583] = {-9'd4,-10'd205};
ram[14584] = {-9'd1,-10'd202};
ram[14585] = {9'd2,-10'd198};
ram[14586] = {9'd5,-10'd195};
ram[14587] = {9'd8,-10'd192};
ram[14588] = {9'd11,-10'd189};
ram[14589] = {9'd14,-10'd186};
ram[14590] = {9'd18,-10'd183};
ram[14591] = {9'd21,-10'd180};
ram[14592] = {9'd21,-10'd180};
ram[14593] = {9'd24,-10'd176};
ram[14594] = {9'd27,-10'd173};
ram[14595] = {9'd30,-10'd170};
ram[14596] = {9'd33,-10'd167};
ram[14597] = {9'd36,-10'd164};
ram[14598] = {9'd40,-10'd161};
ram[14599] = {9'd43,-10'd158};
ram[14600] = {9'd46,-10'd154};
ram[14601] = {9'd49,-10'd151};
ram[14602] = {9'd52,-10'd148};
ram[14603] = {9'd55,-10'd145};
ram[14604] = {9'd58,-10'd142};
ram[14605] = {9'd62,-10'd139};
ram[14606] = {9'd65,-10'd136};
ram[14607] = {9'd68,-10'd132};
ram[14608] = {9'd71,-10'd129};
ram[14609] = {9'd74,-10'd126};
ram[14610] = {9'd77,-10'd123};
ram[14611] = {9'd80,-10'd120};
ram[14612] = {9'd84,-10'd117};
ram[14613] = {9'd87,-10'd114};
ram[14614] = {9'd90,-10'd110};
ram[14615] = {9'd93,-10'd107};
ram[14616] = {9'd96,-10'd104};
ram[14617] = {9'd99,-10'd101};
ram[14618] = {-9'd98,-10'd98};
ram[14619] = {-9'd95,-10'd95};
ram[14620] = {-9'd92,-10'd92};
ram[14621] = {-9'd88,-10'd88};
ram[14622] = {-9'd85,-10'd85};
ram[14623] = {-9'd82,-10'd82};
ram[14624] = {-9'd79,-10'd79};
ram[14625] = {-9'd76,-10'd76};
ram[14626] = {-9'd73,-10'd73};
ram[14627] = {-9'd70,-10'd70};
ram[14628] = {-9'd66,-10'd66};
ram[14629] = {-9'd63,-10'd63};
ram[14630] = {-9'd60,-10'd60};
ram[14631] = {-9'd57,-10'd57};
ram[14632] = {-9'd54,-10'd54};
ram[14633] = {-9'd51,-10'd51};
ram[14634] = {-9'd48,-10'd48};
ram[14635] = {-9'd44,-10'd44};
ram[14636] = {-9'd41,-10'd41};
ram[14637] = {-9'd38,-10'd38};
ram[14638] = {-9'd35,-10'd35};
ram[14639] = {-9'd32,-10'd32};
ram[14640] = {-9'd29,-10'd29};
ram[14641] = {-9'd26,-10'd26};
ram[14642] = {-9'd22,-10'd22};
ram[14643] = {-9'd19,-10'd19};
ram[14644] = {-9'd16,-10'd16};
ram[14645] = {-9'd13,-10'd13};
ram[14646] = {-9'd10,-10'd10};
ram[14647] = {-9'd7,-10'd7};
ram[14648] = {-9'd4,-10'd4};
ram[14649] = {9'd0,10'd0};
ram[14650] = {9'd3,10'd3};
ram[14651] = {9'd6,10'd6};
ram[14652] = {9'd9,10'd9};
ram[14653] = {9'd12,10'd12};
ram[14654] = {9'd15,10'd15};
ram[14655] = {9'd18,10'd18};
ram[14656] = {9'd21,10'd21};
ram[14657] = {9'd25,10'd25};
ram[14658] = {9'd28,10'd28};
ram[14659] = {9'd31,10'd31};
ram[14660] = {9'd34,10'd34};
ram[14661] = {9'd37,10'd37};
ram[14662] = {9'd40,10'd40};
ram[14663] = {9'd43,10'd43};
ram[14664] = {9'd47,10'd47};
ram[14665] = {9'd50,10'd50};
ram[14666] = {9'd53,10'd53};
ram[14667] = {9'd56,10'd56};
ram[14668] = {9'd59,10'd59};
ram[14669] = {9'd62,10'd62};
ram[14670] = {9'd65,10'd65};
ram[14671] = {9'd69,10'd69};
ram[14672] = {9'd72,10'd72};
ram[14673] = {9'd75,10'd75};
ram[14674] = {9'd78,10'd78};
ram[14675] = {9'd81,10'd81};
ram[14676] = {9'd84,10'd84};
ram[14677] = {9'd87,10'd87};
ram[14678] = {9'd91,10'd91};
ram[14679] = {9'd94,10'd94};
ram[14680] = {9'd97,10'd97};
ram[14681] = {-9'd100,10'd100};
ram[14682] = {-9'd97,10'd103};
ram[14683] = {-9'd94,10'd106};
ram[14684] = {-9'd91,10'd109};
ram[14685] = {-9'd88,10'd113};
ram[14686] = {-9'd85,10'd116};
ram[14687] = {-9'd81,10'd119};
ram[14688] = {-9'd78,10'd122};
ram[14689] = {-9'd75,10'd125};
ram[14690] = {-9'd72,10'd128};
ram[14691] = {-9'd69,10'd131};
ram[14692] = {-9'd66,10'd135};
ram[14693] = {-9'd63,10'd138};
ram[14694] = {-9'd59,10'd141};
ram[14695] = {-9'd56,10'd144};
ram[14696] = {-9'd53,10'd147};
ram[14697] = {-9'd50,10'd150};
ram[14698] = {-9'd47,10'd153};
ram[14699] = {-9'd44,10'd157};
ram[14700] = {-9'd41,10'd160};
ram[14701] = {-9'd37,10'd163};
ram[14702] = {-9'd34,10'd166};
ram[14703] = {-9'd31,10'd169};
ram[14704] = {-9'd28,10'd172};
ram[14705] = {-9'd25,10'd175};
ram[14706] = {-9'd22,10'd179};
ram[14707] = {-9'd19,10'd182};
ram[14708] = {-9'd15,10'd185};
ram[14709] = {-9'd12,10'd188};
ram[14710] = {-9'd9,10'd191};
ram[14711] = {-9'd6,10'd194};
ram[14712] = {-9'd3,10'd197};
ram[14713] = {9'd0,10'd201};
ram[14714] = {9'd3,10'd204};
ram[14715] = {9'd7,10'd207};
ram[14716] = {9'd10,10'd210};
ram[14717] = {9'd13,10'd213};
ram[14718] = {9'd16,10'd216};
ram[14719] = {9'd19,10'd219};
ram[14720] = {9'd19,10'd219};
ram[14721] = {9'd22,10'd223};
ram[14722] = {9'd25,10'd226};
ram[14723] = {9'd29,10'd229};
ram[14724] = {9'd32,10'd232};
ram[14725] = {9'd35,10'd235};
ram[14726] = {9'd38,10'd238};
ram[14727] = {9'd41,10'd241};
ram[14728] = {9'd44,10'd245};
ram[14729] = {9'd47,10'd248};
ram[14730] = {9'd51,10'd251};
ram[14731] = {9'd54,10'd254};
ram[14732] = {9'd57,10'd257};
ram[14733] = {9'd60,10'd260};
ram[14734] = {9'd63,10'd263};
ram[14735] = {9'd66,10'd267};
ram[14736] = {9'd69,10'd270};
ram[14737] = {9'd73,10'd273};
ram[14738] = {9'd76,10'd276};
ram[14739] = {9'd79,10'd279};
ram[14740] = {9'd82,10'd282};
ram[14741] = {9'd85,10'd285};
ram[14742] = {9'd88,10'd289};
ram[14743] = {9'd91,10'd292};
ram[14744] = {9'd95,10'd295};
ram[14745] = {9'd98,10'd298};
ram[14746] = {-9'd99,10'd301};
ram[14747] = {-9'd96,10'd304};
ram[14748] = {-9'd93,10'd307};
ram[14749] = {-9'd90,10'd311};
ram[14750] = {-9'd87,10'd314};
ram[14751] = {-9'd84,10'd317};
ram[14752] = {-9'd81,10'd320};
ram[14753] = {-9'd77,10'd323};
ram[14754] = {-9'd74,10'd326};
ram[14755] = {-9'd71,10'd329};
ram[14756] = {-9'd68,10'd333};
ram[14757] = {-9'd65,10'd336};
ram[14758] = {-9'd62,10'd339};
ram[14759] = {-9'd59,10'd342};
ram[14760] = {-9'd55,10'd345};
ram[14761] = {-9'd52,10'd348};
ram[14762] = {-9'd49,10'd351};
ram[14763] = {-9'd46,10'd354};
ram[14764] = {-9'd43,10'd358};
ram[14765] = {-9'd40,10'd361};
ram[14766] = {-9'd37,10'd364};
ram[14767] = {-9'd33,10'd367};
ram[14768] = {-9'd30,10'd370};
ram[14769] = {-9'd27,10'd373};
ram[14770] = {-9'd24,10'd376};
ram[14771] = {-9'd21,10'd380};
ram[14772] = {-9'd18,10'd383};
ram[14773] = {-9'd15,10'd386};
ram[14774] = {-9'd11,10'd389};
ram[14775] = {-9'd8,10'd392};
ram[14776] = {-9'd5,10'd395};
ram[14777] = {-9'd2,10'd398};
ram[14778] = {9'd1,-10'd399};
ram[14779] = {9'd4,-10'd396};
ram[14780] = {9'd7,-10'd393};
ram[14781] = {9'd10,-10'd390};
ram[14782] = {9'd14,-10'd387};
ram[14783] = {9'd17,-10'd384};
ram[14784] = {9'd20,-10'd381};
ram[14785] = {9'd23,-10'd377};
ram[14786] = {9'd26,-10'd374};
ram[14787] = {9'd29,-10'd371};
ram[14788] = {9'd32,-10'd368};
ram[14789] = {9'd36,-10'd365};
ram[14790] = {9'd39,-10'd362};
ram[14791] = {9'd42,-10'd359};
ram[14792] = {9'd45,-10'd355};
ram[14793] = {9'd48,-10'd352};
ram[14794] = {9'd51,-10'd349};
ram[14795] = {9'd54,-10'd346};
ram[14796] = {9'd58,-10'd343};
ram[14797] = {9'd61,-10'd340};
ram[14798] = {9'd64,-10'd337};
ram[14799] = {9'd67,-10'd334};
ram[14800] = {9'd70,-10'd330};
ram[14801] = {9'd73,-10'd327};
ram[14802] = {9'd76,-10'd324};
ram[14803] = {9'd80,-10'd321};
ram[14804] = {9'd83,-10'd318};
ram[14805] = {9'd86,-10'd315};
ram[14806] = {9'd89,-10'd312};
ram[14807] = {9'd92,-10'd308};
ram[14808] = {9'd95,-10'd305};
ram[14809] = {9'd98,-10'd302};
ram[14810] = {-9'd99,-10'd299};
ram[14811] = {-9'd96,-10'd296};
ram[14812] = {-9'd92,-10'd293};
ram[14813] = {-9'd89,-10'd290};
ram[14814] = {-9'd86,-10'd286};
ram[14815] = {-9'd83,-10'd283};
ram[14816] = {-9'd80,-10'd280};
ram[14817] = {-9'd77,-10'd277};
ram[14818] = {-9'd74,-10'd274};
ram[14819] = {-9'd70,-10'd271};
ram[14820] = {-9'd67,-10'd268};
ram[14821] = {-9'd64,-10'd264};
ram[14822] = {-9'd61,-10'd261};
ram[14823] = {-9'd58,-10'd258};
ram[14824] = {-9'd55,-10'd255};
ram[14825] = {-9'd52,-10'd252};
ram[14826] = {-9'd48,-10'd249};
ram[14827] = {-9'd45,-10'd246};
ram[14828] = {-9'd42,-10'd242};
ram[14829] = {-9'd39,-10'd239};
ram[14830] = {-9'd36,-10'd236};
ram[14831] = {-9'd33,-10'd233};
ram[14832] = {-9'd30,-10'd230};
ram[14833] = {-9'd26,-10'd227};
ram[14834] = {-9'd23,-10'd224};
ram[14835] = {-9'd20,-10'd220};
ram[14836] = {-9'd17,-10'd217};
ram[14837] = {-9'd14,-10'd214};
ram[14838] = {-9'd11,-10'd211};
ram[14839] = {-9'd8,-10'd208};
ram[14840] = {-9'd4,-10'd205};
ram[14841] = {-9'd1,-10'd202};
ram[14842] = {9'd2,-10'd198};
ram[14843] = {9'd5,-10'd195};
ram[14844] = {9'd8,-10'd192};
ram[14845] = {9'd11,-10'd189};
ram[14846] = {9'd14,-10'd186};
ram[14847] = {9'd18,-10'd183};
ram[14848] = {9'd18,-10'd183};
ram[14849] = {9'd21,-10'd180};
ram[14850] = {9'd24,-10'd176};
ram[14851] = {9'd27,-10'd173};
ram[14852] = {9'd30,-10'd170};
ram[14853] = {9'd33,-10'd167};
ram[14854] = {9'd36,-10'd164};
ram[14855] = {9'd40,-10'd161};
ram[14856] = {9'd43,-10'd158};
ram[14857] = {9'd46,-10'd154};
ram[14858] = {9'd49,-10'd151};
ram[14859] = {9'd52,-10'd148};
ram[14860] = {9'd55,-10'd145};
ram[14861] = {9'd58,-10'd142};
ram[14862] = {9'd62,-10'd139};
ram[14863] = {9'd65,-10'd136};
ram[14864] = {9'd68,-10'd132};
ram[14865] = {9'd71,-10'd129};
ram[14866] = {9'd74,-10'd126};
ram[14867] = {9'd77,-10'd123};
ram[14868] = {9'd80,-10'd120};
ram[14869] = {9'd84,-10'd117};
ram[14870] = {9'd87,-10'd114};
ram[14871] = {9'd90,-10'd110};
ram[14872] = {9'd93,-10'd107};
ram[14873] = {9'd96,-10'd104};
ram[14874] = {9'd99,-10'd101};
ram[14875] = {-9'd98,-10'd98};
ram[14876] = {-9'd95,-10'd95};
ram[14877] = {-9'd92,-10'd92};
ram[14878] = {-9'd88,-10'd88};
ram[14879] = {-9'd85,-10'd85};
ram[14880] = {-9'd82,-10'd82};
ram[14881] = {-9'd79,-10'd79};
ram[14882] = {-9'd76,-10'd76};
ram[14883] = {-9'd73,-10'd73};
ram[14884] = {-9'd70,-10'd70};
ram[14885] = {-9'd66,-10'd66};
ram[14886] = {-9'd63,-10'd63};
ram[14887] = {-9'd60,-10'd60};
ram[14888] = {-9'd57,-10'd57};
ram[14889] = {-9'd54,-10'd54};
ram[14890] = {-9'd51,-10'd51};
ram[14891] = {-9'd48,-10'd48};
ram[14892] = {-9'd44,-10'd44};
ram[14893] = {-9'd41,-10'd41};
ram[14894] = {-9'd38,-10'd38};
ram[14895] = {-9'd35,-10'd35};
ram[14896] = {-9'd32,-10'd32};
ram[14897] = {-9'd29,-10'd29};
ram[14898] = {-9'd26,-10'd26};
ram[14899] = {-9'd22,-10'd22};
ram[14900] = {-9'd19,-10'd19};
ram[14901] = {-9'd16,-10'd16};
ram[14902] = {-9'd13,-10'd13};
ram[14903] = {-9'd10,-10'd10};
ram[14904] = {-9'd7,-10'd7};
ram[14905] = {-9'd4,-10'd4};
ram[14906] = {9'd0,10'd0};
ram[14907] = {9'd3,10'd3};
ram[14908] = {9'd6,10'd6};
ram[14909] = {9'd9,10'd9};
ram[14910] = {9'd12,10'd12};
ram[14911] = {9'd15,10'd15};
ram[14912] = {9'd18,10'd18};
ram[14913] = {9'd21,10'd21};
ram[14914] = {9'd25,10'd25};
ram[14915] = {9'd28,10'd28};
ram[14916] = {9'd31,10'd31};
ram[14917] = {9'd34,10'd34};
ram[14918] = {9'd37,10'd37};
ram[14919] = {9'd40,10'd40};
ram[14920] = {9'd43,10'd43};
ram[14921] = {9'd47,10'd47};
ram[14922] = {9'd50,10'd50};
ram[14923] = {9'd53,10'd53};
ram[14924] = {9'd56,10'd56};
ram[14925] = {9'd59,10'd59};
ram[14926] = {9'd62,10'd62};
ram[14927] = {9'd65,10'd65};
ram[14928] = {9'd69,10'd69};
ram[14929] = {9'd72,10'd72};
ram[14930] = {9'd75,10'd75};
ram[14931] = {9'd78,10'd78};
ram[14932] = {9'd81,10'd81};
ram[14933] = {9'd84,10'd84};
ram[14934] = {9'd87,10'd87};
ram[14935] = {9'd91,10'd91};
ram[14936] = {9'd94,10'd94};
ram[14937] = {9'd97,10'd97};
ram[14938] = {-9'd100,10'd100};
ram[14939] = {-9'd97,10'd103};
ram[14940] = {-9'd94,10'd106};
ram[14941] = {-9'd91,10'd109};
ram[14942] = {-9'd88,10'd113};
ram[14943] = {-9'd85,10'd116};
ram[14944] = {-9'd81,10'd119};
ram[14945] = {-9'd78,10'd122};
ram[14946] = {-9'd75,10'd125};
ram[14947] = {-9'd72,10'd128};
ram[14948] = {-9'd69,10'd131};
ram[14949] = {-9'd66,10'd135};
ram[14950] = {-9'd63,10'd138};
ram[14951] = {-9'd59,10'd141};
ram[14952] = {-9'd56,10'd144};
ram[14953] = {-9'd53,10'd147};
ram[14954] = {-9'd50,10'd150};
ram[14955] = {-9'd47,10'd153};
ram[14956] = {-9'd44,10'd157};
ram[14957] = {-9'd41,10'd160};
ram[14958] = {-9'd37,10'd163};
ram[14959] = {-9'd34,10'd166};
ram[14960] = {-9'd31,10'd169};
ram[14961] = {-9'd28,10'd172};
ram[14962] = {-9'd25,10'd175};
ram[14963] = {-9'd22,10'd179};
ram[14964] = {-9'd19,10'd182};
ram[14965] = {-9'd15,10'd185};
ram[14966] = {-9'd12,10'd188};
ram[14967] = {-9'd9,10'd191};
ram[14968] = {-9'd6,10'd194};
ram[14969] = {-9'd3,10'd197};
ram[14970] = {9'd0,10'd201};
ram[14971] = {9'd3,10'd204};
ram[14972] = {9'd7,10'd207};
ram[14973] = {9'd10,10'd210};
ram[14974] = {9'd13,10'd213};
ram[14975] = {9'd16,10'd216};
ram[14976] = {9'd16,10'd216};
ram[14977] = {9'd19,10'd219};
ram[14978] = {9'd22,10'd223};
ram[14979] = {9'd25,10'd226};
ram[14980] = {9'd29,10'd229};
ram[14981] = {9'd32,10'd232};
ram[14982] = {9'd35,10'd235};
ram[14983] = {9'd38,10'd238};
ram[14984] = {9'd41,10'd241};
ram[14985] = {9'd44,10'd245};
ram[14986] = {9'd47,10'd248};
ram[14987] = {9'd51,10'd251};
ram[14988] = {9'd54,10'd254};
ram[14989] = {9'd57,10'd257};
ram[14990] = {9'd60,10'd260};
ram[14991] = {9'd63,10'd263};
ram[14992] = {9'd66,10'd267};
ram[14993] = {9'd69,10'd270};
ram[14994] = {9'd73,10'd273};
ram[14995] = {9'd76,10'd276};
ram[14996] = {9'd79,10'd279};
ram[14997] = {9'd82,10'd282};
ram[14998] = {9'd85,10'd285};
ram[14999] = {9'd88,10'd289};
ram[15000] = {9'd91,10'd292};
ram[15001] = {9'd95,10'd295};
ram[15002] = {9'd98,10'd298};
ram[15003] = {-9'd99,10'd301};
ram[15004] = {-9'd96,10'd304};
ram[15005] = {-9'd93,10'd307};
ram[15006] = {-9'd90,10'd311};
ram[15007] = {-9'd87,10'd314};
ram[15008] = {-9'd84,10'd317};
ram[15009] = {-9'd81,10'd320};
ram[15010] = {-9'd77,10'd323};
ram[15011] = {-9'd74,10'd326};
ram[15012] = {-9'd71,10'd329};
ram[15013] = {-9'd68,10'd333};
ram[15014] = {-9'd65,10'd336};
ram[15015] = {-9'd62,10'd339};
ram[15016] = {-9'd59,10'd342};
ram[15017] = {-9'd55,10'd345};
ram[15018] = {-9'd52,10'd348};
ram[15019] = {-9'd49,10'd351};
ram[15020] = {-9'd46,10'd354};
ram[15021] = {-9'd43,10'd358};
ram[15022] = {-9'd40,10'd361};
ram[15023] = {-9'd37,10'd364};
ram[15024] = {-9'd33,10'd367};
ram[15025] = {-9'd30,10'd370};
ram[15026] = {-9'd27,10'd373};
ram[15027] = {-9'd24,10'd376};
ram[15028] = {-9'd21,10'd380};
ram[15029] = {-9'd18,10'd383};
ram[15030] = {-9'd15,10'd386};
ram[15031] = {-9'd11,10'd389};
ram[15032] = {-9'd8,10'd392};
ram[15033] = {-9'd5,10'd395};
ram[15034] = {-9'd2,10'd398};
ram[15035] = {9'd1,-10'd399};
ram[15036] = {9'd4,-10'd396};
ram[15037] = {9'd7,-10'd393};
ram[15038] = {9'd10,-10'd390};
ram[15039] = {9'd14,-10'd387};
ram[15040] = {9'd17,-10'd384};
ram[15041] = {9'd20,-10'd381};
ram[15042] = {9'd23,-10'd377};
ram[15043] = {9'd26,-10'd374};
ram[15044] = {9'd29,-10'd371};
ram[15045] = {9'd32,-10'd368};
ram[15046] = {9'd36,-10'd365};
ram[15047] = {9'd39,-10'd362};
ram[15048] = {9'd42,-10'd359};
ram[15049] = {9'd45,-10'd355};
ram[15050] = {9'd48,-10'd352};
ram[15051] = {9'd51,-10'd349};
ram[15052] = {9'd54,-10'd346};
ram[15053] = {9'd58,-10'd343};
ram[15054] = {9'd61,-10'd340};
ram[15055] = {9'd64,-10'd337};
ram[15056] = {9'd67,-10'd334};
ram[15057] = {9'd70,-10'd330};
ram[15058] = {9'd73,-10'd327};
ram[15059] = {9'd76,-10'd324};
ram[15060] = {9'd80,-10'd321};
ram[15061] = {9'd83,-10'd318};
ram[15062] = {9'd86,-10'd315};
ram[15063] = {9'd89,-10'd312};
ram[15064] = {9'd92,-10'd308};
ram[15065] = {9'd95,-10'd305};
ram[15066] = {9'd98,-10'd302};
ram[15067] = {-9'd99,-10'd299};
ram[15068] = {-9'd96,-10'd296};
ram[15069] = {-9'd92,-10'd293};
ram[15070] = {-9'd89,-10'd290};
ram[15071] = {-9'd86,-10'd286};
ram[15072] = {-9'd83,-10'd283};
ram[15073] = {-9'd80,-10'd280};
ram[15074] = {-9'd77,-10'd277};
ram[15075] = {-9'd74,-10'd274};
ram[15076] = {-9'd70,-10'd271};
ram[15077] = {-9'd67,-10'd268};
ram[15078] = {-9'd64,-10'd264};
ram[15079] = {-9'd61,-10'd261};
ram[15080] = {-9'd58,-10'd258};
ram[15081] = {-9'd55,-10'd255};
ram[15082] = {-9'd52,-10'd252};
ram[15083] = {-9'd48,-10'd249};
ram[15084] = {-9'd45,-10'd246};
ram[15085] = {-9'd42,-10'd242};
ram[15086] = {-9'd39,-10'd239};
ram[15087] = {-9'd36,-10'd236};
ram[15088] = {-9'd33,-10'd233};
ram[15089] = {-9'd30,-10'd230};
ram[15090] = {-9'd26,-10'd227};
ram[15091] = {-9'd23,-10'd224};
ram[15092] = {-9'd20,-10'd220};
ram[15093] = {-9'd17,-10'd217};
ram[15094] = {-9'd14,-10'd214};
ram[15095] = {-9'd11,-10'd211};
ram[15096] = {-9'd8,-10'd208};
ram[15097] = {-9'd4,-10'd205};
ram[15098] = {-9'd1,-10'd202};
ram[15099] = {9'd2,-10'd198};
ram[15100] = {9'd5,-10'd195};
ram[15101] = {9'd8,-10'd192};
ram[15102] = {9'd11,-10'd189};
ram[15103] = {9'd14,-10'd186};
ram[15104] = {9'd14,-10'd186};
ram[15105] = {9'd18,-10'd183};
ram[15106] = {9'd21,-10'd180};
ram[15107] = {9'd24,-10'd176};
ram[15108] = {9'd27,-10'd173};
ram[15109] = {9'd30,-10'd170};
ram[15110] = {9'd33,-10'd167};
ram[15111] = {9'd36,-10'd164};
ram[15112] = {9'd40,-10'd161};
ram[15113] = {9'd43,-10'd158};
ram[15114] = {9'd46,-10'd154};
ram[15115] = {9'd49,-10'd151};
ram[15116] = {9'd52,-10'd148};
ram[15117] = {9'd55,-10'd145};
ram[15118] = {9'd58,-10'd142};
ram[15119] = {9'd62,-10'd139};
ram[15120] = {9'd65,-10'd136};
ram[15121] = {9'd68,-10'd132};
ram[15122] = {9'd71,-10'd129};
ram[15123] = {9'd74,-10'd126};
ram[15124] = {9'd77,-10'd123};
ram[15125] = {9'd80,-10'd120};
ram[15126] = {9'd84,-10'd117};
ram[15127] = {9'd87,-10'd114};
ram[15128] = {9'd90,-10'd110};
ram[15129] = {9'd93,-10'd107};
ram[15130] = {9'd96,-10'd104};
ram[15131] = {9'd99,-10'd101};
ram[15132] = {-9'd98,-10'd98};
ram[15133] = {-9'd95,-10'd95};
ram[15134] = {-9'd92,-10'd92};
ram[15135] = {-9'd88,-10'd88};
ram[15136] = {-9'd85,-10'd85};
ram[15137] = {-9'd82,-10'd82};
ram[15138] = {-9'd79,-10'd79};
ram[15139] = {-9'd76,-10'd76};
ram[15140] = {-9'd73,-10'd73};
ram[15141] = {-9'd70,-10'd70};
ram[15142] = {-9'd66,-10'd66};
ram[15143] = {-9'd63,-10'd63};
ram[15144] = {-9'd60,-10'd60};
ram[15145] = {-9'd57,-10'd57};
ram[15146] = {-9'd54,-10'd54};
ram[15147] = {-9'd51,-10'd51};
ram[15148] = {-9'd48,-10'd48};
ram[15149] = {-9'd44,-10'd44};
ram[15150] = {-9'd41,-10'd41};
ram[15151] = {-9'd38,-10'd38};
ram[15152] = {-9'd35,-10'd35};
ram[15153] = {-9'd32,-10'd32};
ram[15154] = {-9'd29,-10'd29};
ram[15155] = {-9'd26,-10'd26};
ram[15156] = {-9'd22,-10'd22};
ram[15157] = {-9'd19,-10'd19};
ram[15158] = {-9'd16,-10'd16};
ram[15159] = {-9'd13,-10'd13};
ram[15160] = {-9'd10,-10'd10};
ram[15161] = {-9'd7,-10'd7};
ram[15162] = {-9'd4,-10'd4};
ram[15163] = {9'd0,10'd0};
ram[15164] = {9'd3,10'd3};
ram[15165] = {9'd6,10'd6};
ram[15166] = {9'd9,10'd9};
ram[15167] = {9'd12,10'd12};
ram[15168] = {9'd15,10'd15};
ram[15169] = {9'd18,10'd18};
ram[15170] = {9'd21,10'd21};
ram[15171] = {9'd25,10'd25};
ram[15172] = {9'd28,10'd28};
ram[15173] = {9'd31,10'd31};
ram[15174] = {9'd34,10'd34};
ram[15175] = {9'd37,10'd37};
ram[15176] = {9'd40,10'd40};
ram[15177] = {9'd43,10'd43};
ram[15178] = {9'd47,10'd47};
ram[15179] = {9'd50,10'd50};
ram[15180] = {9'd53,10'd53};
ram[15181] = {9'd56,10'd56};
ram[15182] = {9'd59,10'd59};
ram[15183] = {9'd62,10'd62};
ram[15184] = {9'd65,10'd65};
ram[15185] = {9'd69,10'd69};
ram[15186] = {9'd72,10'd72};
ram[15187] = {9'd75,10'd75};
ram[15188] = {9'd78,10'd78};
ram[15189] = {9'd81,10'd81};
ram[15190] = {9'd84,10'd84};
ram[15191] = {9'd87,10'd87};
ram[15192] = {9'd91,10'd91};
ram[15193] = {9'd94,10'd94};
ram[15194] = {9'd97,10'd97};
ram[15195] = {-9'd100,10'd100};
ram[15196] = {-9'd97,10'd103};
ram[15197] = {-9'd94,10'd106};
ram[15198] = {-9'd91,10'd109};
ram[15199] = {-9'd88,10'd113};
ram[15200] = {-9'd85,10'd116};
ram[15201] = {-9'd81,10'd119};
ram[15202] = {-9'd78,10'd122};
ram[15203] = {-9'd75,10'd125};
ram[15204] = {-9'd72,10'd128};
ram[15205] = {-9'd69,10'd131};
ram[15206] = {-9'd66,10'd135};
ram[15207] = {-9'd63,10'd138};
ram[15208] = {-9'd59,10'd141};
ram[15209] = {-9'd56,10'd144};
ram[15210] = {-9'd53,10'd147};
ram[15211] = {-9'd50,10'd150};
ram[15212] = {-9'd47,10'd153};
ram[15213] = {-9'd44,10'd157};
ram[15214] = {-9'd41,10'd160};
ram[15215] = {-9'd37,10'd163};
ram[15216] = {-9'd34,10'd166};
ram[15217] = {-9'd31,10'd169};
ram[15218] = {-9'd28,10'd172};
ram[15219] = {-9'd25,10'd175};
ram[15220] = {-9'd22,10'd179};
ram[15221] = {-9'd19,10'd182};
ram[15222] = {-9'd15,10'd185};
ram[15223] = {-9'd12,10'd188};
ram[15224] = {-9'd9,10'd191};
ram[15225] = {-9'd6,10'd194};
ram[15226] = {-9'd3,10'd197};
ram[15227] = {9'd0,10'd201};
ram[15228] = {9'd3,10'd204};
ram[15229] = {9'd7,10'd207};
ram[15230] = {9'd10,10'd210};
ram[15231] = {9'd13,10'd213};
ram[15232] = {9'd13,10'd213};
ram[15233] = {9'd16,10'd216};
ram[15234] = {9'd19,10'd219};
ram[15235] = {9'd22,10'd223};
ram[15236] = {9'd25,10'd226};
ram[15237] = {9'd29,10'd229};
ram[15238] = {9'd32,10'd232};
ram[15239] = {9'd35,10'd235};
ram[15240] = {9'd38,10'd238};
ram[15241] = {9'd41,10'd241};
ram[15242] = {9'd44,10'd245};
ram[15243] = {9'd47,10'd248};
ram[15244] = {9'd51,10'd251};
ram[15245] = {9'd54,10'd254};
ram[15246] = {9'd57,10'd257};
ram[15247] = {9'd60,10'd260};
ram[15248] = {9'd63,10'd263};
ram[15249] = {9'd66,10'd267};
ram[15250] = {9'd69,10'd270};
ram[15251] = {9'd73,10'd273};
ram[15252] = {9'd76,10'd276};
ram[15253] = {9'd79,10'd279};
ram[15254] = {9'd82,10'd282};
ram[15255] = {9'd85,10'd285};
ram[15256] = {9'd88,10'd289};
ram[15257] = {9'd91,10'd292};
ram[15258] = {9'd95,10'd295};
ram[15259] = {9'd98,10'd298};
ram[15260] = {-9'd99,10'd301};
ram[15261] = {-9'd96,10'd304};
ram[15262] = {-9'd93,10'd307};
ram[15263] = {-9'd90,10'd311};
ram[15264] = {-9'd87,10'd314};
ram[15265] = {-9'd84,10'd317};
ram[15266] = {-9'd81,10'd320};
ram[15267] = {-9'd77,10'd323};
ram[15268] = {-9'd74,10'd326};
ram[15269] = {-9'd71,10'd329};
ram[15270] = {-9'd68,10'd333};
ram[15271] = {-9'd65,10'd336};
ram[15272] = {-9'd62,10'd339};
ram[15273] = {-9'd59,10'd342};
ram[15274] = {-9'd55,10'd345};
ram[15275] = {-9'd52,10'd348};
ram[15276] = {-9'd49,10'd351};
ram[15277] = {-9'd46,10'd354};
ram[15278] = {-9'd43,10'd358};
ram[15279] = {-9'd40,10'd361};
ram[15280] = {-9'd37,10'd364};
ram[15281] = {-9'd33,10'd367};
ram[15282] = {-9'd30,10'd370};
ram[15283] = {-9'd27,10'd373};
ram[15284] = {-9'd24,10'd376};
ram[15285] = {-9'd21,10'd380};
ram[15286] = {-9'd18,10'd383};
ram[15287] = {-9'd15,10'd386};
ram[15288] = {-9'd11,10'd389};
ram[15289] = {-9'd8,10'd392};
ram[15290] = {-9'd5,10'd395};
ram[15291] = {-9'd2,10'd398};
ram[15292] = {9'd1,-10'd399};
ram[15293] = {9'd4,-10'd396};
ram[15294] = {9'd7,-10'd393};
ram[15295] = {9'd10,-10'd390};
ram[15296] = {9'd14,-10'd387};
ram[15297] = {9'd17,-10'd384};
ram[15298] = {9'd20,-10'd381};
ram[15299] = {9'd23,-10'd377};
ram[15300] = {9'd26,-10'd374};
ram[15301] = {9'd29,-10'd371};
ram[15302] = {9'd32,-10'd368};
ram[15303] = {9'd36,-10'd365};
ram[15304] = {9'd39,-10'd362};
ram[15305] = {9'd42,-10'd359};
ram[15306] = {9'd45,-10'd355};
ram[15307] = {9'd48,-10'd352};
ram[15308] = {9'd51,-10'd349};
ram[15309] = {9'd54,-10'd346};
ram[15310] = {9'd58,-10'd343};
ram[15311] = {9'd61,-10'd340};
ram[15312] = {9'd64,-10'd337};
ram[15313] = {9'd67,-10'd334};
ram[15314] = {9'd70,-10'd330};
ram[15315] = {9'd73,-10'd327};
ram[15316] = {9'd76,-10'd324};
ram[15317] = {9'd80,-10'd321};
ram[15318] = {9'd83,-10'd318};
ram[15319] = {9'd86,-10'd315};
ram[15320] = {9'd89,-10'd312};
ram[15321] = {9'd92,-10'd308};
ram[15322] = {9'd95,-10'd305};
ram[15323] = {9'd98,-10'd302};
ram[15324] = {-9'd99,-10'd299};
ram[15325] = {-9'd96,-10'd296};
ram[15326] = {-9'd92,-10'd293};
ram[15327] = {-9'd89,-10'd290};
ram[15328] = {-9'd86,-10'd286};
ram[15329] = {-9'd83,-10'd283};
ram[15330] = {-9'd80,-10'd280};
ram[15331] = {-9'd77,-10'd277};
ram[15332] = {-9'd74,-10'd274};
ram[15333] = {-9'd70,-10'd271};
ram[15334] = {-9'd67,-10'd268};
ram[15335] = {-9'd64,-10'd264};
ram[15336] = {-9'd61,-10'd261};
ram[15337] = {-9'd58,-10'd258};
ram[15338] = {-9'd55,-10'd255};
ram[15339] = {-9'd52,-10'd252};
ram[15340] = {-9'd48,-10'd249};
ram[15341] = {-9'd45,-10'd246};
ram[15342] = {-9'd42,-10'd242};
ram[15343] = {-9'd39,-10'd239};
ram[15344] = {-9'd36,-10'd236};
ram[15345] = {-9'd33,-10'd233};
ram[15346] = {-9'd30,-10'd230};
ram[15347] = {-9'd26,-10'd227};
ram[15348] = {-9'd23,-10'd224};
ram[15349] = {-9'd20,-10'd220};
ram[15350] = {-9'd17,-10'd217};
ram[15351] = {-9'd14,-10'd214};
ram[15352] = {-9'd11,-10'd211};
ram[15353] = {-9'd8,-10'd208};
ram[15354] = {-9'd4,-10'd205};
ram[15355] = {-9'd1,-10'd202};
ram[15356] = {9'd2,-10'd198};
ram[15357] = {9'd5,-10'd195};
ram[15358] = {9'd8,-10'd192};
ram[15359] = {9'd11,-10'd189};
ram[15360] = {9'd11,-10'd189};
ram[15361] = {9'd14,-10'd186};
ram[15362] = {9'd18,-10'd183};
ram[15363] = {9'd21,-10'd180};
ram[15364] = {9'd24,-10'd176};
ram[15365] = {9'd27,-10'd173};
ram[15366] = {9'd30,-10'd170};
ram[15367] = {9'd33,-10'd167};
ram[15368] = {9'd36,-10'd164};
ram[15369] = {9'd40,-10'd161};
ram[15370] = {9'd43,-10'd158};
ram[15371] = {9'd46,-10'd154};
ram[15372] = {9'd49,-10'd151};
ram[15373] = {9'd52,-10'd148};
ram[15374] = {9'd55,-10'd145};
ram[15375] = {9'd58,-10'd142};
ram[15376] = {9'd62,-10'd139};
ram[15377] = {9'd65,-10'd136};
ram[15378] = {9'd68,-10'd132};
ram[15379] = {9'd71,-10'd129};
ram[15380] = {9'd74,-10'd126};
ram[15381] = {9'd77,-10'd123};
ram[15382] = {9'd80,-10'd120};
ram[15383] = {9'd84,-10'd117};
ram[15384] = {9'd87,-10'd114};
ram[15385] = {9'd90,-10'd110};
ram[15386] = {9'd93,-10'd107};
ram[15387] = {9'd96,-10'd104};
ram[15388] = {9'd99,-10'd101};
ram[15389] = {-9'd98,-10'd98};
ram[15390] = {-9'd95,-10'd95};
ram[15391] = {-9'd92,-10'd92};
ram[15392] = {-9'd88,-10'd88};
ram[15393] = {-9'd85,-10'd85};
ram[15394] = {-9'd82,-10'd82};
ram[15395] = {-9'd79,-10'd79};
ram[15396] = {-9'd76,-10'd76};
ram[15397] = {-9'd73,-10'd73};
ram[15398] = {-9'd70,-10'd70};
ram[15399] = {-9'd66,-10'd66};
ram[15400] = {-9'd63,-10'd63};
ram[15401] = {-9'd60,-10'd60};
ram[15402] = {-9'd57,-10'd57};
ram[15403] = {-9'd54,-10'd54};
ram[15404] = {-9'd51,-10'd51};
ram[15405] = {-9'd48,-10'd48};
ram[15406] = {-9'd44,-10'd44};
ram[15407] = {-9'd41,-10'd41};
ram[15408] = {-9'd38,-10'd38};
ram[15409] = {-9'd35,-10'd35};
ram[15410] = {-9'd32,-10'd32};
ram[15411] = {-9'd29,-10'd29};
ram[15412] = {-9'd26,-10'd26};
ram[15413] = {-9'd22,-10'd22};
ram[15414] = {-9'd19,-10'd19};
ram[15415] = {-9'd16,-10'd16};
ram[15416] = {-9'd13,-10'd13};
ram[15417] = {-9'd10,-10'd10};
ram[15418] = {-9'd7,-10'd7};
ram[15419] = {-9'd4,-10'd4};
ram[15420] = {9'd0,10'd0};
ram[15421] = {9'd3,10'd3};
ram[15422] = {9'd6,10'd6};
ram[15423] = {9'd9,10'd9};
ram[15424] = {9'd12,10'd12};
ram[15425] = {9'd15,10'd15};
ram[15426] = {9'd18,10'd18};
ram[15427] = {9'd21,10'd21};
ram[15428] = {9'd25,10'd25};
ram[15429] = {9'd28,10'd28};
ram[15430] = {9'd31,10'd31};
ram[15431] = {9'd34,10'd34};
ram[15432] = {9'd37,10'd37};
ram[15433] = {9'd40,10'd40};
ram[15434] = {9'd43,10'd43};
ram[15435] = {9'd47,10'd47};
ram[15436] = {9'd50,10'd50};
ram[15437] = {9'd53,10'd53};
ram[15438] = {9'd56,10'd56};
ram[15439] = {9'd59,10'd59};
ram[15440] = {9'd62,10'd62};
ram[15441] = {9'd65,10'd65};
ram[15442] = {9'd69,10'd69};
ram[15443] = {9'd72,10'd72};
ram[15444] = {9'd75,10'd75};
ram[15445] = {9'd78,10'd78};
ram[15446] = {9'd81,10'd81};
ram[15447] = {9'd84,10'd84};
ram[15448] = {9'd87,10'd87};
ram[15449] = {9'd91,10'd91};
ram[15450] = {9'd94,10'd94};
ram[15451] = {9'd97,10'd97};
ram[15452] = {-9'd100,10'd100};
ram[15453] = {-9'd97,10'd103};
ram[15454] = {-9'd94,10'd106};
ram[15455] = {-9'd91,10'd109};
ram[15456] = {-9'd88,10'd113};
ram[15457] = {-9'd85,10'd116};
ram[15458] = {-9'd81,10'd119};
ram[15459] = {-9'd78,10'd122};
ram[15460] = {-9'd75,10'd125};
ram[15461] = {-9'd72,10'd128};
ram[15462] = {-9'd69,10'd131};
ram[15463] = {-9'd66,10'd135};
ram[15464] = {-9'd63,10'd138};
ram[15465] = {-9'd59,10'd141};
ram[15466] = {-9'd56,10'd144};
ram[15467] = {-9'd53,10'd147};
ram[15468] = {-9'd50,10'd150};
ram[15469] = {-9'd47,10'd153};
ram[15470] = {-9'd44,10'd157};
ram[15471] = {-9'd41,10'd160};
ram[15472] = {-9'd37,10'd163};
ram[15473] = {-9'd34,10'd166};
ram[15474] = {-9'd31,10'd169};
ram[15475] = {-9'd28,10'd172};
ram[15476] = {-9'd25,10'd175};
ram[15477] = {-9'd22,10'd179};
ram[15478] = {-9'd19,10'd182};
ram[15479] = {-9'd15,10'd185};
ram[15480] = {-9'd12,10'd188};
ram[15481] = {-9'd9,10'd191};
ram[15482] = {-9'd6,10'd194};
ram[15483] = {-9'd3,10'd197};
ram[15484] = {9'd0,10'd201};
ram[15485] = {9'd3,10'd204};
ram[15486] = {9'd7,10'd207};
ram[15487] = {9'd10,10'd210};
ram[15488] = {9'd10,10'd210};
ram[15489] = {9'd13,10'd213};
ram[15490] = {9'd16,10'd216};
ram[15491] = {9'd19,10'd219};
ram[15492] = {9'd22,10'd223};
ram[15493] = {9'd25,10'd226};
ram[15494] = {9'd29,10'd229};
ram[15495] = {9'd32,10'd232};
ram[15496] = {9'd35,10'd235};
ram[15497] = {9'd38,10'd238};
ram[15498] = {9'd41,10'd241};
ram[15499] = {9'd44,10'd245};
ram[15500] = {9'd47,10'd248};
ram[15501] = {9'd51,10'd251};
ram[15502] = {9'd54,10'd254};
ram[15503] = {9'd57,10'd257};
ram[15504] = {9'd60,10'd260};
ram[15505] = {9'd63,10'd263};
ram[15506] = {9'd66,10'd267};
ram[15507] = {9'd69,10'd270};
ram[15508] = {9'd73,10'd273};
ram[15509] = {9'd76,10'd276};
ram[15510] = {9'd79,10'd279};
ram[15511] = {9'd82,10'd282};
ram[15512] = {9'd85,10'd285};
ram[15513] = {9'd88,10'd289};
ram[15514] = {9'd91,10'd292};
ram[15515] = {9'd95,10'd295};
ram[15516] = {9'd98,10'd298};
ram[15517] = {-9'd99,10'd301};
ram[15518] = {-9'd96,10'd304};
ram[15519] = {-9'd93,10'd307};
ram[15520] = {-9'd90,10'd311};
ram[15521] = {-9'd87,10'd314};
ram[15522] = {-9'd84,10'd317};
ram[15523] = {-9'd81,10'd320};
ram[15524] = {-9'd77,10'd323};
ram[15525] = {-9'd74,10'd326};
ram[15526] = {-9'd71,10'd329};
ram[15527] = {-9'd68,10'd333};
ram[15528] = {-9'd65,10'd336};
ram[15529] = {-9'd62,10'd339};
ram[15530] = {-9'd59,10'd342};
ram[15531] = {-9'd55,10'd345};
ram[15532] = {-9'd52,10'd348};
ram[15533] = {-9'd49,10'd351};
ram[15534] = {-9'd46,10'd354};
ram[15535] = {-9'd43,10'd358};
ram[15536] = {-9'd40,10'd361};
ram[15537] = {-9'd37,10'd364};
ram[15538] = {-9'd33,10'd367};
ram[15539] = {-9'd30,10'd370};
ram[15540] = {-9'd27,10'd373};
ram[15541] = {-9'd24,10'd376};
ram[15542] = {-9'd21,10'd380};
ram[15543] = {-9'd18,10'd383};
ram[15544] = {-9'd15,10'd386};
ram[15545] = {-9'd11,10'd389};
ram[15546] = {-9'd8,10'd392};
ram[15547] = {-9'd5,10'd395};
ram[15548] = {-9'd2,10'd398};
ram[15549] = {9'd1,-10'd399};
ram[15550] = {9'd4,-10'd396};
ram[15551] = {9'd7,-10'd393};
ram[15552] = {9'd10,-10'd390};
ram[15553] = {9'd14,-10'd387};
ram[15554] = {9'd17,-10'd384};
ram[15555] = {9'd20,-10'd381};
ram[15556] = {9'd23,-10'd377};
ram[15557] = {9'd26,-10'd374};
ram[15558] = {9'd29,-10'd371};
ram[15559] = {9'd32,-10'd368};
ram[15560] = {9'd36,-10'd365};
ram[15561] = {9'd39,-10'd362};
ram[15562] = {9'd42,-10'd359};
ram[15563] = {9'd45,-10'd355};
ram[15564] = {9'd48,-10'd352};
ram[15565] = {9'd51,-10'd349};
ram[15566] = {9'd54,-10'd346};
ram[15567] = {9'd58,-10'd343};
ram[15568] = {9'd61,-10'd340};
ram[15569] = {9'd64,-10'd337};
ram[15570] = {9'd67,-10'd334};
ram[15571] = {9'd70,-10'd330};
ram[15572] = {9'd73,-10'd327};
ram[15573] = {9'd76,-10'd324};
ram[15574] = {9'd80,-10'd321};
ram[15575] = {9'd83,-10'd318};
ram[15576] = {9'd86,-10'd315};
ram[15577] = {9'd89,-10'd312};
ram[15578] = {9'd92,-10'd308};
ram[15579] = {9'd95,-10'd305};
ram[15580] = {9'd98,-10'd302};
ram[15581] = {-9'd99,-10'd299};
ram[15582] = {-9'd96,-10'd296};
ram[15583] = {-9'd92,-10'd293};
ram[15584] = {-9'd89,-10'd290};
ram[15585] = {-9'd86,-10'd286};
ram[15586] = {-9'd83,-10'd283};
ram[15587] = {-9'd80,-10'd280};
ram[15588] = {-9'd77,-10'd277};
ram[15589] = {-9'd74,-10'd274};
ram[15590] = {-9'd70,-10'd271};
ram[15591] = {-9'd67,-10'd268};
ram[15592] = {-9'd64,-10'd264};
ram[15593] = {-9'd61,-10'd261};
ram[15594] = {-9'd58,-10'd258};
ram[15595] = {-9'd55,-10'd255};
ram[15596] = {-9'd52,-10'd252};
ram[15597] = {-9'd48,-10'd249};
ram[15598] = {-9'd45,-10'd246};
ram[15599] = {-9'd42,-10'd242};
ram[15600] = {-9'd39,-10'd239};
ram[15601] = {-9'd36,-10'd236};
ram[15602] = {-9'd33,-10'd233};
ram[15603] = {-9'd30,-10'd230};
ram[15604] = {-9'd26,-10'd227};
ram[15605] = {-9'd23,-10'd224};
ram[15606] = {-9'd20,-10'd220};
ram[15607] = {-9'd17,-10'd217};
ram[15608] = {-9'd14,-10'd214};
ram[15609] = {-9'd11,-10'd211};
ram[15610] = {-9'd8,-10'd208};
ram[15611] = {-9'd4,-10'd205};
ram[15612] = {-9'd1,-10'd202};
ram[15613] = {9'd2,-10'd198};
ram[15614] = {9'd5,-10'd195};
ram[15615] = {9'd8,-10'd192};
ram[15616] = {9'd8,-10'd192};
ram[15617] = {9'd11,-10'd189};
ram[15618] = {9'd14,-10'd186};
ram[15619] = {9'd18,-10'd183};
ram[15620] = {9'd21,-10'd180};
ram[15621] = {9'd24,-10'd176};
ram[15622] = {9'd27,-10'd173};
ram[15623] = {9'd30,-10'd170};
ram[15624] = {9'd33,-10'd167};
ram[15625] = {9'd36,-10'd164};
ram[15626] = {9'd40,-10'd161};
ram[15627] = {9'd43,-10'd158};
ram[15628] = {9'd46,-10'd154};
ram[15629] = {9'd49,-10'd151};
ram[15630] = {9'd52,-10'd148};
ram[15631] = {9'd55,-10'd145};
ram[15632] = {9'd58,-10'd142};
ram[15633] = {9'd62,-10'd139};
ram[15634] = {9'd65,-10'd136};
ram[15635] = {9'd68,-10'd132};
ram[15636] = {9'd71,-10'd129};
ram[15637] = {9'd74,-10'd126};
ram[15638] = {9'd77,-10'd123};
ram[15639] = {9'd80,-10'd120};
ram[15640] = {9'd84,-10'd117};
ram[15641] = {9'd87,-10'd114};
ram[15642] = {9'd90,-10'd110};
ram[15643] = {9'd93,-10'd107};
ram[15644] = {9'd96,-10'd104};
ram[15645] = {9'd99,-10'd101};
ram[15646] = {-9'd98,-10'd98};
ram[15647] = {-9'd95,-10'd95};
ram[15648] = {-9'd92,-10'd92};
ram[15649] = {-9'd88,-10'd88};
ram[15650] = {-9'd85,-10'd85};
ram[15651] = {-9'd82,-10'd82};
ram[15652] = {-9'd79,-10'd79};
ram[15653] = {-9'd76,-10'd76};
ram[15654] = {-9'd73,-10'd73};
ram[15655] = {-9'd70,-10'd70};
ram[15656] = {-9'd66,-10'd66};
ram[15657] = {-9'd63,-10'd63};
ram[15658] = {-9'd60,-10'd60};
ram[15659] = {-9'd57,-10'd57};
ram[15660] = {-9'd54,-10'd54};
ram[15661] = {-9'd51,-10'd51};
ram[15662] = {-9'd48,-10'd48};
ram[15663] = {-9'd44,-10'd44};
ram[15664] = {-9'd41,-10'd41};
ram[15665] = {-9'd38,-10'd38};
ram[15666] = {-9'd35,-10'd35};
ram[15667] = {-9'd32,-10'd32};
ram[15668] = {-9'd29,-10'd29};
ram[15669] = {-9'd26,-10'd26};
ram[15670] = {-9'd22,-10'd22};
ram[15671] = {-9'd19,-10'd19};
ram[15672] = {-9'd16,-10'd16};
ram[15673] = {-9'd13,-10'd13};
ram[15674] = {-9'd10,-10'd10};
ram[15675] = {-9'd7,-10'd7};
ram[15676] = {-9'd4,-10'd4};
ram[15677] = {9'd0,10'd0};
ram[15678] = {9'd3,10'd3};
ram[15679] = {9'd6,10'd6};
ram[15680] = {9'd9,10'd9};
ram[15681] = {9'd12,10'd12};
ram[15682] = {9'd15,10'd15};
ram[15683] = {9'd18,10'd18};
ram[15684] = {9'd21,10'd21};
ram[15685] = {9'd25,10'd25};
ram[15686] = {9'd28,10'd28};
ram[15687] = {9'd31,10'd31};
ram[15688] = {9'd34,10'd34};
ram[15689] = {9'd37,10'd37};
ram[15690] = {9'd40,10'd40};
ram[15691] = {9'd43,10'd43};
ram[15692] = {9'd47,10'd47};
ram[15693] = {9'd50,10'd50};
ram[15694] = {9'd53,10'd53};
ram[15695] = {9'd56,10'd56};
ram[15696] = {9'd59,10'd59};
ram[15697] = {9'd62,10'd62};
ram[15698] = {9'd65,10'd65};
ram[15699] = {9'd69,10'd69};
ram[15700] = {9'd72,10'd72};
ram[15701] = {9'd75,10'd75};
ram[15702] = {9'd78,10'd78};
ram[15703] = {9'd81,10'd81};
ram[15704] = {9'd84,10'd84};
ram[15705] = {9'd87,10'd87};
ram[15706] = {9'd91,10'd91};
ram[15707] = {9'd94,10'd94};
ram[15708] = {9'd97,10'd97};
ram[15709] = {-9'd100,10'd100};
ram[15710] = {-9'd97,10'd103};
ram[15711] = {-9'd94,10'd106};
ram[15712] = {-9'd91,10'd109};
ram[15713] = {-9'd88,10'd113};
ram[15714] = {-9'd85,10'd116};
ram[15715] = {-9'd81,10'd119};
ram[15716] = {-9'd78,10'd122};
ram[15717] = {-9'd75,10'd125};
ram[15718] = {-9'd72,10'd128};
ram[15719] = {-9'd69,10'd131};
ram[15720] = {-9'd66,10'd135};
ram[15721] = {-9'd63,10'd138};
ram[15722] = {-9'd59,10'd141};
ram[15723] = {-9'd56,10'd144};
ram[15724] = {-9'd53,10'd147};
ram[15725] = {-9'd50,10'd150};
ram[15726] = {-9'd47,10'd153};
ram[15727] = {-9'd44,10'd157};
ram[15728] = {-9'd41,10'd160};
ram[15729] = {-9'd37,10'd163};
ram[15730] = {-9'd34,10'd166};
ram[15731] = {-9'd31,10'd169};
ram[15732] = {-9'd28,10'd172};
ram[15733] = {-9'd25,10'd175};
ram[15734] = {-9'd22,10'd179};
ram[15735] = {-9'd19,10'd182};
ram[15736] = {-9'd15,10'd185};
ram[15737] = {-9'd12,10'd188};
ram[15738] = {-9'd9,10'd191};
ram[15739] = {-9'd6,10'd194};
ram[15740] = {-9'd3,10'd197};
ram[15741] = {9'd0,10'd201};
ram[15742] = {9'd3,10'd204};
ram[15743] = {9'd7,10'd207};
ram[15744] = {9'd7,10'd207};
ram[15745] = {9'd10,10'd210};
ram[15746] = {9'd13,10'd213};
ram[15747] = {9'd16,10'd216};
ram[15748] = {9'd19,10'd219};
ram[15749] = {9'd22,10'd223};
ram[15750] = {9'd25,10'd226};
ram[15751] = {9'd29,10'd229};
ram[15752] = {9'd32,10'd232};
ram[15753] = {9'd35,10'd235};
ram[15754] = {9'd38,10'd238};
ram[15755] = {9'd41,10'd241};
ram[15756] = {9'd44,10'd245};
ram[15757] = {9'd47,10'd248};
ram[15758] = {9'd51,10'd251};
ram[15759] = {9'd54,10'd254};
ram[15760] = {9'd57,10'd257};
ram[15761] = {9'd60,10'd260};
ram[15762] = {9'd63,10'd263};
ram[15763] = {9'd66,10'd267};
ram[15764] = {9'd69,10'd270};
ram[15765] = {9'd73,10'd273};
ram[15766] = {9'd76,10'd276};
ram[15767] = {9'd79,10'd279};
ram[15768] = {9'd82,10'd282};
ram[15769] = {9'd85,10'd285};
ram[15770] = {9'd88,10'd289};
ram[15771] = {9'd91,10'd292};
ram[15772] = {9'd95,10'd295};
ram[15773] = {9'd98,10'd298};
ram[15774] = {-9'd99,10'd301};
ram[15775] = {-9'd96,10'd304};
ram[15776] = {-9'd93,10'd307};
ram[15777] = {-9'd90,10'd311};
ram[15778] = {-9'd87,10'd314};
ram[15779] = {-9'd84,10'd317};
ram[15780] = {-9'd81,10'd320};
ram[15781] = {-9'd77,10'd323};
ram[15782] = {-9'd74,10'd326};
ram[15783] = {-9'd71,10'd329};
ram[15784] = {-9'd68,10'd333};
ram[15785] = {-9'd65,10'd336};
ram[15786] = {-9'd62,10'd339};
ram[15787] = {-9'd59,10'd342};
ram[15788] = {-9'd55,10'd345};
ram[15789] = {-9'd52,10'd348};
ram[15790] = {-9'd49,10'd351};
ram[15791] = {-9'd46,10'd354};
ram[15792] = {-9'd43,10'd358};
ram[15793] = {-9'd40,10'd361};
ram[15794] = {-9'd37,10'd364};
ram[15795] = {-9'd33,10'd367};
ram[15796] = {-9'd30,10'd370};
ram[15797] = {-9'd27,10'd373};
ram[15798] = {-9'd24,10'd376};
ram[15799] = {-9'd21,10'd380};
ram[15800] = {-9'd18,10'd383};
ram[15801] = {-9'd15,10'd386};
ram[15802] = {-9'd11,10'd389};
ram[15803] = {-9'd8,10'd392};
ram[15804] = {-9'd5,10'd395};
ram[15805] = {-9'd2,10'd398};
ram[15806] = {9'd1,-10'd399};
ram[15807] = {9'd4,-10'd396};
ram[15808] = {9'd7,-10'd393};
ram[15809] = {9'd10,-10'd390};
ram[15810] = {9'd14,-10'd387};
ram[15811] = {9'd17,-10'd384};
ram[15812] = {9'd20,-10'd381};
ram[15813] = {9'd23,-10'd377};
ram[15814] = {9'd26,-10'd374};
ram[15815] = {9'd29,-10'd371};
ram[15816] = {9'd32,-10'd368};
ram[15817] = {9'd36,-10'd365};
ram[15818] = {9'd39,-10'd362};
ram[15819] = {9'd42,-10'd359};
ram[15820] = {9'd45,-10'd355};
ram[15821] = {9'd48,-10'd352};
ram[15822] = {9'd51,-10'd349};
ram[15823] = {9'd54,-10'd346};
ram[15824] = {9'd58,-10'd343};
ram[15825] = {9'd61,-10'd340};
ram[15826] = {9'd64,-10'd337};
ram[15827] = {9'd67,-10'd334};
ram[15828] = {9'd70,-10'd330};
ram[15829] = {9'd73,-10'd327};
ram[15830] = {9'd76,-10'd324};
ram[15831] = {9'd80,-10'd321};
ram[15832] = {9'd83,-10'd318};
ram[15833] = {9'd86,-10'd315};
ram[15834] = {9'd89,-10'd312};
ram[15835] = {9'd92,-10'd308};
ram[15836] = {9'd95,-10'd305};
ram[15837] = {9'd98,-10'd302};
ram[15838] = {-9'd99,-10'd299};
ram[15839] = {-9'd96,-10'd296};
ram[15840] = {-9'd92,-10'd293};
ram[15841] = {-9'd89,-10'd290};
ram[15842] = {-9'd86,-10'd286};
ram[15843] = {-9'd83,-10'd283};
ram[15844] = {-9'd80,-10'd280};
ram[15845] = {-9'd77,-10'd277};
ram[15846] = {-9'd74,-10'd274};
ram[15847] = {-9'd70,-10'd271};
ram[15848] = {-9'd67,-10'd268};
ram[15849] = {-9'd64,-10'd264};
ram[15850] = {-9'd61,-10'd261};
ram[15851] = {-9'd58,-10'd258};
ram[15852] = {-9'd55,-10'd255};
ram[15853] = {-9'd52,-10'd252};
ram[15854] = {-9'd48,-10'd249};
ram[15855] = {-9'd45,-10'd246};
ram[15856] = {-9'd42,-10'd242};
ram[15857] = {-9'd39,-10'd239};
ram[15858] = {-9'd36,-10'd236};
ram[15859] = {-9'd33,-10'd233};
ram[15860] = {-9'd30,-10'd230};
ram[15861] = {-9'd26,-10'd227};
ram[15862] = {-9'd23,-10'd224};
ram[15863] = {-9'd20,-10'd220};
ram[15864] = {-9'd17,-10'd217};
ram[15865] = {-9'd14,-10'd214};
ram[15866] = {-9'd11,-10'd211};
ram[15867] = {-9'd8,-10'd208};
ram[15868] = {-9'd4,-10'd205};
ram[15869] = {-9'd1,-10'd202};
ram[15870] = {9'd2,-10'd198};
ram[15871] = {9'd5,-10'd195};
ram[15872] = {9'd5,-10'd195};
ram[15873] = {9'd8,-10'd192};
ram[15874] = {9'd11,-10'd189};
ram[15875] = {9'd14,-10'd186};
ram[15876] = {9'd18,-10'd183};
ram[15877] = {9'd21,-10'd180};
ram[15878] = {9'd24,-10'd176};
ram[15879] = {9'd27,-10'd173};
ram[15880] = {9'd30,-10'd170};
ram[15881] = {9'd33,-10'd167};
ram[15882] = {9'd36,-10'd164};
ram[15883] = {9'd40,-10'd161};
ram[15884] = {9'd43,-10'd158};
ram[15885] = {9'd46,-10'd154};
ram[15886] = {9'd49,-10'd151};
ram[15887] = {9'd52,-10'd148};
ram[15888] = {9'd55,-10'd145};
ram[15889] = {9'd58,-10'd142};
ram[15890] = {9'd62,-10'd139};
ram[15891] = {9'd65,-10'd136};
ram[15892] = {9'd68,-10'd132};
ram[15893] = {9'd71,-10'd129};
ram[15894] = {9'd74,-10'd126};
ram[15895] = {9'd77,-10'd123};
ram[15896] = {9'd80,-10'd120};
ram[15897] = {9'd84,-10'd117};
ram[15898] = {9'd87,-10'd114};
ram[15899] = {9'd90,-10'd110};
ram[15900] = {9'd93,-10'd107};
ram[15901] = {9'd96,-10'd104};
ram[15902] = {9'd99,-10'd101};
ram[15903] = {-9'd98,-10'd98};
ram[15904] = {-9'd95,-10'd95};
ram[15905] = {-9'd92,-10'd92};
ram[15906] = {-9'd88,-10'd88};
ram[15907] = {-9'd85,-10'd85};
ram[15908] = {-9'd82,-10'd82};
ram[15909] = {-9'd79,-10'd79};
ram[15910] = {-9'd76,-10'd76};
ram[15911] = {-9'd73,-10'd73};
ram[15912] = {-9'd70,-10'd70};
ram[15913] = {-9'd66,-10'd66};
ram[15914] = {-9'd63,-10'd63};
ram[15915] = {-9'd60,-10'd60};
ram[15916] = {-9'd57,-10'd57};
ram[15917] = {-9'd54,-10'd54};
ram[15918] = {-9'd51,-10'd51};
ram[15919] = {-9'd48,-10'd48};
ram[15920] = {-9'd44,-10'd44};
ram[15921] = {-9'd41,-10'd41};
ram[15922] = {-9'd38,-10'd38};
ram[15923] = {-9'd35,-10'd35};
ram[15924] = {-9'd32,-10'd32};
ram[15925] = {-9'd29,-10'd29};
ram[15926] = {-9'd26,-10'd26};
ram[15927] = {-9'd22,-10'd22};
ram[15928] = {-9'd19,-10'd19};
ram[15929] = {-9'd16,-10'd16};
ram[15930] = {-9'd13,-10'd13};
ram[15931] = {-9'd10,-10'd10};
ram[15932] = {-9'd7,-10'd7};
ram[15933] = {-9'd4,-10'd4};
ram[15934] = {9'd0,10'd0};
ram[15935] = {9'd3,10'd3};
ram[15936] = {9'd6,10'd6};
ram[15937] = {9'd9,10'd9};
ram[15938] = {9'd12,10'd12};
ram[15939] = {9'd15,10'd15};
ram[15940] = {9'd18,10'd18};
ram[15941] = {9'd21,10'd21};
ram[15942] = {9'd25,10'd25};
ram[15943] = {9'd28,10'd28};
ram[15944] = {9'd31,10'd31};
ram[15945] = {9'd34,10'd34};
ram[15946] = {9'd37,10'd37};
ram[15947] = {9'd40,10'd40};
ram[15948] = {9'd43,10'd43};
ram[15949] = {9'd47,10'd47};
ram[15950] = {9'd50,10'd50};
ram[15951] = {9'd53,10'd53};
ram[15952] = {9'd56,10'd56};
ram[15953] = {9'd59,10'd59};
ram[15954] = {9'd62,10'd62};
ram[15955] = {9'd65,10'd65};
ram[15956] = {9'd69,10'd69};
ram[15957] = {9'd72,10'd72};
ram[15958] = {9'd75,10'd75};
ram[15959] = {9'd78,10'd78};
ram[15960] = {9'd81,10'd81};
ram[15961] = {9'd84,10'd84};
ram[15962] = {9'd87,10'd87};
ram[15963] = {9'd91,10'd91};
ram[15964] = {9'd94,10'd94};
ram[15965] = {9'd97,10'd97};
ram[15966] = {-9'd100,10'd100};
ram[15967] = {-9'd97,10'd103};
ram[15968] = {-9'd94,10'd106};
ram[15969] = {-9'd91,10'd109};
ram[15970] = {-9'd88,10'd113};
ram[15971] = {-9'd85,10'd116};
ram[15972] = {-9'd81,10'd119};
ram[15973] = {-9'd78,10'd122};
ram[15974] = {-9'd75,10'd125};
ram[15975] = {-9'd72,10'd128};
ram[15976] = {-9'd69,10'd131};
ram[15977] = {-9'd66,10'd135};
ram[15978] = {-9'd63,10'd138};
ram[15979] = {-9'd59,10'd141};
ram[15980] = {-9'd56,10'd144};
ram[15981] = {-9'd53,10'd147};
ram[15982] = {-9'd50,10'd150};
ram[15983] = {-9'd47,10'd153};
ram[15984] = {-9'd44,10'd157};
ram[15985] = {-9'd41,10'd160};
ram[15986] = {-9'd37,10'd163};
ram[15987] = {-9'd34,10'd166};
ram[15988] = {-9'd31,10'd169};
ram[15989] = {-9'd28,10'd172};
ram[15990] = {-9'd25,10'd175};
ram[15991] = {-9'd22,10'd179};
ram[15992] = {-9'd19,10'd182};
ram[15993] = {-9'd15,10'd185};
ram[15994] = {-9'd12,10'd188};
ram[15995] = {-9'd9,10'd191};
ram[15996] = {-9'd6,10'd194};
ram[15997] = {-9'd3,10'd197};
ram[15998] = {9'd0,10'd201};
ram[15999] = {9'd3,10'd204};
ram[16000] = {9'd3,10'd204};
ram[16001] = {9'd7,10'd207};
ram[16002] = {9'd10,10'd210};
ram[16003] = {9'd13,10'd213};
ram[16004] = {9'd16,10'd216};
ram[16005] = {9'd19,10'd219};
ram[16006] = {9'd22,10'd223};
ram[16007] = {9'd25,10'd226};
ram[16008] = {9'd29,10'd229};
ram[16009] = {9'd32,10'd232};
ram[16010] = {9'd35,10'd235};
ram[16011] = {9'd38,10'd238};
ram[16012] = {9'd41,10'd241};
ram[16013] = {9'd44,10'd245};
ram[16014] = {9'd47,10'd248};
ram[16015] = {9'd51,10'd251};
ram[16016] = {9'd54,10'd254};
ram[16017] = {9'd57,10'd257};
ram[16018] = {9'd60,10'd260};
ram[16019] = {9'd63,10'd263};
ram[16020] = {9'd66,10'd267};
ram[16021] = {9'd69,10'd270};
ram[16022] = {9'd73,10'd273};
ram[16023] = {9'd76,10'd276};
ram[16024] = {9'd79,10'd279};
ram[16025] = {9'd82,10'd282};
ram[16026] = {9'd85,10'd285};
ram[16027] = {9'd88,10'd289};
ram[16028] = {9'd91,10'd292};
ram[16029] = {9'd95,10'd295};
ram[16030] = {9'd98,10'd298};
ram[16031] = {-9'd99,10'd301};
ram[16032] = {-9'd96,10'd304};
ram[16033] = {-9'd93,10'd307};
ram[16034] = {-9'd90,10'd311};
ram[16035] = {-9'd87,10'd314};
ram[16036] = {-9'd84,10'd317};
ram[16037] = {-9'd81,10'd320};
ram[16038] = {-9'd77,10'd323};
ram[16039] = {-9'd74,10'd326};
ram[16040] = {-9'd71,10'd329};
ram[16041] = {-9'd68,10'd333};
ram[16042] = {-9'd65,10'd336};
ram[16043] = {-9'd62,10'd339};
ram[16044] = {-9'd59,10'd342};
ram[16045] = {-9'd55,10'd345};
ram[16046] = {-9'd52,10'd348};
ram[16047] = {-9'd49,10'd351};
ram[16048] = {-9'd46,10'd354};
ram[16049] = {-9'd43,10'd358};
ram[16050] = {-9'd40,10'd361};
ram[16051] = {-9'd37,10'd364};
ram[16052] = {-9'd33,10'd367};
ram[16053] = {-9'd30,10'd370};
ram[16054] = {-9'd27,10'd373};
ram[16055] = {-9'd24,10'd376};
ram[16056] = {-9'd21,10'd380};
ram[16057] = {-9'd18,10'd383};
ram[16058] = {-9'd15,10'd386};
ram[16059] = {-9'd11,10'd389};
ram[16060] = {-9'd8,10'd392};
ram[16061] = {-9'd5,10'd395};
ram[16062] = {-9'd2,10'd398};
ram[16063] = {9'd1,-10'd399};
ram[16064] = {9'd4,-10'd396};
ram[16065] = {9'd7,-10'd393};
ram[16066] = {9'd10,-10'd390};
ram[16067] = {9'd14,-10'd387};
ram[16068] = {9'd17,-10'd384};
ram[16069] = {9'd20,-10'd381};
ram[16070] = {9'd23,-10'd377};
ram[16071] = {9'd26,-10'd374};
ram[16072] = {9'd29,-10'd371};
ram[16073] = {9'd32,-10'd368};
ram[16074] = {9'd36,-10'd365};
ram[16075] = {9'd39,-10'd362};
ram[16076] = {9'd42,-10'd359};
ram[16077] = {9'd45,-10'd355};
ram[16078] = {9'd48,-10'd352};
ram[16079] = {9'd51,-10'd349};
ram[16080] = {9'd54,-10'd346};
ram[16081] = {9'd58,-10'd343};
ram[16082] = {9'd61,-10'd340};
ram[16083] = {9'd64,-10'd337};
ram[16084] = {9'd67,-10'd334};
ram[16085] = {9'd70,-10'd330};
ram[16086] = {9'd73,-10'd327};
ram[16087] = {9'd76,-10'd324};
ram[16088] = {9'd80,-10'd321};
ram[16089] = {9'd83,-10'd318};
ram[16090] = {9'd86,-10'd315};
ram[16091] = {9'd89,-10'd312};
ram[16092] = {9'd92,-10'd308};
ram[16093] = {9'd95,-10'd305};
ram[16094] = {9'd98,-10'd302};
ram[16095] = {-9'd99,-10'd299};
ram[16096] = {-9'd96,-10'd296};
ram[16097] = {-9'd92,-10'd293};
ram[16098] = {-9'd89,-10'd290};
ram[16099] = {-9'd86,-10'd286};
ram[16100] = {-9'd83,-10'd283};
ram[16101] = {-9'd80,-10'd280};
ram[16102] = {-9'd77,-10'd277};
ram[16103] = {-9'd74,-10'd274};
ram[16104] = {-9'd70,-10'd271};
ram[16105] = {-9'd67,-10'd268};
ram[16106] = {-9'd64,-10'd264};
ram[16107] = {-9'd61,-10'd261};
ram[16108] = {-9'd58,-10'd258};
ram[16109] = {-9'd55,-10'd255};
ram[16110] = {-9'd52,-10'd252};
ram[16111] = {-9'd48,-10'd249};
ram[16112] = {-9'd45,-10'd246};
ram[16113] = {-9'd42,-10'd242};
ram[16114] = {-9'd39,-10'd239};
ram[16115] = {-9'd36,-10'd236};
ram[16116] = {-9'd33,-10'd233};
ram[16117] = {-9'd30,-10'd230};
ram[16118] = {-9'd26,-10'd227};
ram[16119] = {-9'd23,-10'd224};
ram[16120] = {-9'd20,-10'd220};
ram[16121] = {-9'd17,-10'd217};
ram[16122] = {-9'd14,-10'd214};
ram[16123] = {-9'd11,-10'd211};
ram[16124] = {-9'd8,-10'd208};
ram[16125] = {-9'd4,-10'd205};
ram[16126] = {-9'd1,-10'd202};
ram[16127] = {9'd2,-10'd198};
ram[16128] = {9'd2,-10'd198};
ram[16129] = {9'd5,-10'd195};
ram[16130] = {9'd8,-10'd192};
ram[16131] = {9'd11,-10'd189};
ram[16132] = {9'd14,-10'd186};
ram[16133] = {9'd18,-10'd183};
ram[16134] = {9'd21,-10'd180};
ram[16135] = {9'd24,-10'd176};
ram[16136] = {9'd27,-10'd173};
ram[16137] = {9'd30,-10'd170};
ram[16138] = {9'd33,-10'd167};
ram[16139] = {9'd36,-10'd164};
ram[16140] = {9'd40,-10'd161};
ram[16141] = {9'd43,-10'd158};
ram[16142] = {9'd46,-10'd154};
ram[16143] = {9'd49,-10'd151};
ram[16144] = {9'd52,-10'd148};
ram[16145] = {9'd55,-10'd145};
ram[16146] = {9'd58,-10'd142};
ram[16147] = {9'd62,-10'd139};
ram[16148] = {9'd65,-10'd136};
ram[16149] = {9'd68,-10'd132};
ram[16150] = {9'd71,-10'd129};
ram[16151] = {9'd74,-10'd126};
ram[16152] = {9'd77,-10'd123};
ram[16153] = {9'd80,-10'd120};
ram[16154] = {9'd84,-10'd117};
ram[16155] = {9'd87,-10'd114};
ram[16156] = {9'd90,-10'd110};
ram[16157] = {9'd93,-10'd107};
ram[16158] = {9'd96,-10'd104};
ram[16159] = {9'd99,-10'd101};
ram[16160] = {-9'd98,-10'd98};
ram[16161] = {-9'd95,-10'd95};
ram[16162] = {-9'd92,-10'd92};
ram[16163] = {-9'd88,-10'd88};
ram[16164] = {-9'd85,-10'd85};
ram[16165] = {-9'd82,-10'd82};
ram[16166] = {-9'd79,-10'd79};
ram[16167] = {-9'd76,-10'd76};
ram[16168] = {-9'd73,-10'd73};
ram[16169] = {-9'd70,-10'd70};
ram[16170] = {-9'd66,-10'd66};
ram[16171] = {-9'd63,-10'd63};
ram[16172] = {-9'd60,-10'd60};
ram[16173] = {-9'd57,-10'd57};
ram[16174] = {-9'd54,-10'd54};
ram[16175] = {-9'd51,-10'd51};
ram[16176] = {-9'd48,-10'd48};
ram[16177] = {-9'd44,-10'd44};
ram[16178] = {-9'd41,-10'd41};
ram[16179] = {-9'd38,-10'd38};
ram[16180] = {-9'd35,-10'd35};
ram[16181] = {-9'd32,-10'd32};
ram[16182] = {-9'd29,-10'd29};
ram[16183] = {-9'd26,-10'd26};
ram[16184] = {-9'd22,-10'd22};
ram[16185] = {-9'd19,-10'd19};
ram[16186] = {-9'd16,-10'd16};
ram[16187] = {-9'd13,-10'd13};
ram[16188] = {-9'd10,-10'd10};
ram[16189] = {-9'd7,-10'd7};
ram[16190] = {-9'd4,-10'd4};
ram[16191] = {9'd0,10'd0};
ram[16192] = {9'd3,10'd3};
ram[16193] = {9'd6,10'd6};
ram[16194] = {9'd9,10'd9};
ram[16195] = {9'd12,10'd12};
ram[16196] = {9'd15,10'd15};
ram[16197] = {9'd18,10'd18};
ram[16198] = {9'd21,10'd21};
ram[16199] = {9'd25,10'd25};
ram[16200] = {9'd28,10'd28};
ram[16201] = {9'd31,10'd31};
ram[16202] = {9'd34,10'd34};
ram[16203] = {9'd37,10'd37};
ram[16204] = {9'd40,10'd40};
ram[16205] = {9'd43,10'd43};
ram[16206] = {9'd47,10'd47};
ram[16207] = {9'd50,10'd50};
ram[16208] = {9'd53,10'd53};
ram[16209] = {9'd56,10'd56};
ram[16210] = {9'd59,10'd59};
ram[16211] = {9'd62,10'd62};
ram[16212] = {9'd65,10'd65};
ram[16213] = {9'd69,10'd69};
ram[16214] = {9'd72,10'd72};
ram[16215] = {9'd75,10'd75};
ram[16216] = {9'd78,10'd78};
ram[16217] = {9'd81,10'd81};
ram[16218] = {9'd84,10'd84};
ram[16219] = {9'd87,10'd87};
ram[16220] = {9'd91,10'd91};
ram[16221] = {9'd94,10'd94};
ram[16222] = {9'd97,10'd97};
ram[16223] = {-9'd100,10'd100};
ram[16224] = {-9'd97,10'd103};
ram[16225] = {-9'd94,10'd106};
ram[16226] = {-9'd91,10'd109};
ram[16227] = {-9'd88,10'd113};
ram[16228] = {-9'd85,10'd116};
ram[16229] = {-9'd81,10'd119};
ram[16230] = {-9'd78,10'd122};
ram[16231] = {-9'd75,10'd125};
ram[16232] = {-9'd72,10'd128};
ram[16233] = {-9'd69,10'd131};
ram[16234] = {-9'd66,10'd135};
ram[16235] = {-9'd63,10'd138};
ram[16236] = {-9'd59,10'd141};
ram[16237] = {-9'd56,10'd144};
ram[16238] = {-9'd53,10'd147};
ram[16239] = {-9'd50,10'd150};
ram[16240] = {-9'd47,10'd153};
ram[16241] = {-9'd44,10'd157};
ram[16242] = {-9'd41,10'd160};
ram[16243] = {-9'd37,10'd163};
ram[16244] = {-9'd34,10'd166};
ram[16245] = {-9'd31,10'd169};
ram[16246] = {-9'd28,10'd172};
ram[16247] = {-9'd25,10'd175};
ram[16248] = {-9'd22,10'd179};
ram[16249] = {-9'd19,10'd182};
ram[16250] = {-9'd15,10'd185};
ram[16251] = {-9'd12,10'd188};
ram[16252] = {-9'd9,10'd191};
ram[16253] = {-9'd6,10'd194};
ram[16254] = {-9'd3,10'd197};
ram[16255] = {9'd0,10'd201};
ram[16256] = {9'd0,10'd201};
ram[16257] = {9'd3,10'd204};
ram[16258] = {9'd7,10'd207};
ram[16259] = {9'd10,10'd210};
ram[16260] = {9'd13,10'd213};
ram[16261] = {9'd16,10'd216};
ram[16262] = {9'd19,10'd219};
ram[16263] = {9'd22,10'd223};
ram[16264] = {9'd25,10'd226};
ram[16265] = {9'd29,10'd229};
ram[16266] = {9'd32,10'd232};
ram[16267] = {9'd35,10'd235};
ram[16268] = {9'd38,10'd238};
ram[16269] = {9'd41,10'd241};
ram[16270] = {9'd44,10'd245};
ram[16271] = {9'd47,10'd248};
ram[16272] = {9'd51,10'd251};
ram[16273] = {9'd54,10'd254};
ram[16274] = {9'd57,10'd257};
ram[16275] = {9'd60,10'd260};
ram[16276] = {9'd63,10'd263};
ram[16277] = {9'd66,10'd267};
ram[16278] = {9'd69,10'd270};
ram[16279] = {9'd73,10'd273};
ram[16280] = {9'd76,10'd276};
ram[16281] = {9'd79,10'd279};
ram[16282] = {9'd82,10'd282};
ram[16283] = {9'd85,10'd285};
ram[16284] = {9'd88,10'd289};
ram[16285] = {9'd91,10'd292};
ram[16286] = {9'd95,10'd295};
ram[16287] = {9'd98,10'd298};
ram[16288] = {-9'd99,10'd301};
ram[16289] = {-9'd96,10'd304};
ram[16290] = {-9'd93,10'd307};
ram[16291] = {-9'd90,10'd311};
ram[16292] = {-9'd87,10'd314};
ram[16293] = {-9'd84,10'd317};
ram[16294] = {-9'd81,10'd320};
ram[16295] = {-9'd77,10'd323};
ram[16296] = {-9'd74,10'd326};
ram[16297] = {-9'd71,10'd329};
ram[16298] = {-9'd68,10'd333};
ram[16299] = {-9'd65,10'd336};
ram[16300] = {-9'd62,10'd339};
ram[16301] = {-9'd59,10'd342};
ram[16302] = {-9'd55,10'd345};
ram[16303] = {-9'd52,10'd348};
ram[16304] = {-9'd49,10'd351};
ram[16305] = {-9'd46,10'd354};
ram[16306] = {-9'd43,10'd358};
ram[16307] = {-9'd40,10'd361};
ram[16308] = {-9'd37,10'd364};
ram[16309] = {-9'd33,10'd367};
ram[16310] = {-9'd30,10'd370};
ram[16311] = {-9'd27,10'd373};
ram[16312] = {-9'd24,10'd376};
ram[16313] = {-9'd21,10'd380};
ram[16314] = {-9'd18,10'd383};
ram[16315] = {-9'd15,10'd386};
ram[16316] = {-9'd11,10'd389};
ram[16317] = {-9'd8,10'd392};
ram[16318] = {-9'd5,10'd395};
ram[16319] = {-9'd2,10'd398};
ram[16320] = {9'd1,-10'd399};
ram[16321] = {9'd4,-10'd396};
ram[16322] = {9'd7,-10'd393};
ram[16323] = {9'd10,-10'd390};
ram[16324] = {9'd14,-10'd387};
ram[16325] = {9'd17,-10'd384};
ram[16326] = {9'd20,-10'd381};
ram[16327] = {9'd23,-10'd377};
ram[16328] = {9'd26,-10'd374};
ram[16329] = {9'd29,-10'd371};
ram[16330] = {9'd32,-10'd368};
ram[16331] = {9'd36,-10'd365};
ram[16332] = {9'd39,-10'd362};
ram[16333] = {9'd42,-10'd359};
ram[16334] = {9'd45,-10'd355};
ram[16335] = {9'd48,-10'd352};
ram[16336] = {9'd51,-10'd349};
ram[16337] = {9'd54,-10'd346};
ram[16338] = {9'd58,-10'd343};
ram[16339] = {9'd61,-10'd340};
ram[16340] = {9'd64,-10'd337};
ram[16341] = {9'd67,-10'd334};
ram[16342] = {9'd70,-10'd330};
ram[16343] = {9'd73,-10'd327};
ram[16344] = {9'd76,-10'd324};
ram[16345] = {9'd80,-10'd321};
ram[16346] = {9'd83,-10'd318};
ram[16347] = {9'd86,-10'd315};
ram[16348] = {9'd89,-10'd312};
ram[16349] = {9'd92,-10'd308};
ram[16350] = {9'd95,-10'd305};
ram[16351] = {9'd98,-10'd302};
ram[16352] = {-9'd99,-10'd299};
ram[16353] = {-9'd96,-10'd296};
ram[16354] = {-9'd92,-10'd293};
ram[16355] = {-9'd89,-10'd290};
ram[16356] = {-9'd86,-10'd286};
ram[16357] = {-9'd83,-10'd283};
ram[16358] = {-9'd80,-10'd280};
ram[16359] = {-9'd77,-10'd277};
ram[16360] = {-9'd74,-10'd274};
ram[16361] = {-9'd70,-10'd271};
ram[16362] = {-9'd67,-10'd268};
ram[16363] = {-9'd64,-10'd264};
ram[16364] = {-9'd61,-10'd261};
ram[16365] = {-9'd58,-10'd258};
ram[16366] = {-9'd55,-10'd255};
ram[16367] = {-9'd52,-10'd252};
ram[16368] = {-9'd48,-10'd249};
ram[16369] = {-9'd45,-10'd246};
ram[16370] = {-9'd42,-10'd242};
ram[16371] = {-9'd39,-10'd239};
ram[16372] = {-9'd36,-10'd236};
ram[16373] = {-9'd33,-10'd233};
ram[16374] = {-9'd30,-10'd230};
ram[16375] = {-9'd26,-10'd227};
ram[16376] = {-9'd23,-10'd224};
ram[16377] = {-9'd20,-10'd220};
ram[16378] = {-9'd17,-10'd217};
ram[16379] = {-9'd14,-10'd214};
ram[16380] = {-9'd11,-10'd211};
ram[16381] = {-9'd8,-10'd208};
ram[16382] = {-9'd4,-10'd205};
ram[16383] = {-9'd1,-10'd202};
ram[16384] = {-9'd1,-10'd202};
ram[16385] = {9'd2,-10'd198};
ram[16386] = {9'd5,-10'd195};
ram[16387] = {9'd8,-10'd192};
ram[16388] = {9'd11,-10'd189};
ram[16389] = {9'd14,-10'd186};
ram[16390] = {9'd18,-10'd183};
ram[16391] = {9'd21,-10'd180};
ram[16392] = {9'd24,-10'd176};
ram[16393] = {9'd27,-10'd173};
ram[16394] = {9'd30,-10'd170};
ram[16395] = {9'd33,-10'd167};
ram[16396] = {9'd36,-10'd164};
ram[16397] = {9'd40,-10'd161};
ram[16398] = {9'd43,-10'd158};
ram[16399] = {9'd46,-10'd154};
ram[16400] = {9'd49,-10'd151};
ram[16401] = {9'd52,-10'd148};
ram[16402] = {9'd55,-10'd145};
ram[16403] = {9'd58,-10'd142};
ram[16404] = {9'd62,-10'd139};
ram[16405] = {9'd65,-10'd136};
ram[16406] = {9'd68,-10'd132};
ram[16407] = {9'd71,-10'd129};
ram[16408] = {9'd74,-10'd126};
ram[16409] = {9'd77,-10'd123};
ram[16410] = {9'd80,-10'd120};
ram[16411] = {9'd84,-10'd117};
ram[16412] = {9'd87,-10'd114};
ram[16413] = {9'd90,-10'd110};
ram[16414] = {9'd93,-10'd107};
ram[16415] = {9'd96,-10'd104};
ram[16416] = {9'd99,-10'd101};
ram[16417] = {-9'd98,-10'd98};
ram[16418] = {-9'd95,-10'd95};
ram[16419] = {-9'd92,-10'd92};
ram[16420] = {-9'd88,-10'd88};
ram[16421] = {-9'd85,-10'd85};
ram[16422] = {-9'd82,-10'd82};
ram[16423] = {-9'd79,-10'd79};
ram[16424] = {-9'd76,-10'd76};
ram[16425] = {-9'd73,-10'd73};
ram[16426] = {-9'd70,-10'd70};
ram[16427] = {-9'd66,-10'd66};
ram[16428] = {-9'd63,-10'd63};
ram[16429] = {-9'd60,-10'd60};
ram[16430] = {-9'd57,-10'd57};
ram[16431] = {-9'd54,-10'd54};
ram[16432] = {-9'd51,-10'd51};
ram[16433] = {-9'd48,-10'd48};
ram[16434] = {-9'd44,-10'd44};
ram[16435] = {-9'd41,-10'd41};
ram[16436] = {-9'd38,-10'd38};
ram[16437] = {-9'd35,-10'd35};
ram[16438] = {-9'd32,-10'd32};
ram[16439] = {-9'd29,-10'd29};
ram[16440] = {-9'd26,-10'd26};
ram[16441] = {-9'd22,-10'd22};
ram[16442] = {-9'd19,-10'd19};
ram[16443] = {-9'd16,-10'd16};
ram[16444] = {-9'd13,-10'd13};
ram[16445] = {-9'd10,-10'd10};
ram[16446] = {-9'd7,-10'd7};
ram[16447] = {-9'd4,-10'd4};
ram[16448] = {9'd0,10'd0};
ram[16449] = {9'd3,10'd3};
ram[16450] = {9'd6,10'd6};
ram[16451] = {9'd9,10'd9};
ram[16452] = {9'd12,10'd12};
ram[16453] = {9'd15,10'd15};
ram[16454] = {9'd18,10'd18};
ram[16455] = {9'd21,10'd21};
ram[16456] = {9'd25,10'd25};
ram[16457] = {9'd28,10'd28};
ram[16458] = {9'd31,10'd31};
ram[16459] = {9'd34,10'd34};
ram[16460] = {9'd37,10'd37};
ram[16461] = {9'd40,10'd40};
ram[16462] = {9'd43,10'd43};
ram[16463] = {9'd47,10'd47};
ram[16464] = {9'd50,10'd50};
ram[16465] = {9'd53,10'd53};
ram[16466] = {9'd56,10'd56};
ram[16467] = {9'd59,10'd59};
ram[16468] = {9'd62,10'd62};
ram[16469] = {9'd65,10'd65};
ram[16470] = {9'd69,10'd69};
ram[16471] = {9'd72,10'd72};
ram[16472] = {9'd75,10'd75};
ram[16473] = {9'd78,10'd78};
ram[16474] = {9'd81,10'd81};
ram[16475] = {9'd84,10'd84};
ram[16476] = {9'd87,10'd87};
ram[16477] = {9'd91,10'd91};
ram[16478] = {9'd94,10'd94};
ram[16479] = {9'd97,10'd97};
ram[16480] = {-9'd100,10'd100};
ram[16481] = {-9'd97,10'd103};
ram[16482] = {-9'd94,10'd106};
ram[16483] = {-9'd91,10'd109};
ram[16484] = {-9'd88,10'd113};
ram[16485] = {-9'd85,10'd116};
ram[16486] = {-9'd81,10'd119};
ram[16487] = {-9'd78,10'd122};
ram[16488] = {-9'd75,10'd125};
ram[16489] = {-9'd72,10'd128};
ram[16490] = {-9'd69,10'd131};
ram[16491] = {-9'd66,10'd135};
ram[16492] = {-9'd63,10'd138};
ram[16493] = {-9'd59,10'd141};
ram[16494] = {-9'd56,10'd144};
ram[16495] = {-9'd53,10'd147};
ram[16496] = {-9'd50,10'd150};
ram[16497] = {-9'd47,10'd153};
ram[16498] = {-9'd44,10'd157};
ram[16499] = {-9'd41,10'd160};
ram[16500] = {-9'd37,10'd163};
ram[16501] = {-9'd34,10'd166};
ram[16502] = {-9'd31,10'd169};
ram[16503] = {-9'd28,10'd172};
ram[16504] = {-9'd25,10'd175};
ram[16505] = {-9'd22,10'd179};
ram[16506] = {-9'd19,10'd182};
ram[16507] = {-9'd15,10'd185};
ram[16508] = {-9'd12,10'd188};
ram[16509] = {-9'd9,10'd191};
ram[16510] = {-9'd6,10'd194};
ram[16511] = {-9'd3,10'd197};
ram[16512] = {-9'd3,10'd197};
ram[16513] = {9'd0,10'd201};
ram[16514] = {9'd3,10'd204};
ram[16515] = {9'd7,10'd207};
ram[16516] = {9'd10,10'd210};
ram[16517] = {9'd13,10'd213};
ram[16518] = {9'd16,10'd216};
ram[16519] = {9'd19,10'd219};
ram[16520] = {9'd22,10'd223};
ram[16521] = {9'd25,10'd226};
ram[16522] = {9'd29,10'd229};
ram[16523] = {9'd32,10'd232};
ram[16524] = {9'd35,10'd235};
ram[16525] = {9'd38,10'd238};
ram[16526] = {9'd41,10'd241};
ram[16527] = {9'd44,10'd245};
ram[16528] = {9'd47,10'd248};
ram[16529] = {9'd51,10'd251};
ram[16530] = {9'd54,10'd254};
ram[16531] = {9'd57,10'd257};
ram[16532] = {9'd60,10'd260};
ram[16533] = {9'd63,10'd263};
ram[16534] = {9'd66,10'd267};
ram[16535] = {9'd69,10'd270};
ram[16536] = {9'd73,10'd273};
ram[16537] = {9'd76,10'd276};
ram[16538] = {9'd79,10'd279};
ram[16539] = {9'd82,10'd282};
ram[16540] = {9'd85,10'd285};
ram[16541] = {9'd88,10'd289};
ram[16542] = {9'd91,10'd292};
ram[16543] = {9'd95,10'd295};
ram[16544] = {9'd98,10'd298};
ram[16545] = {-9'd99,10'd301};
ram[16546] = {-9'd96,10'd304};
ram[16547] = {-9'd93,10'd307};
ram[16548] = {-9'd90,10'd311};
ram[16549] = {-9'd87,10'd314};
ram[16550] = {-9'd84,10'd317};
ram[16551] = {-9'd81,10'd320};
ram[16552] = {-9'd77,10'd323};
ram[16553] = {-9'd74,10'd326};
ram[16554] = {-9'd71,10'd329};
ram[16555] = {-9'd68,10'd333};
ram[16556] = {-9'd65,10'd336};
ram[16557] = {-9'd62,10'd339};
ram[16558] = {-9'd59,10'd342};
ram[16559] = {-9'd55,10'd345};
ram[16560] = {-9'd52,10'd348};
ram[16561] = {-9'd49,10'd351};
ram[16562] = {-9'd46,10'd354};
ram[16563] = {-9'd43,10'd358};
ram[16564] = {-9'd40,10'd361};
ram[16565] = {-9'd37,10'd364};
ram[16566] = {-9'd33,10'd367};
ram[16567] = {-9'd30,10'd370};
ram[16568] = {-9'd27,10'd373};
ram[16569] = {-9'd24,10'd376};
ram[16570] = {-9'd21,10'd380};
ram[16571] = {-9'd18,10'd383};
ram[16572] = {-9'd15,10'd386};
ram[16573] = {-9'd11,10'd389};
ram[16574] = {-9'd8,10'd392};
ram[16575] = {-9'd5,10'd395};
ram[16576] = {-9'd2,10'd398};
ram[16577] = {9'd1,-10'd399};
ram[16578] = {9'd4,-10'd396};
ram[16579] = {9'd7,-10'd393};
ram[16580] = {9'd10,-10'd390};
ram[16581] = {9'd14,-10'd387};
ram[16582] = {9'd17,-10'd384};
ram[16583] = {9'd20,-10'd381};
ram[16584] = {9'd23,-10'd377};
ram[16585] = {9'd26,-10'd374};
ram[16586] = {9'd29,-10'd371};
ram[16587] = {9'd32,-10'd368};
ram[16588] = {9'd36,-10'd365};
ram[16589] = {9'd39,-10'd362};
ram[16590] = {9'd42,-10'd359};
ram[16591] = {9'd45,-10'd355};
ram[16592] = {9'd48,-10'd352};
ram[16593] = {9'd51,-10'd349};
ram[16594] = {9'd54,-10'd346};
ram[16595] = {9'd58,-10'd343};
ram[16596] = {9'd61,-10'd340};
ram[16597] = {9'd64,-10'd337};
ram[16598] = {9'd67,-10'd334};
ram[16599] = {9'd70,-10'd330};
ram[16600] = {9'd73,-10'd327};
ram[16601] = {9'd76,-10'd324};
ram[16602] = {9'd80,-10'd321};
ram[16603] = {9'd83,-10'd318};
ram[16604] = {9'd86,-10'd315};
ram[16605] = {9'd89,-10'd312};
ram[16606] = {9'd92,-10'd308};
ram[16607] = {9'd95,-10'd305};
ram[16608] = {9'd98,-10'd302};
ram[16609] = {-9'd99,-10'd299};
ram[16610] = {-9'd96,-10'd296};
ram[16611] = {-9'd92,-10'd293};
ram[16612] = {-9'd89,-10'd290};
ram[16613] = {-9'd86,-10'd286};
ram[16614] = {-9'd83,-10'd283};
ram[16615] = {-9'd80,-10'd280};
ram[16616] = {-9'd77,-10'd277};
ram[16617] = {-9'd74,-10'd274};
ram[16618] = {-9'd70,-10'd271};
ram[16619] = {-9'd67,-10'd268};
ram[16620] = {-9'd64,-10'd264};
ram[16621] = {-9'd61,-10'd261};
ram[16622] = {-9'd58,-10'd258};
ram[16623] = {-9'd55,-10'd255};
ram[16624] = {-9'd52,-10'd252};
ram[16625] = {-9'd48,-10'd249};
ram[16626] = {-9'd45,-10'd246};
ram[16627] = {-9'd42,-10'd242};
ram[16628] = {-9'd39,-10'd239};
ram[16629] = {-9'd36,-10'd236};
ram[16630] = {-9'd33,-10'd233};
ram[16631] = {-9'd30,-10'd230};
ram[16632] = {-9'd26,-10'd227};
ram[16633] = {-9'd23,-10'd224};
ram[16634] = {-9'd20,-10'd220};
ram[16635] = {-9'd17,-10'd217};
ram[16636] = {-9'd14,-10'd214};
ram[16637] = {-9'd11,-10'd211};
ram[16638] = {-9'd8,-10'd208};
ram[16639] = {-9'd4,-10'd205};
ram[16640] = {-9'd4,-10'd205};
ram[16641] = {-9'd1,-10'd202};
ram[16642] = {9'd2,-10'd198};
ram[16643] = {9'd5,-10'd195};
ram[16644] = {9'd8,-10'd192};
ram[16645] = {9'd11,-10'd189};
ram[16646] = {9'd14,-10'd186};
ram[16647] = {9'd18,-10'd183};
ram[16648] = {9'd21,-10'd180};
ram[16649] = {9'd24,-10'd176};
ram[16650] = {9'd27,-10'd173};
ram[16651] = {9'd30,-10'd170};
ram[16652] = {9'd33,-10'd167};
ram[16653] = {9'd36,-10'd164};
ram[16654] = {9'd40,-10'd161};
ram[16655] = {9'd43,-10'd158};
ram[16656] = {9'd46,-10'd154};
ram[16657] = {9'd49,-10'd151};
ram[16658] = {9'd52,-10'd148};
ram[16659] = {9'd55,-10'd145};
ram[16660] = {9'd58,-10'd142};
ram[16661] = {9'd62,-10'd139};
ram[16662] = {9'd65,-10'd136};
ram[16663] = {9'd68,-10'd132};
ram[16664] = {9'd71,-10'd129};
ram[16665] = {9'd74,-10'd126};
ram[16666] = {9'd77,-10'd123};
ram[16667] = {9'd80,-10'd120};
ram[16668] = {9'd84,-10'd117};
ram[16669] = {9'd87,-10'd114};
ram[16670] = {9'd90,-10'd110};
ram[16671] = {9'd93,-10'd107};
ram[16672] = {9'd96,-10'd104};
ram[16673] = {9'd99,-10'd101};
ram[16674] = {-9'd98,-10'd98};
ram[16675] = {-9'd95,-10'd95};
ram[16676] = {-9'd92,-10'd92};
ram[16677] = {-9'd88,-10'd88};
ram[16678] = {-9'd85,-10'd85};
ram[16679] = {-9'd82,-10'd82};
ram[16680] = {-9'd79,-10'd79};
ram[16681] = {-9'd76,-10'd76};
ram[16682] = {-9'd73,-10'd73};
ram[16683] = {-9'd70,-10'd70};
ram[16684] = {-9'd66,-10'd66};
ram[16685] = {-9'd63,-10'd63};
ram[16686] = {-9'd60,-10'd60};
ram[16687] = {-9'd57,-10'd57};
ram[16688] = {-9'd54,-10'd54};
ram[16689] = {-9'd51,-10'd51};
ram[16690] = {-9'd48,-10'd48};
ram[16691] = {-9'd44,-10'd44};
ram[16692] = {-9'd41,-10'd41};
ram[16693] = {-9'd38,-10'd38};
ram[16694] = {-9'd35,-10'd35};
ram[16695] = {-9'd32,-10'd32};
ram[16696] = {-9'd29,-10'd29};
ram[16697] = {-9'd26,-10'd26};
ram[16698] = {-9'd22,-10'd22};
ram[16699] = {-9'd19,-10'd19};
ram[16700] = {-9'd16,-10'd16};
ram[16701] = {-9'd13,-10'd13};
ram[16702] = {-9'd10,-10'd10};
ram[16703] = {-9'd7,-10'd7};
ram[16704] = {-9'd4,-10'd4};
ram[16705] = {9'd0,10'd0};
ram[16706] = {9'd3,10'd3};
ram[16707] = {9'd6,10'd6};
ram[16708] = {9'd9,10'd9};
ram[16709] = {9'd12,10'd12};
ram[16710] = {9'd15,10'd15};
ram[16711] = {9'd18,10'd18};
ram[16712] = {9'd21,10'd21};
ram[16713] = {9'd25,10'd25};
ram[16714] = {9'd28,10'd28};
ram[16715] = {9'd31,10'd31};
ram[16716] = {9'd34,10'd34};
ram[16717] = {9'd37,10'd37};
ram[16718] = {9'd40,10'd40};
ram[16719] = {9'd43,10'd43};
ram[16720] = {9'd47,10'd47};
ram[16721] = {9'd50,10'd50};
ram[16722] = {9'd53,10'd53};
ram[16723] = {9'd56,10'd56};
ram[16724] = {9'd59,10'd59};
ram[16725] = {9'd62,10'd62};
ram[16726] = {9'd65,10'd65};
ram[16727] = {9'd69,10'd69};
ram[16728] = {9'd72,10'd72};
ram[16729] = {9'd75,10'd75};
ram[16730] = {9'd78,10'd78};
ram[16731] = {9'd81,10'd81};
ram[16732] = {9'd84,10'd84};
ram[16733] = {9'd87,10'd87};
ram[16734] = {9'd91,10'd91};
ram[16735] = {9'd94,10'd94};
ram[16736] = {9'd97,10'd97};
ram[16737] = {-9'd100,10'd100};
ram[16738] = {-9'd97,10'd103};
ram[16739] = {-9'd94,10'd106};
ram[16740] = {-9'd91,10'd109};
ram[16741] = {-9'd88,10'd113};
ram[16742] = {-9'd85,10'd116};
ram[16743] = {-9'd81,10'd119};
ram[16744] = {-9'd78,10'd122};
ram[16745] = {-9'd75,10'd125};
ram[16746] = {-9'd72,10'd128};
ram[16747] = {-9'd69,10'd131};
ram[16748] = {-9'd66,10'd135};
ram[16749] = {-9'd63,10'd138};
ram[16750] = {-9'd59,10'd141};
ram[16751] = {-9'd56,10'd144};
ram[16752] = {-9'd53,10'd147};
ram[16753] = {-9'd50,10'd150};
ram[16754] = {-9'd47,10'd153};
ram[16755] = {-9'd44,10'd157};
ram[16756] = {-9'd41,10'd160};
ram[16757] = {-9'd37,10'd163};
ram[16758] = {-9'd34,10'd166};
ram[16759] = {-9'd31,10'd169};
ram[16760] = {-9'd28,10'd172};
ram[16761] = {-9'd25,10'd175};
ram[16762] = {-9'd22,10'd179};
ram[16763] = {-9'd19,10'd182};
ram[16764] = {-9'd15,10'd185};
ram[16765] = {-9'd12,10'd188};
ram[16766] = {-9'd9,10'd191};
ram[16767] = {-9'd6,10'd194};
ram[16768] = {-9'd6,10'd194};
ram[16769] = {-9'd3,10'd197};
ram[16770] = {9'd0,10'd201};
ram[16771] = {9'd3,10'd204};
ram[16772] = {9'd7,10'd207};
ram[16773] = {9'd10,10'd210};
ram[16774] = {9'd13,10'd213};
ram[16775] = {9'd16,10'd216};
ram[16776] = {9'd19,10'd219};
ram[16777] = {9'd22,10'd223};
ram[16778] = {9'd25,10'd226};
ram[16779] = {9'd29,10'd229};
ram[16780] = {9'd32,10'd232};
ram[16781] = {9'd35,10'd235};
ram[16782] = {9'd38,10'd238};
ram[16783] = {9'd41,10'd241};
ram[16784] = {9'd44,10'd245};
ram[16785] = {9'd47,10'd248};
ram[16786] = {9'd51,10'd251};
ram[16787] = {9'd54,10'd254};
ram[16788] = {9'd57,10'd257};
ram[16789] = {9'd60,10'd260};
ram[16790] = {9'd63,10'd263};
ram[16791] = {9'd66,10'd267};
ram[16792] = {9'd69,10'd270};
ram[16793] = {9'd73,10'd273};
ram[16794] = {9'd76,10'd276};
ram[16795] = {9'd79,10'd279};
ram[16796] = {9'd82,10'd282};
ram[16797] = {9'd85,10'd285};
ram[16798] = {9'd88,10'd289};
ram[16799] = {9'd91,10'd292};
ram[16800] = {9'd95,10'd295};
ram[16801] = {9'd98,10'd298};
ram[16802] = {-9'd99,10'd301};
ram[16803] = {-9'd96,10'd304};
ram[16804] = {-9'd93,10'd307};
ram[16805] = {-9'd90,10'd311};
ram[16806] = {-9'd87,10'd314};
ram[16807] = {-9'd84,10'd317};
ram[16808] = {-9'd81,10'd320};
ram[16809] = {-9'd77,10'd323};
ram[16810] = {-9'd74,10'd326};
ram[16811] = {-9'd71,10'd329};
ram[16812] = {-9'd68,10'd333};
ram[16813] = {-9'd65,10'd336};
ram[16814] = {-9'd62,10'd339};
ram[16815] = {-9'd59,10'd342};
ram[16816] = {-9'd55,10'd345};
ram[16817] = {-9'd52,10'd348};
ram[16818] = {-9'd49,10'd351};
ram[16819] = {-9'd46,10'd354};
ram[16820] = {-9'd43,10'd358};
ram[16821] = {-9'd40,10'd361};
ram[16822] = {-9'd37,10'd364};
ram[16823] = {-9'd33,10'd367};
ram[16824] = {-9'd30,10'd370};
ram[16825] = {-9'd27,10'd373};
ram[16826] = {-9'd24,10'd376};
ram[16827] = {-9'd21,10'd380};
ram[16828] = {-9'd18,10'd383};
ram[16829] = {-9'd15,10'd386};
ram[16830] = {-9'd11,10'd389};
ram[16831] = {-9'd8,10'd392};
ram[16832] = {-9'd5,10'd395};
ram[16833] = {-9'd2,10'd398};
ram[16834] = {9'd1,-10'd399};
ram[16835] = {9'd4,-10'd396};
ram[16836] = {9'd7,-10'd393};
ram[16837] = {9'd10,-10'd390};
ram[16838] = {9'd14,-10'd387};
ram[16839] = {9'd17,-10'd384};
ram[16840] = {9'd20,-10'd381};
ram[16841] = {9'd23,-10'd377};
ram[16842] = {9'd26,-10'd374};
ram[16843] = {9'd29,-10'd371};
ram[16844] = {9'd32,-10'd368};
ram[16845] = {9'd36,-10'd365};
ram[16846] = {9'd39,-10'd362};
ram[16847] = {9'd42,-10'd359};
ram[16848] = {9'd45,-10'd355};
ram[16849] = {9'd48,-10'd352};
ram[16850] = {9'd51,-10'd349};
ram[16851] = {9'd54,-10'd346};
ram[16852] = {9'd58,-10'd343};
ram[16853] = {9'd61,-10'd340};
ram[16854] = {9'd64,-10'd337};
ram[16855] = {9'd67,-10'd334};
ram[16856] = {9'd70,-10'd330};
ram[16857] = {9'd73,-10'd327};
ram[16858] = {9'd76,-10'd324};
ram[16859] = {9'd80,-10'd321};
ram[16860] = {9'd83,-10'd318};
ram[16861] = {9'd86,-10'd315};
ram[16862] = {9'd89,-10'd312};
ram[16863] = {9'd92,-10'd308};
ram[16864] = {9'd95,-10'd305};
ram[16865] = {9'd98,-10'd302};
ram[16866] = {-9'd99,-10'd299};
ram[16867] = {-9'd96,-10'd296};
ram[16868] = {-9'd92,-10'd293};
ram[16869] = {-9'd89,-10'd290};
ram[16870] = {-9'd86,-10'd286};
ram[16871] = {-9'd83,-10'd283};
ram[16872] = {-9'd80,-10'd280};
ram[16873] = {-9'd77,-10'd277};
ram[16874] = {-9'd74,-10'd274};
ram[16875] = {-9'd70,-10'd271};
ram[16876] = {-9'd67,-10'd268};
ram[16877] = {-9'd64,-10'd264};
ram[16878] = {-9'd61,-10'd261};
ram[16879] = {-9'd58,-10'd258};
ram[16880] = {-9'd55,-10'd255};
ram[16881] = {-9'd52,-10'd252};
ram[16882] = {-9'd48,-10'd249};
ram[16883] = {-9'd45,-10'd246};
ram[16884] = {-9'd42,-10'd242};
ram[16885] = {-9'd39,-10'd239};
ram[16886] = {-9'd36,-10'd236};
ram[16887] = {-9'd33,-10'd233};
ram[16888] = {-9'd30,-10'd230};
ram[16889] = {-9'd26,-10'd227};
ram[16890] = {-9'd23,-10'd224};
ram[16891] = {-9'd20,-10'd220};
ram[16892] = {-9'd17,-10'd217};
ram[16893] = {-9'd14,-10'd214};
ram[16894] = {-9'd11,-10'd211};
ram[16895] = {-9'd8,-10'd208};
ram[16896] = {-9'd8,-10'd208};
ram[16897] = {-9'd4,-10'd205};
ram[16898] = {-9'd1,-10'd202};
ram[16899] = {9'd2,-10'd198};
ram[16900] = {9'd5,-10'd195};
ram[16901] = {9'd8,-10'd192};
ram[16902] = {9'd11,-10'd189};
ram[16903] = {9'd14,-10'd186};
ram[16904] = {9'd18,-10'd183};
ram[16905] = {9'd21,-10'd180};
ram[16906] = {9'd24,-10'd176};
ram[16907] = {9'd27,-10'd173};
ram[16908] = {9'd30,-10'd170};
ram[16909] = {9'd33,-10'd167};
ram[16910] = {9'd36,-10'd164};
ram[16911] = {9'd40,-10'd161};
ram[16912] = {9'd43,-10'd158};
ram[16913] = {9'd46,-10'd154};
ram[16914] = {9'd49,-10'd151};
ram[16915] = {9'd52,-10'd148};
ram[16916] = {9'd55,-10'd145};
ram[16917] = {9'd58,-10'd142};
ram[16918] = {9'd62,-10'd139};
ram[16919] = {9'd65,-10'd136};
ram[16920] = {9'd68,-10'd132};
ram[16921] = {9'd71,-10'd129};
ram[16922] = {9'd74,-10'd126};
ram[16923] = {9'd77,-10'd123};
ram[16924] = {9'd80,-10'd120};
ram[16925] = {9'd84,-10'd117};
ram[16926] = {9'd87,-10'd114};
ram[16927] = {9'd90,-10'd110};
ram[16928] = {9'd93,-10'd107};
ram[16929] = {9'd96,-10'd104};
ram[16930] = {9'd99,-10'd101};
ram[16931] = {-9'd98,-10'd98};
ram[16932] = {-9'd95,-10'd95};
ram[16933] = {-9'd92,-10'd92};
ram[16934] = {-9'd88,-10'd88};
ram[16935] = {-9'd85,-10'd85};
ram[16936] = {-9'd82,-10'd82};
ram[16937] = {-9'd79,-10'd79};
ram[16938] = {-9'd76,-10'd76};
ram[16939] = {-9'd73,-10'd73};
ram[16940] = {-9'd70,-10'd70};
ram[16941] = {-9'd66,-10'd66};
ram[16942] = {-9'd63,-10'd63};
ram[16943] = {-9'd60,-10'd60};
ram[16944] = {-9'd57,-10'd57};
ram[16945] = {-9'd54,-10'd54};
ram[16946] = {-9'd51,-10'd51};
ram[16947] = {-9'd48,-10'd48};
ram[16948] = {-9'd44,-10'd44};
ram[16949] = {-9'd41,-10'd41};
ram[16950] = {-9'd38,-10'd38};
ram[16951] = {-9'd35,-10'd35};
ram[16952] = {-9'd32,-10'd32};
ram[16953] = {-9'd29,-10'd29};
ram[16954] = {-9'd26,-10'd26};
ram[16955] = {-9'd22,-10'd22};
ram[16956] = {-9'd19,-10'd19};
ram[16957] = {-9'd16,-10'd16};
ram[16958] = {-9'd13,-10'd13};
ram[16959] = {-9'd10,-10'd10};
ram[16960] = {-9'd7,-10'd7};
ram[16961] = {-9'd4,-10'd4};
ram[16962] = {9'd0,10'd0};
ram[16963] = {9'd3,10'd3};
ram[16964] = {9'd6,10'd6};
ram[16965] = {9'd9,10'd9};
ram[16966] = {9'd12,10'd12};
ram[16967] = {9'd15,10'd15};
ram[16968] = {9'd18,10'd18};
ram[16969] = {9'd21,10'd21};
ram[16970] = {9'd25,10'd25};
ram[16971] = {9'd28,10'd28};
ram[16972] = {9'd31,10'd31};
ram[16973] = {9'd34,10'd34};
ram[16974] = {9'd37,10'd37};
ram[16975] = {9'd40,10'd40};
ram[16976] = {9'd43,10'd43};
ram[16977] = {9'd47,10'd47};
ram[16978] = {9'd50,10'd50};
ram[16979] = {9'd53,10'd53};
ram[16980] = {9'd56,10'd56};
ram[16981] = {9'd59,10'd59};
ram[16982] = {9'd62,10'd62};
ram[16983] = {9'd65,10'd65};
ram[16984] = {9'd69,10'd69};
ram[16985] = {9'd72,10'd72};
ram[16986] = {9'd75,10'd75};
ram[16987] = {9'd78,10'd78};
ram[16988] = {9'd81,10'd81};
ram[16989] = {9'd84,10'd84};
ram[16990] = {9'd87,10'd87};
ram[16991] = {9'd91,10'd91};
ram[16992] = {9'd94,10'd94};
ram[16993] = {9'd97,10'd97};
ram[16994] = {-9'd100,10'd100};
ram[16995] = {-9'd97,10'd103};
ram[16996] = {-9'd94,10'd106};
ram[16997] = {-9'd91,10'd109};
ram[16998] = {-9'd88,10'd113};
ram[16999] = {-9'd85,10'd116};
ram[17000] = {-9'd81,10'd119};
ram[17001] = {-9'd78,10'd122};
ram[17002] = {-9'd75,10'd125};
ram[17003] = {-9'd72,10'd128};
ram[17004] = {-9'd69,10'd131};
ram[17005] = {-9'd66,10'd135};
ram[17006] = {-9'd63,10'd138};
ram[17007] = {-9'd59,10'd141};
ram[17008] = {-9'd56,10'd144};
ram[17009] = {-9'd53,10'd147};
ram[17010] = {-9'd50,10'd150};
ram[17011] = {-9'd47,10'd153};
ram[17012] = {-9'd44,10'd157};
ram[17013] = {-9'd41,10'd160};
ram[17014] = {-9'd37,10'd163};
ram[17015] = {-9'd34,10'd166};
ram[17016] = {-9'd31,10'd169};
ram[17017] = {-9'd28,10'd172};
ram[17018] = {-9'd25,10'd175};
ram[17019] = {-9'd22,10'd179};
ram[17020] = {-9'd19,10'd182};
ram[17021] = {-9'd15,10'd185};
ram[17022] = {-9'd12,10'd188};
ram[17023] = {-9'd9,10'd191};
ram[17024] = {-9'd9,10'd191};
ram[17025] = {-9'd6,10'd194};
ram[17026] = {-9'd3,10'd197};
ram[17027] = {9'd0,10'd201};
ram[17028] = {9'd3,10'd204};
ram[17029] = {9'd7,10'd207};
ram[17030] = {9'd10,10'd210};
ram[17031] = {9'd13,10'd213};
ram[17032] = {9'd16,10'd216};
ram[17033] = {9'd19,10'd219};
ram[17034] = {9'd22,10'd223};
ram[17035] = {9'd25,10'd226};
ram[17036] = {9'd29,10'd229};
ram[17037] = {9'd32,10'd232};
ram[17038] = {9'd35,10'd235};
ram[17039] = {9'd38,10'd238};
ram[17040] = {9'd41,10'd241};
ram[17041] = {9'd44,10'd245};
ram[17042] = {9'd47,10'd248};
ram[17043] = {9'd51,10'd251};
ram[17044] = {9'd54,10'd254};
ram[17045] = {9'd57,10'd257};
ram[17046] = {9'd60,10'd260};
ram[17047] = {9'd63,10'd263};
ram[17048] = {9'd66,10'd267};
ram[17049] = {9'd69,10'd270};
ram[17050] = {9'd73,10'd273};
ram[17051] = {9'd76,10'd276};
ram[17052] = {9'd79,10'd279};
ram[17053] = {9'd82,10'd282};
ram[17054] = {9'd85,10'd285};
ram[17055] = {9'd88,10'd289};
ram[17056] = {9'd91,10'd292};
ram[17057] = {9'd95,10'd295};
ram[17058] = {9'd98,10'd298};
ram[17059] = {-9'd99,10'd301};
ram[17060] = {-9'd96,10'd304};
ram[17061] = {-9'd93,10'd307};
ram[17062] = {-9'd90,10'd311};
ram[17063] = {-9'd87,10'd314};
ram[17064] = {-9'd84,10'd317};
ram[17065] = {-9'd81,10'd320};
ram[17066] = {-9'd77,10'd323};
ram[17067] = {-9'd74,10'd326};
ram[17068] = {-9'd71,10'd329};
ram[17069] = {-9'd68,10'd333};
ram[17070] = {-9'd65,10'd336};
ram[17071] = {-9'd62,10'd339};
ram[17072] = {-9'd59,10'd342};
ram[17073] = {-9'd55,10'd345};
ram[17074] = {-9'd52,10'd348};
ram[17075] = {-9'd49,10'd351};
ram[17076] = {-9'd46,10'd354};
ram[17077] = {-9'd43,10'd358};
ram[17078] = {-9'd40,10'd361};
ram[17079] = {-9'd37,10'd364};
ram[17080] = {-9'd33,10'd367};
ram[17081] = {-9'd30,10'd370};
ram[17082] = {-9'd27,10'd373};
ram[17083] = {-9'd24,10'd376};
ram[17084] = {-9'd21,10'd380};
ram[17085] = {-9'd18,10'd383};
ram[17086] = {-9'd15,10'd386};
ram[17087] = {-9'd11,10'd389};
ram[17088] = {-9'd8,10'd392};
ram[17089] = {-9'd5,10'd395};
ram[17090] = {-9'd2,10'd398};
ram[17091] = {9'd1,-10'd399};
ram[17092] = {9'd4,-10'd396};
ram[17093] = {9'd7,-10'd393};
ram[17094] = {9'd10,-10'd390};
ram[17095] = {9'd14,-10'd387};
ram[17096] = {9'd17,-10'd384};
ram[17097] = {9'd20,-10'd381};
ram[17098] = {9'd23,-10'd377};
ram[17099] = {9'd26,-10'd374};
ram[17100] = {9'd29,-10'd371};
ram[17101] = {9'd32,-10'd368};
ram[17102] = {9'd36,-10'd365};
ram[17103] = {9'd39,-10'd362};
ram[17104] = {9'd42,-10'd359};
ram[17105] = {9'd45,-10'd355};
ram[17106] = {9'd48,-10'd352};
ram[17107] = {9'd51,-10'd349};
ram[17108] = {9'd54,-10'd346};
ram[17109] = {9'd58,-10'd343};
ram[17110] = {9'd61,-10'd340};
ram[17111] = {9'd64,-10'd337};
ram[17112] = {9'd67,-10'd334};
ram[17113] = {9'd70,-10'd330};
ram[17114] = {9'd73,-10'd327};
ram[17115] = {9'd76,-10'd324};
ram[17116] = {9'd80,-10'd321};
ram[17117] = {9'd83,-10'd318};
ram[17118] = {9'd86,-10'd315};
ram[17119] = {9'd89,-10'd312};
ram[17120] = {9'd92,-10'd308};
ram[17121] = {9'd95,-10'd305};
ram[17122] = {9'd98,-10'd302};
ram[17123] = {-9'd99,-10'd299};
ram[17124] = {-9'd96,-10'd296};
ram[17125] = {-9'd92,-10'd293};
ram[17126] = {-9'd89,-10'd290};
ram[17127] = {-9'd86,-10'd286};
ram[17128] = {-9'd83,-10'd283};
ram[17129] = {-9'd80,-10'd280};
ram[17130] = {-9'd77,-10'd277};
ram[17131] = {-9'd74,-10'd274};
ram[17132] = {-9'd70,-10'd271};
ram[17133] = {-9'd67,-10'd268};
ram[17134] = {-9'd64,-10'd264};
ram[17135] = {-9'd61,-10'd261};
ram[17136] = {-9'd58,-10'd258};
ram[17137] = {-9'd55,-10'd255};
ram[17138] = {-9'd52,-10'd252};
ram[17139] = {-9'd48,-10'd249};
ram[17140] = {-9'd45,-10'd246};
ram[17141] = {-9'd42,-10'd242};
ram[17142] = {-9'd39,-10'd239};
ram[17143] = {-9'd36,-10'd236};
ram[17144] = {-9'd33,-10'd233};
ram[17145] = {-9'd30,-10'd230};
ram[17146] = {-9'd26,-10'd227};
ram[17147] = {-9'd23,-10'd224};
ram[17148] = {-9'd20,-10'd220};
ram[17149] = {-9'd17,-10'd217};
ram[17150] = {-9'd14,-10'd214};
ram[17151] = {-9'd11,-10'd211};
ram[17152] = {-9'd11,-10'd211};
ram[17153] = {-9'd8,-10'd208};
ram[17154] = {-9'd4,-10'd205};
ram[17155] = {-9'd1,-10'd202};
ram[17156] = {9'd2,-10'd198};
ram[17157] = {9'd5,-10'd195};
ram[17158] = {9'd8,-10'd192};
ram[17159] = {9'd11,-10'd189};
ram[17160] = {9'd14,-10'd186};
ram[17161] = {9'd18,-10'd183};
ram[17162] = {9'd21,-10'd180};
ram[17163] = {9'd24,-10'd176};
ram[17164] = {9'd27,-10'd173};
ram[17165] = {9'd30,-10'd170};
ram[17166] = {9'd33,-10'd167};
ram[17167] = {9'd36,-10'd164};
ram[17168] = {9'd40,-10'd161};
ram[17169] = {9'd43,-10'd158};
ram[17170] = {9'd46,-10'd154};
ram[17171] = {9'd49,-10'd151};
ram[17172] = {9'd52,-10'd148};
ram[17173] = {9'd55,-10'd145};
ram[17174] = {9'd58,-10'd142};
ram[17175] = {9'd62,-10'd139};
ram[17176] = {9'd65,-10'd136};
ram[17177] = {9'd68,-10'd132};
ram[17178] = {9'd71,-10'd129};
ram[17179] = {9'd74,-10'd126};
ram[17180] = {9'd77,-10'd123};
ram[17181] = {9'd80,-10'd120};
ram[17182] = {9'd84,-10'd117};
ram[17183] = {9'd87,-10'd114};
ram[17184] = {9'd90,-10'd110};
ram[17185] = {9'd93,-10'd107};
ram[17186] = {9'd96,-10'd104};
ram[17187] = {9'd99,-10'd101};
ram[17188] = {-9'd98,-10'd98};
ram[17189] = {-9'd95,-10'd95};
ram[17190] = {-9'd92,-10'd92};
ram[17191] = {-9'd88,-10'd88};
ram[17192] = {-9'd85,-10'd85};
ram[17193] = {-9'd82,-10'd82};
ram[17194] = {-9'd79,-10'd79};
ram[17195] = {-9'd76,-10'd76};
ram[17196] = {-9'd73,-10'd73};
ram[17197] = {-9'd70,-10'd70};
ram[17198] = {-9'd66,-10'd66};
ram[17199] = {-9'd63,-10'd63};
ram[17200] = {-9'd60,-10'd60};
ram[17201] = {-9'd57,-10'd57};
ram[17202] = {-9'd54,-10'd54};
ram[17203] = {-9'd51,-10'd51};
ram[17204] = {-9'd48,-10'd48};
ram[17205] = {-9'd44,-10'd44};
ram[17206] = {-9'd41,-10'd41};
ram[17207] = {-9'd38,-10'd38};
ram[17208] = {-9'd35,-10'd35};
ram[17209] = {-9'd32,-10'd32};
ram[17210] = {-9'd29,-10'd29};
ram[17211] = {-9'd26,-10'd26};
ram[17212] = {-9'd22,-10'd22};
ram[17213] = {-9'd19,-10'd19};
ram[17214] = {-9'd16,-10'd16};
ram[17215] = {-9'd13,-10'd13};
ram[17216] = {-9'd10,-10'd10};
ram[17217] = {-9'd7,-10'd7};
ram[17218] = {-9'd4,-10'd4};
ram[17219] = {9'd0,10'd0};
ram[17220] = {9'd3,10'd3};
ram[17221] = {9'd6,10'd6};
ram[17222] = {9'd9,10'd9};
ram[17223] = {9'd12,10'd12};
ram[17224] = {9'd15,10'd15};
ram[17225] = {9'd18,10'd18};
ram[17226] = {9'd21,10'd21};
ram[17227] = {9'd25,10'd25};
ram[17228] = {9'd28,10'd28};
ram[17229] = {9'd31,10'd31};
ram[17230] = {9'd34,10'd34};
ram[17231] = {9'd37,10'd37};
ram[17232] = {9'd40,10'd40};
ram[17233] = {9'd43,10'd43};
ram[17234] = {9'd47,10'd47};
ram[17235] = {9'd50,10'd50};
ram[17236] = {9'd53,10'd53};
ram[17237] = {9'd56,10'd56};
ram[17238] = {9'd59,10'd59};
ram[17239] = {9'd62,10'd62};
ram[17240] = {9'd65,10'd65};
ram[17241] = {9'd69,10'd69};
ram[17242] = {9'd72,10'd72};
ram[17243] = {9'd75,10'd75};
ram[17244] = {9'd78,10'd78};
ram[17245] = {9'd81,10'd81};
ram[17246] = {9'd84,10'd84};
ram[17247] = {9'd87,10'd87};
ram[17248] = {9'd91,10'd91};
ram[17249] = {9'd94,10'd94};
ram[17250] = {9'd97,10'd97};
ram[17251] = {-9'd100,10'd100};
ram[17252] = {-9'd97,10'd103};
ram[17253] = {-9'd94,10'd106};
ram[17254] = {-9'd91,10'd109};
ram[17255] = {-9'd88,10'd113};
ram[17256] = {-9'd85,10'd116};
ram[17257] = {-9'd81,10'd119};
ram[17258] = {-9'd78,10'd122};
ram[17259] = {-9'd75,10'd125};
ram[17260] = {-9'd72,10'd128};
ram[17261] = {-9'd69,10'd131};
ram[17262] = {-9'd66,10'd135};
ram[17263] = {-9'd63,10'd138};
ram[17264] = {-9'd59,10'd141};
ram[17265] = {-9'd56,10'd144};
ram[17266] = {-9'd53,10'd147};
ram[17267] = {-9'd50,10'd150};
ram[17268] = {-9'd47,10'd153};
ram[17269] = {-9'd44,10'd157};
ram[17270] = {-9'd41,10'd160};
ram[17271] = {-9'd37,10'd163};
ram[17272] = {-9'd34,10'd166};
ram[17273] = {-9'd31,10'd169};
ram[17274] = {-9'd28,10'd172};
ram[17275] = {-9'd25,10'd175};
ram[17276] = {-9'd22,10'd179};
ram[17277] = {-9'd19,10'd182};
ram[17278] = {-9'd15,10'd185};
ram[17279] = {-9'd12,10'd188};
ram[17280] = {-9'd12,10'd188};
ram[17281] = {-9'd9,10'd191};
ram[17282] = {-9'd6,10'd194};
ram[17283] = {-9'd3,10'd197};
ram[17284] = {9'd0,10'd201};
ram[17285] = {9'd3,10'd204};
ram[17286] = {9'd7,10'd207};
ram[17287] = {9'd10,10'd210};
ram[17288] = {9'd13,10'd213};
ram[17289] = {9'd16,10'd216};
ram[17290] = {9'd19,10'd219};
ram[17291] = {9'd22,10'd223};
ram[17292] = {9'd25,10'd226};
ram[17293] = {9'd29,10'd229};
ram[17294] = {9'd32,10'd232};
ram[17295] = {9'd35,10'd235};
ram[17296] = {9'd38,10'd238};
ram[17297] = {9'd41,10'd241};
ram[17298] = {9'd44,10'd245};
ram[17299] = {9'd47,10'd248};
ram[17300] = {9'd51,10'd251};
ram[17301] = {9'd54,10'd254};
ram[17302] = {9'd57,10'd257};
ram[17303] = {9'd60,10'd260};
ram[17304] = {9'd63,10'd263};
ram[17305] = {9'd66,10'd267};
ram[17306] = {9'd69,10'd270};
ram[17307] = {9'd73,10'd273};
ram[17308] = {9'd76,10'd276};
ram[17309] = {9'd79,10'd279};
ram[17310] = {9'd82,10'd282};
ram[17311] = {9'd85,10'd285};
ram[17312] = {9'd88,10'd289};
ram[17313] = {9'd91,10'd292};
ram[17314] = {9'd95,10'd295};
ram[17315] = {9'd98,10'd298};
ram[17316] = {-9'd99,10'd301};
ram[17317] = {-9'd96,10'd304};
ram[17318] = {-9'd93,10'd307};
ram[17319] = {-9'd90,10'd311};
ram[17320] = {-9'd87,10'd314};
ram[17321] = {-9'd84,10'd317};
ram[17322] = {-9'd81,10'd320};
ram[17323] = {-9'd77,10'd323};
ram[17324] = {-9'd74,10'd326};
ram[17325] = {-9'd71,10'd329};
ram[17326] = {-9'd68,10'd333};
ram[17327] = {-9'd65,10'd336};
ram[17328] = {-9'd62,10'd339};
ram[17329] = {-9'd59,10'd342};
ram[17330] = {-9'd55,10'd345};
ram[17331] = {-9'd52,10'd348};
ram[17332] = {-9'd49,10'd351};
ram[17333] = {-9'd46,10'd354};
ram[17334] = {-9'd43,10'd358};
ram[17335] = {-9'd40,10'd361};
ram[17336] = {-9'd37,10'd364};
ram[17337] = {-9'd33,10'd367};
ram[17338] = {-9'd30,10'd370};
ram[17339] = {-9'd27,10'd373};
ram[17340] = {-9'd24,10'd376};
ram[17341] = {-9'd21,10'd380};
ram[17342] = {-9'd18,10'd383};
ram[17343] = {-9'd15,10'd386};
ram[17344] = {-9'd11,10'd389};
ram[17345] = {-9'd8,10'd392};
ram[17346] = {-9'd5,10'd395};
ram[17347] = {-9'd2,10'd398};
ram[17348] = {9'd1,-10'd399};
ram[17349] = {9'd4,-10'd396};
ram[17350] = {9'd7,-10'd393};
ram[17351] = {9'd10,-10'd390};
ram[17352] = {9'd14,-10'd387};
ram[17353] = {9'd17,-10'd384};
ram[17354] = {9'd20,-10'd381};
ram[17355] = {9'd23,-10'd377};
ram[17356] = {9'd26,-10'd374};
ram[17357] = {9'd29,-10'd371};
ram[17358] = {9'd32,-10'd368};
ram[17359] = {9'd36,-10'd365};
ram[17360] = {9'd39,-10'd362};
ram[17361] = {9'd42,-10'd359};
ram[17362] = {9'd45,-10'd355};
ram[17363] = {9'd48,-10'd352};
ram[17364] = {9'd51,-10'd349};
ram[17365] = {9'd54,-10'd346};
ram[17366] = {9'd58,-10'd343};
ram[17367] = {9'd61,-10'd340};
ram[17368] = {9'd64,-10'd337};
ram[17369] = {9'd67,-10'd334};
ram[17370] = {9'd70,-10'd330};
ram[17371] = {9'd73,-10'd327};
ram[17372] = {9'd76,-10'd324};
ram[17373] = {9'd80,-10'd321};
ram[17374] = {9'd83,-10'd318};
ram[17375] = {9'd86,-10'd315};
ram[17376] = {9'd89,-10'd312};
ram[17377] = {9'd92,-10'd308};
ram[17378] = {9'd95,-10'd305};
ram[17379] = {9'd98,-10'd302};
ram[17380] = {-9'd99,-10'd299};
ram[17381] = {-9'd96,-10'd296};
ram[17382] = {-9'd92,-10'd293};
ram[17383] = {-9'd89,-10'd290};
ram[17384] = {-9'd86,-10'd286};
ram[17385] = {-9'd83,-10'd283};
ram[17386] = {-9'd80,-10'd280};
ram[17387] = {-9'd77,-10'd277};
ram[17388] = {-9'd74,-10'd274};
ram[17389] = {-9'd70,-10'd271};
ram[17390] = {-9'd67,-10'd268};
ram[17391] = {-9'd64,-10'd264};
ram[17392] = {-9'd61,-10'd261};
ram[17393] = {-9'd58,-10'd258};
ram[17394] = {-9'd55,-10'd255};
ram[17395] = {-9'd52,-10'd252};
ram[17396] = {-9'd48,-10'd249};
ram[17397] = {-9'd45,-10'd246};
ram[17398] = {-9'd42,-10'd242};
ram[17399] = {-9'd39,-10'd239};
ram[17400] = {-9'd36,-10'd236};
ram[17401] = {-9'd33,-10'd233};
ram[17402] = {-9'd30,-10'd230};
ram[17403] = {-9'd26,-10'd227};
ram[17404] = {-9'd23,-10'd224};
ram[17405] = {-9'd20,-10'd220};
ram[17406] = {-9'd17,-10'd217};
ram[17407] = {-9'd14,-10'd214};
ram[17408] = {-9'd14,-10'd214};
ram[17409] = {-9'd11,-10'd211};
ram[17410] = {-9'd8,-10'd208};
ram[17411] = {-9'd4,-10'd205};
ram[17412] = {-9'd1,-10'd202};
ram[17413] = {9'd2,-10'd198};
ram[17414] = {9'd5,-10'd195};
ram[17415] = {9'd8,-10'd192};
ram[17416] = {9'd11,-10'd189};
ram[17417] = {9'd14,-10'd186};
ram[17418] = {9'd18,-10'd183};
ram[17419] = {9'd21,-10'd180};
ram[17420] = {9'd24,-10'd176};
ram[17421] = {9'd27,-10'd173};
ram[17422] = {9'd30,-10'd170};
ram[17423] = {9'd33,-10'd167};
ram[17424] = {9'd36,-10'd164};
ram[17425] = {9'd40,-10'd161};
ram[17426] = {9'd43,-10'd158};
ram[17427] = {9'd46,-10'd154};
ram[17428] = {9'd49,-10'd151};
ram[17429] = {9'd52,-10'd148};
ram[17430] = {9'd55,-10'd145};
ram[17431] = {9'd58,-10'd142};
ram[17432] = {9'd62,-10'd139};
ram[17433] = {9'd65,-10'd136};
ram[17434] = {9'd68,-10'd132};
ram[17435] = {9'd71,-10'd129};
ram[17436] = {9'd74,-10'd126};
ram[17437] = {9'd77,-10'd123};
ram[17438] = {9'd80,-10'd120};
ram[17439] = {9'd84,-10'd117};
ram[17440] = {9'd87,-10'd114};
ram[17441] = {9'd90,-10'd110};
ram[17442] = {9'd93,-10'd107};
ram[17443] = {9'd96,-10'd104};
ram[17444] = {9'd99,-10'd101};
ram[17445] = {-9'd98,-10'd98};
ram[17446] = {-9'd95,-10'd95};
ram[17447] = {-9'd92,-10'd92};
ram[17448] = {-9'd88,-10'd88};
ram[17449] = {-9'd85,-10'd85};
ram[17450] = {-9'd82,-10'd82};
ram[17451] = {-9'd79,-10'd79};
ram[17452] = {-9'd76,-10'd76};
ram[17453] = {-9'd73,-10'd73};
ram[17454] = {-9'd70,-10'd70};
ram[17455] = {-9'd66,-10'd66};
ram[17456] = {-9'd63,-10'd63};
ram[17457] = {-9'd60,-10'd60};
ram[17458] = {-9'd57,-10'd57};
ram[17459] = {-9'd54,-10'd54};
ram[17460] = {-9'd51,-10'd51};
ram[17461] = {-9'd48,-10'd48};
ram[17462] = {-9'd44,-10'd44};
ram[17463] = {-9'd41,-10'd41};
ram[17464] = {-9'd38,-10'd38};
ram[17465] = {-9'd35,-10'd35};
ram[17466] = {-9'd32,-10'd32};
ram[17467] = {-9'd29,-10'd29};
ram[17468] = {-9'd26,-10'd26};
ram[17469] = {-9'd22,-10'd22};
ram[17470] = {-9'd19,-10'd19};
ram[17471] = {-9'd16,-10'd16};
ram[17472] = {-9'd13,-10'd13};
ram[17473] = {-9'd10,-10'd10};
ram[17474] = {-9'd7,-10'd7};
ram[17475] = {-9'd4,-10'd4};
ram[17476] = {9'd0,10'd0};
ram[17477] = {9'd3,10'd3};
ram[17478] = {9'd6,10'd6};
ram[17479] = {9'd9,10'd9};
ram[17480] = {9'd12,10'd12};
ram[17481] = {9'd15,10'd15};
ram[17482] = {9'd18,10'd18};
ram[17483] = {9'd21,10'd21};
ram[17484] = {9'd25,10'd25};
ram[17485] = {9'd28,10'd28};
ram[17486] = {9'd31,10'd31};
ram[17487] = {9'd34,10'd34};
ram[17488] = {9'd37,10'd37};
ram[17489] = {9'd40,10'd40};
ram[17490] = {9'd43,10'd43};
ram[17491] = {9'd47,10'd47};
ram[17492] = {9'd50,10'd50};
ram[17493] = {9'd53,10'd53};
ram[17494] = {9'd56,10'd56};
ram[17495] = {9'd59,10'd59};
ram[17496] = {9'd62,10'd62};
ram[17497] = {9'd65,10'd65};
ram[17498] = {9'd69,10'd69};
ram[17499] = {9'd72,10'd72};
ram[17500] = {9'd75,10'd75};
ram[17501] = {9'd78,10'd78};
ram[17502] = {9'd81,10'd81};
ram[17503] = {9'd84,10'd84};
ram[17504] = {9'd87,10'd87};
ram[17505] = {9'd91,10'd91};
ram[17506] = {9'd94,10'd94};
ram[17507] = {9'd97,10'd97};
ram[17508] = {-9'd100,10'd100};
ram[17509] = {-9'd97,10'd103};
ram[17510] = {-9'd94,10'd106};
ram[17511] = {-9'd91,10'd109};
ram[17512] = {-9'd88,10'd113};
ram[17513] = {-9'd85,10'd116};
ram[17514] = {-9'd81,10'd119};
ram[17515] = {-9'd78,10'd122};
ram[17516] = {-9'd75,10'd125};
ram[17517] = {-9'd72,10'd128};
ram[17518] = {-9'd69,10'd131};
ram[17519] = {-9'd66,10'd135};
ram[17520] = {-9'd63,10'd138};
ram[17521] = {-9'd59,10'd141};
ram[17522] = {-9'd56,10'd144};
ram[17523] = {-9'd53,10'd147};
ram[17524] = {-9'd50,10'd150};
ram[17525] = {-9'd47,10'd153};
ram[17526] = {-9'd44,10'd157};
ram[17527] = {-9'd41,10'd160};
ram[17528] = {-9'd37,10'd163};
ram[17529] = {-9'd34,10'd166};
ram[17530] = {-9'd31,10'd169};
ram[17531] = {-9'd28,10'd172};
ram[17532] = {-9'd25,10'd175};
ram[17533] = {-9'd22,10'd179};
ram[17534] = {-9'd19,10'd182};
ram[17535] = {-9'd15,10'd185};
ram[17536] = {-9'd15,10'd185};
ram[17537] = {-9'd12,10'd188};
ram[17538] = {-9'd9,10'd191};
ram[17539] = {-9'd6,10'd194};
ram[17540] = {-9'd3,10'd197};
ram[17541] = {9'd0,10'd201};
ram[17542] = {9'd3,10'd204};
ram[17543] = {9'd7,10'd207};
ram[17544] = {9'd10,10'd210};
ram[17545] = {9'd13,10'd213};
ram[17546] = {9'd16,10'd216};
ram[17547] = {9'd19,10'd219};
ram[17548] = {9'd22,10'd223};
ram[17549] = {9'd25,10'd226};
ram[17550] = {9'd29,10'd229};
ram[17551] = {9'd32,10'd232};
ram[17552] = {9'd35,10'd235};
ram[17553] = {9'd38,10'd238};
ram[17554] = {9'd41,10'd241};
ram[17555] = {9'd44,10'd245};
ram[17556] = {9'd47,10'd248};
ram[17557] = {9'd51,10'd251};
ram[17558] = {9'd54,10'd254};
ram[17559] = {9'd57,10'd257};
ram[17560] = {9'd60,10'd260};
ram[17561] = {9'd63,10'd263};
ram[17562] = {9'd66,10'd267};
ram[17563] = {9'd69,10'd270};
ram[17564] = {9'd73,10'd273};
ram[17565] = {9'd76,10'd276};
ram[17566] = {9'd79,10'd279};
ram[17567] = {9'd82,10'd282};
ram[17568] = {9'd85,10'd285};
ram[17569] = {9'd88,10'd289};
ram[17570] = {9'd91,10'd292};
ram[17571] = {9'd95,10'd295};
ram[17572] = {9'd98,10'd298};
ram[17573] = {-9'd99,10'd301};
ram[17574] = {-9'd96,10'd304};
ram[17575] = {-9'd93,10'd307};
ram[17576] = {-9'd90,10'd311};
ram[17577] = {-9'd87,10'd314};
ram[17578] = {-9'd84,10'd317};
ram[17579] = {-9'd81,10'd320};
ram[17580] = {-9'd77,10'd323};
ram[17581] = {-9'd74,10'd326};
ram[17582] = {-9'd71,10'd329};
ram[17583] = {-9'd68,10'd333};
ram[17584] = {-9'd65,10'd336};
ram[17585] = {-9'd62,10'd339};
ram[17586] = {-9'd59,10'd342};
ram[17587] = {-9'd55,10'd345};
ram[17588] = {-9'd52,10'd348};
ram[17589] = {-9'd49,10'd351};
ram[17590] = {-9'd46,10'd354};
ram[17591] = {-9'd43,10'd358};
ram[17592] = {-9'd40,10'd361};
ram[17593] = {-9'd37,10'd364};
ram[17594] = {-9'd33,10'd367};
ram[17595] = {-9'd30,10'd370};
ram[17596] = {-9'd27,10'd373};
ram[17597] = {-9'd24,10'd376};
ram[17598] = {-9'd21,10'd380};
ram[17599] = {-9'd18,10'd383};
ram[17600] = {-9'd15,10'd386};
ram[17601] = {-9'd11,10'd389};
ram[17602] = {-9'd8,10'd392};
ram[17603] = {-9'd5,10'd395};
ram[17604] = {-9'd2,10'd398};
ram[17605] = {9'd1,-10'd399};
ram[17606] = {9'd4,-10'd396};
ram[17607] = {9'd7,-10'd393};
ram[17608] = {9'd10,-10'd390};
ram[17609] = {9'd14,-10'd387};
ram[17610] = {9'd17,-10'd384};
ram[17611] = {9'd20,-10'd381};
ram[17612] = {9'd23,-10'd377};
ram[17613] = {9'd26,-10'd374};
ram[17614] = {9'd29,-10'd371};
ram[17615] = {9'd32,-10'd368};
ram[17616] = {9'd36,-10'd365};
ram[17617] = {9'd39,-10'd362};
ram[17618] = {9'd42,-10'd359};
ram[17619] = {9'd45,-10'd355};
ram[17620] = {9'd48,-10'd352};
ram[17621] = {9'd51,-10'd349};
ram[17622] = {9'd54,-10'd346};
ram[17623] = {9'd58,-10'd343};
ram[17624] = {9'd61,-10'd340};
ram[17625] = {9'd64,-10'd337};
ram[17626] = {9'd67,-10'd334};
ram[17627] = {9'd70,-10'd330};
ram[17628] = {9'd73,-10'd327};
ram[17629] = {9'd76,-10'd324};
ram[17630] = {9'd80,-10'd321};
ram[17631] = {9'd83,-10'd318};
ram[17632] = {9'd86,-10'd315};
ram[17633] = {9'd89,-10'd312};
ram[17634] = {9'd92,-10'd308};
ram[17635] = {9'd95,-10'd305};
ram[17636] = {9'd98,-10'd302};
ram[17637] = {-9'd99,-10'd299};
ram[17638] = {-9'd96,-10'd296};
ram[17639] = {-9'd92,-10'd293};
ram[17640] = {-9'd89,-10'd290};
ram[17641] = {-9'd86,-10'd286};
ram[17642] = {-9'd83,-10'd283};
ram[17643] = {-9'd80,-10'd280};
ram[17644] = {-9'd77,-10'd277};
ram[17645] = {-9'd74,-10'd274};
ram[17646] = {-9'd70,-10'd271};
ram[17647] = {-9'd67,-10'd268};
ram[17648] = {-9'd64,-10'd264};
ram[17649] = {-9'd61,-10'd261};
ram[17650] = {-9'd58,-10'd258};
ram[17651] = {-9'd55,-10'd255};
ram[17652] = {-9'd52,-10'd252};
ram[17653] = {-9'd48,-10'd249};
ram[17654] = {-9'd45,-10'd246};
ram[17655] = {-9'd42,-10'd242};
ram[17656] = {-9'd39,-10'd239};
ram[17657] = {-9'd36,-10'd236};
ram[17658] = {-9'd33,-10'd233};
ram[17659] = {-9'd30,-10'd230};
ram[17660] = {-9'd26,-10'd227};
ram[17661] = {-9'd23,-10'd224};
ram[17662] = {-9'd20,-10'd220};
ram[17663] = {-9'd17,-10'd217};
ram[17664] = {-9'd17,-10'd217};
ram[17665] = {-9'd14,-10'd214};
ram[17666] = {-9'd11,-10'd211};
ram[17667] = {-9'd8,-10'd208};
ram[17668] = {-9'd4,-10'd205};
ram[17669] = {-9'd1,-10'd202};
ram[17670] = {9'd2,-10'd198};
ram[17671] = {9'd5,-10'd195};
ram[17672] = {9'd8,-10'd192};
ram[17673] = {9'd11,-10'd189};
ram[17674] = {9'd14,-10'd186};
ram[17675] = {9'd18,-10'd183};
ram[17676] = {9'd21,-10'd180};
ram[17677] = {9'd24,-10'd176};
ram[17678] = {9'd27,-10'd173};
ram[17679] = {9'd30,-10'd170};
ram[17680] = {9'd33,-10'd167};
ram[17681] = {9'd36,-10'd164};
ram[17682] = {9'd40,-10'd161};
ram[17683] = {9'd43,-10'd158};
ram[17684] = {9'd46,-10'd154};
ram[17685] = {9'd49,-10'd151};
ram[17686] = {9'd52,-10'd148};
ram[17687] = {9'd55,-10'd145};
ram[17688] = {9'd58,-10'd142};
ram[17689] = {9'd62,-10'd139};
ram[17690] = {9'd65,-10'd136};
ram[17691] = {9'd68,-10'd132};
ram[17692] = {9'd71,-10'd129};
ram[17693] = {9'd74,-10'd126};
ram[17694] = {9'd77,-10'd123};
ram[17695] = {9'd80,-10'd120};
ram[17696] = {9'd84,-10'd117};
ram[17697] = {9'd87,-10'd114};
ram[17698] = {9'd90,-10'd110};
ram[17699] = {9'd93,-10'd107};
ram[17700] = {9'd96,-10'd104};
ram[17701] = {9'd99,-10'd101};
ram[17702] = {-9'd98,-10'd98};
ram[17703] = {-9'd95,-10'd95};
ram[17704] = {-9'd92,-10'd92};
ram[17705] = {-9'd88,-10'd88};
ram[17706] = {-9'd85,-10'd85};
ram[17707] = {-9'd82,-10'd82};
ram[17708] = {-9'd79,-10'd79};
ram[17709] = {-9'd76,-10'd76};
ram[17710] = {-9'd73,-10'd73};
ram[17711] = {-9'd70,-10'd70};
ram[17712] = {-9'd66,-10'd66};
ram[17713] = {-9'd63,-10'd63};
ram[17714] = {-9'd60,-10'd60};
ram[17715] = {-9'd57,-10'd57};
ram[17716] = {-9'd54,-10'd54};
ram[17717] = {-9'd51,-10'd51};
ram[17718] = {-9'd48,-10'd48};
ram[17719] = {-9'd44,-10'd44};
ram[17720] = {-9'd41,-10'd41};
ram[17721] = {-9'd38,-10'd38};
ram[17722] = {-9'd35,-10'd35};
ram[17723] = {-9'd32,-10'd32};
ram[17724] = {-9'd29,-10'd29};
ram[17725] = {-9'd26,-10'd26};
ram[17726] = {-9'd22,-10'd22};
ram[17727] = {-9'd19,-10'd19};
ram[17728] = {-9'd16,-10'd16};
ram[17729] = {-9'd13,-10'd13};
ram[17730] = {-9'd10,-10'd10};
ram[17731] = {-9'd7,-10'd7};
ram[17732] = {-9'd4,-10'd4};
ram[17733] = {9'd0,10'd0};
ram[17734] = {9'd3,10'd3};
ram[17735] = {9'd6,10'd6};
ram[17736] = {9'd9,10'd9};
ram[17737] = {9'd12,10'd12};
ram[17738] = {9'd15,10'd15};
ram[17739] = {9'd18,10'd18};
ram[17740] = {9'd21,10'd21};
ram[17741] = {9'd25,10'd25};
ram[17742] = {9'd28,10'd28};
ram[17743] = {9'd31,10'd31};
ram[17744] = {9'd34,10'd34};
ram[17745] = {9'd37,10'd37};
ram[17746] = {9'd40,10'd40};
ram[17747] = {9'd43,10'd43};
ram[17748] = {9'd47,10'd47};
ram[17749] = {9'd50,10'd50};
ram[17750] = {9'd53,10'd53};
ram[17751] = {9'd56,10'd56};
ram[17752] = {9'd59,10'd59};
ram[17753] = {9'd62,10'd62};
ram[17754] = {9'd65,10'd65};
ram[17755] = {9'd69,10'd69};
ram[17756] = {9'd72,10'd72};
ram[17757] = {9'd75,10'd75};
ram[17758] = {9'd78,10'd78};
ram[17759] = {9'd81,10'd81};
ram[17760] = {9'd84,10'd84};
ram[17761] = {9'd87,10'd87};
ram[17762] = {9'd91,10'd91};
ram[17763] = {9'd94,10'd94};
ram[17764] = {9'd97,10'd97};
ram[17765] = {-9'd100,10'd100};
ram[17766] = {-9'd97,10'd103};
ram[17767] = {-9'd94,10'd106};
ram[17768] = {-9'd91,10'd109};
ram[17769] = {-9'd88,10'd113};
ram[17770] = {-9'd85,10'd116};
ram[17771] = {-9'd81,10'd119};
ram[17772] = {-9'd78,10'd122};
ram[17773] = {-9'd75,10'd125};
ram[17774] = {-9'd72,10'd128};
ram[17775] = {-9'd69,10'd131};
ram[17776] = {-9'd66,10'd135};
ram[17777] = {-9'd63,10'd138};
ram[17778] = {-9'd59,10'd141};
ram[17779] = {-9'd56,10'd144};
ram[17780] = {-9'd53,10'd147};
ram[17781] = {-9'd50,10'd150};
ram[17782] = {-9'd47,10'd153};
ram[17783] = {-9'd44,10'd157};
ram[17784] = {-9'd41,10'd160};
ram[17785] = {-9'd37,10'd163};
ram[17786] = {-9'd34,10'd166};
ram[17787] = {-9'd31,10'd169};
ram[17788] = {-9'd28,10'd172};
ram[17789] = {-9'd25,10'd175};
ram[17790] = {-9'd22,10'd179};
ram[17791] = {-9'd19,10'd182};
ram[17792] = {-9'd19,10'd182};
ram[17793] = {-9'd15,10'd185};
ram[17794] = {-9'd12,10'd188};
ram[17795] = {-9'd9,10'd191};
ram[17796] = {-9'd6,10'd194};
ram[17797] = {-9'd3,10'd197};
ram[17798] = {9'd0,10'd201};
ram[17799] = {9'd3,10'd204};
ram[17800] = {9'd7,10'd207};
ram[17801] = {9'd10,10'd210};
ram[17802] = {9'd13,10'd213};
ram[17803] = {9'd16,10'd216};
ram[17804] = {9'd19,10'd219};
ram[17805] = {9'd22,10'd223};
ram[17806] = {9'd25,10'd226};
ram[17807] = {9'd29,10'd229};
ram[17808] = {9'd32,10'd232};
ram[17809] = {9'd35,10'd235};
ram[17810] = {9'd38,10'd238};
ram[17811] = {9'd41,10'd241};
ram[17812] = {9'd44,10'd245};
ram[17813] = {9'd47,10'd248};
ram[17814] = {9'd51,10'd251};
ram[17815] = {9'd54,10'd254};
ram[17816] = {9'd57,10'd257};
ram[17817] = {9'd60,10'd260};
ram[17818] = {9'd63,10'd263};
ram[17819] = {9'd66,10'd267};
ram[17820] = {9'd69,10'd270};
ram[17821] = {9'd73,10'd273};
ram[17822] = {9'd76,10'd276};
ram[17823] = {9'd79,10'd279};
ram[17824] = {9'd82,10'd282};
ram[17825] = {9'd85,10'd285};
ram[17826] = {9'd88,10'd289};
ram[17827] = {9'd91,10'd292};
ram[17828] = {9'd95,10'd295};
ram[17829] = {9'd98,10'd298};
ram[17830] = {-9'd99,10'd301};
ram[17831] = {-9'd96,10'd304};
ram[17832] = {-9'd93,10'd307};
ram[17833] = {-9'd90,10'd311};
ram[17834] = {-9'd87,10'd314};
ram[17835] = {-9'd84,10'd317};
ram[17836] = {-9'd81,10'd320};
ram[17837] = {-9'd77,10'd323};
ram[17838] = {-9'd74,10'd326};
ram[17839] = {-9'd71,10'd329};
ram[17840] = {-9'd68,10'd333};
ram[17841] = {-9'd65,10'd336};
ram[17842] = {-9'd62,10'd339};
ram[17843] = {-9'd59,10'd342};
ram[17844] = {-9'd55,10'd345};
ram[17845] = {-9'd52,10'd348};
ram[17846] = {-9'd49,10'd351};
ram[17847] = {-9'd46,10'd354};
ram[17848] = {-9'd43,10'd358};
ram[17849] = {-9'd40,10'd361};
ram[17850] = {-9'd37,10'd364};
ram[17851] = {-9'd33,10'd367};
ram[17852] = {-9'd30,10'd370};
ram[17853] = {-9'd27,10'd373};
ram[17854] = {-9'd24,10'd376};
ram[17855] = {-9'd21,10'd380};
ram[17856] = {-9'd18,10'd383};
ram[17857] = {-9'd15,10'd386};
ram[17858] = {-9'd11,10'd389};
ram[17859] = {-9'd8,10'd392};
ram[17860] = {-9'd5,10'd395};
ram[17861] = {-9'd2,10'd398};
ram[17862] = {9'd1,-10'd399};
ram[17863] = {9'd4,-10'd396};
ram[17864] = {9'd7,-10'd393};
ram[17865] = {9'd10,-10'd390};
ram[17866] = {9'd14,-10'd387};
ram[17867] = {9'd17,-10'd384};
ram[17868] = {9'd20,-10'd381};
ram[17869] = {9'd23,-10'd377};
ram[17870] = {9'd26,-10'd374};
ram[17871] = {9'd29,-10'd371};
ram[17872] = {9'd32,-10'd368};
ram[17873] = {9'd36,-10'd365};
ram[17874] = {9'd39,-10'd362};
ram[17875] = {9'd42,-10'd359};
ram[17876] = {9'd45,-10'd355};
ram[17877] = {9'd48,-10'd352};
ram[17878] = {9'd51,-10'd349};
ram[17879] = {9'd54,-10'd346};
ram[17880] = {9'd58,-10'd343};
ram[17881] = {9'd61,-10'd340};
ram[17882] = {9'd64,-10'd337};
ram[17883] = {9'd67,-10'd334};
ram[17884] = {9'd70,-10'd330};
ram[17885] = {9'd73,-10'd327};
ram[17886] = {9'd76,-10'd324};
ram[17887] = {9'd80,-10'd321};
ram[17888] = {9'd83,-10'd318};
ram[17889] = {9'd86,-10'd315};
ram[17890] = {9'd89,-10'd312};
ram[17891] = {9'd92,-10'd308};
ram[17892] = {9'd95,-10'd305};
ram[17893] = {9'd98,-10'd302};
ram[17894] = {-9'd99,-10'd299};
ram[17895] = {-9'd96,-10'd296};
ram[17896] = {-9'd92,-10'd293};
ram[17897] = {-9'd89,-10'd290};
ram[17898] = {-9'd86,-10'd286};
ram[17899] = {-9'd83,-10'd283};
ram[17900] = {-9'd80,-10'd280};
ram[17901] = {-9'd77,-10'd277};
ram[17902] = {-9'd74,-10'd274};
ram[17903] = {-9'd70,-10'd271};
ram[17904] = {-9'd67,-10'd268};
ram[17905] = {-9'd64,-10'd264};
ram[17906] = {-9'd61,-10'd261};
ram[17907] = {-9'd58,-10'd258};
ram[17908] = {-9'd55,-10'd255};
ram[17909] = {-9'd52,-10'd252};
ram[17910] = {-9'd48,-10'd249};
ram[17911] = {-9'd45,-10'd246};
ram[17912] = {-9'd42,-10'd242};
ram[17913] = {-9'd39,-10'd239};
ram[17914] = {-9'd36,-10'd236};
ram[17915] = {-9'd33,-10'd233};
ram[17916] = {-9'd30,-10'd230};
ram[17917] = {-9'd26,-10'd227};
ram[17918] = {-9'd23,-10'd224};
ram[17919] = {-9'd20,-10'd220};
ram[17920] = {-9'd20,-10'd220};
ram[17921] = {-9'd17,-10'd217};
ram[17922] = {-9'd14,-10'd214};
ram[17923] = {-9'd11,-10'd211};
ram[17924] = {-9'd8,-10'd208};
ram[17925] = {-9'd4,-10'd205};
ram[17926] = {-9'd1,-10'd202};
ram[17927] = {9'd2,-10'd198};
ram[17928] = {9'd5,-10'd195};
ram[17929] = {9'd8,-10'd192};
ram[17930] = {9'd11,-10'd189};
ram[17931] = {9'd14,-10'd186};
ram[17932] = {9'd18,-10'd183};
ram[17933] = {9'd21,-10'd180};
ram[17934] = {9'd24,-10'd176};
ram[17935] = {9'd27,-10'd173};
ram[17936] = {9'd30,-10'd170};
ram[17937] = {9'd33,-10'd167};
ram[17938] = {9'd36,-10'd164};
ram[17939] = {9'd40,-10'd161};
ram[17940] = {9'd43,-10'd158};
ram[17941] = {9'd46,-10'd154};
ram[17942] = {9'd49,-10'd151};
ram[17943] = {9'd52,-10'd148};
ram[17944] = {9'd55,-10'd145};
ram[17945] = {9'd58,-10'd142};
ram[17946] = {9'd62,-10'd139};
ram[17947] = {9'd65,-10'd136};
ram[17948] = {9'd68,-10'd132};
ram[17949] = {9'd71,-10'd129};
ram[17950] = {9'd74,-10'd126};
ram[17951] = {9'd77,-10'd123};
ram[17952] = {9'd80,-10'd120};
ram[17953] = {9'd84,-10'd117};
ram[17954] = {9'd87,-10'd114};
ram[17955] = {9'd90,-10'd110};
ram[17956] = {9'd93,-10'd107};
ram[17957] = {9'd96,-10'd104};
ram[17958] = {9'd99,-10'd101};
ram[17959] = {-9'd98,-10'd98};
ram[17960] = {-9'd95,-10'd95};
ram[17961] = {-9'd92,-10'd92};
ram[17962] = {-9'd88,-10'd88};
ram[17963] = {-9'd85,-10'd85};
ram[17964] = {-9'd82,-10'd82};
ram[17965] = {-9'd79,-10'd79};
ram[17966] = {-9'd76,-10'd76};
ram[17967] = {-9'd73,-10'd73};
ram[17968] = {-9'd70,-10'd70};
ram[17969] = {-9'd66,-10'd66};
ram[17970] = {-9'd63,-10'd63};
ram[17971] = {-9'd60,-10'd60};
ram[17972] = {-9'd57,-10'd57};
ram[17973] = {-9'd54,-10'd54};
ram[17974] = {-9'd51,-10'd51};
ram[17975] = {-9'd48,-10'd48};
ram[17976] = {-9'd44,-10'd44};
ram[17977] = {-9'd41,-10'd41};
ram[17978] = {-9'd38,-10'd38};
ram[17979] = {-9'd35,-10'd35};
ram[17980] = {-9'd32,-10'd32};
ram[17981] = {-9'd29,-10'd29};
ram[17982] = {-9'd26,-10'd26};
ram[17983] = {-9'd22,-10'd22};
ram[17984] = {-9'd19,-10'd19};
ram[17985] = {-9'd16,-10'd16};
ram[17986] = {-9'd13,-10'd13};
ram[17987] = {-9'd10,-10'd10};
ram[17988] = {-9'd7,-10'd7};
ram[17989] = {-9'd4,-10'd4};
ram[17990] = {9'd0,10'd0};
ram[17991] = {9'd3,10'd3};
ram[17992] = {9'd6,10'd6};
ram[17993] = {9'd9,10'd9};
ram[17994] = {9'd12,10'd12};
ram[17995] = {9'd15,10'd15};
ram[17996] = {9'd18,10'd18};
ram[17997] = {9'd21,10'd21};
ram[17998] = {9'd25,10'd25};
ram[17999] = {9'd28,10'd28};
ram[18000] = {9'd31,10'd31};
ram[18001] = {9'd34,10'd34};
ram[18002] = {9'd37,10'd37};
ram[18003] = {9'd40,10'd40};
ram[18004] = {9'd43,10'd43};
ram[18005] = {9'd47,10'd47};
ram[18006] = {9'd50,10'd50};
ram[18007] = {9'd53,10'd53};
ram[18008] = {9'd56,10'd56};
ram[18009] = {9'd59,10'd59};
ram[18010] = {9'd62,10'd62};
ram[18011] = {9'd65,10'd65};
ram[18012] = {9'd69,10'd69};
ram[18013] = {9'd72,10'd72};
ram[18014] = {9'd75,10'd75};
ram[18015] = {9'd78,10'd78};
ram[18016] = {9'd81,10'd81};
ram[18017] = {9'd84,10'd84};
ram[18018] = {9'd87,10'd87};
ram[18019] = {9'd91,10'd91};
ram[18020] = {9'd94,10'd94};
ram[18021] = {9'd97,10'd97};
ram[18022] = {-9'd100,10'd100};
ram[18023] = {-9'd97,10'd103};
ram[18024] = {-9'd94,10'd106};
ram[18025] = {-9'd91,10'd109};
ram[18026] = {-9'd88,10'd113};
ram[18027] = {-9'd85,10'd116};
ram[18028] = {-9'd81,10'd119};
ram[18029] = {-9'd78,10'd122};
ram[18030] = {-9'd75,10'd125};
ram[18031] = {-9'd72,10'd128};
ram[18032] = {-9'd69,10'd131};
ram[18033] = {-9'd66,10'd135};
ram[18034] = {-9'd63,10'd138};
ram[18035] = {-9'd59,10'd141};
ram[18036] = {-9'd56,10'd144};
ram[18037] = {-9'd53,10'd147};
ram[18038] = {-9'd50,10'd150};
ram[18039] = {-9'd47,10'd153};
ram[18040] = {-9'd44,10'd157};
ram[18041] = {-9'd41,10'd160};
ram[18042] = {-9'd37,10'd163};
ram[18043] = {-9'd34,10'd166};
ram[18044] = {-9'd31,10'd169};
ram[18045] = {-9'd28,10'd172};
ram[18046] = {-9'd25,10'd175};
ram[18047] = {-9'd22,10'd179};
ram[18048] = {-9'd22,10'd179};
ram[18049] = {-9'd19,10'd182};
ram[18050] = {-9'd15,10'd185};
ram[18051] = {-9'd12,10'd188};
ram[18052] = {-9'd9,10'd191};
ram[18053] = {-9'd6,10'd194};
ram[18054] = {-9'd3,10'd197};
ram[18055] = {9'd0,10'd201};
ram[18056] = {9'd3,10'd204};
ram[18057] = {9'd7,10'd207};
ram[18058] = {9'd10,10'd210};
ram[18059] = {9'd13,10'd213};
ram[18060] = {9'd16,10'd216};
ram[18061] = {9'd19,10'd219};
ram[18062] = {9'd22,10'd223};
ram[18063] = {9'd25,10'd226};
ram[18064] = {9'd29,10'd229};
ram[18065] = {9'd32,10'd232};
ram[18066] = {9'd35,10'd235};
ram[18067] = {9'd38,10'd238};
ram[18068] = {9'd41,10'd241};
ram[18069] = {9'd44,10'd245};
ram[18070] = {9'd47,10'd248};
ram[18071] = {9'd51,10'd251};
ram[18072] = {9'd54,10'd254};
ram[18073] = {9'd57,10'd257};
ram[18074] = {9'd60,10'd260};
ram[18075] = {9'd63,10'd263};
ram[18076] = {9'd66,10'd267};
ram[18077] = {9'd69,10'd270};
ram[18078] = {9'd73,10'd273};
ram[18079] = {9'd76,10'd276};
ram[18080] = {9'd79,10'd279};
ram[18081] = {9'd82,10'd282};
ram[18082] = {9'd85,10'd285};
ram[18083] = {9'd88,10'd289};
ram[18084] = {9'd91,10'd292};
ram[18085] = {9'd95,10'd295};
ram[18086] = {9'd98,10'd298};
ram[18087] = {-9'd99,10'd301};
ram[18088] = {-9'd96,10'd304};
ram[18089] = {-9'd93,10'd307};
ram[18090] = {-9'd90,10'd311};
ram[18091] = {-9'd87,10'd314};
ram[18092] = {-9'd84,10'd317};
ram[18093] = {-9'd81,10'd320};
ram[18094] = {-9'd77,10'd323};
ram[18095] = {-9'd74,10'd326};
ram[18096] = {-9'd71,10'd329};
ram[18097] = {-9'd68,10'd333};
ram[18098] = {-9'd65,10'd336};
ram[18099] = {-9'd62,10'd339};
ram[18100] = {-9'd59,10'd342};
ram[18101] = {-9'd55,10'd345};
ram[18102] = {-9'd52,10'd348};
ram[18103] = {-9'd49,10'd351};
ram[18104] = {-9'd46,10'd354};
ram[18105] = {-9'd43,10'd358};
ram[18106] = {-9'd40,10'd361};
ram[18107] = {-9'd37,10'd364};
ram[18108] = {-9'd33,10'd367};
ram[18109] = {-9'd30,10'd370};
ram[18110] = {-9'd27,10'd373};
ram[18111] = {-9'd24,10'd376};
ram[18112] = {-9'd21,10'd380};
ram[18113] = {-9'd18,10'd383};
ram[18114] = {-9'd15,10'd386};
ram[18115] = {-9'd11,10'd389};
ram[18116] = {-9'd8,10'd392};
ram[18117] = {-9'd5,10'd395};
ram[18118] = {-9'd2,10'd398};
ram[18119] = {9'd1,-10'd399};
ram[18120] = {9'd4,-10'd396};
ram[18121] = {9'd7,-10'd393};
ram[18122] = {9'd10,-10'd390};
ram[18123] = {9'd14,-10'd387};
ram[18124] = {9'd17,-10'd384};
ram[18125] = {9'd20,-10'd381};
ram[18126] = {9'd23,-10'd377};
ram[18127] = {9'd26,-10'd374};
ram[18128] = {9'd29,-10'd371};
ram[18129] = {9'd32,-10'd368};
ram[18130] = {9'd36,-10'd365};
ram[18131] = {9'd39,-10'd362};
ram[18132] = {9'd42,-10'd359};
ram[18133] = {9'd45,-10'd355};
ram[18134] = {9'd48,-10'd352};
ram[18135] = {9'd51,-10'd349};
ram[18136] = {9'd54,-10'd346};
ram[18137] = {9'd58,-10'd343};
ram[18138] = {9'd61,-10'd340};
ram[18139] = {9'd64,-10'd337};
ram[18140] = {9'd67,-10'd334};
ram[18141] = {9'd70,-10'd330};
ram[18142] = {9'd73,-10'd327};
ram[18143] = {9'd76,-10'd324};
ram[18144] = {9'd80,-10'd321};
ram[18145] = {9'd83,-10'd318};
ram[18146] = {9'd86,-10'd315};
ram[18147] = {9'd89,-10'd312};
ram[18148] = {9'd92,-10'd308};
ram[18149] = {9'd95,-10'd305};
ram[18150] = {9'd98,-10'd302};
ram[18151] = {-9'd99,-10'd299};
ram[18152] = {-9'd96,-10'd296};
ram[18153] = {-9'd92,-10'd293};
ram[18154] = {-9'd89,-10'd290};
ram[18155] = {-9'd86,-10'd286};
ram[18156] = {-9'd83,-10'd283};
ram[18157] = {-9'd80,-10'd280};
ram[18158] = {-9'd77,-10'd277};
ram[18159] = {-9'd74,-10'd274};
ram[18160] = {-9'd70,-10'd271};
ram[18161] = {-9'd67,-10'd268};
ram[18162] = {-9'd64,-10'd264};
ram[18163] = {-9'd61,-10'd261};
ram[18164] = {-9'd58,-10'd258};
ram[18165] = {-9'd55,-10'd255};
ram[18166] = {-9'd52,-10'd252};
ram[18167] = {-9'd48,-10'd249};
ram[18168] = {-9'd45,-10'd246};
ram[18169] = {-9'd42,-10'd242};
ram[18170] = {-9'd39,-10'd239};
ram[18171] = {-9'd36,-10'd236};
ram[18172] = {-9'd33,-10'd233};
ram[18173] = {-9'd30,-10'd230};
ram[18174] = {-9'd26,-10'd227};
ram[18175] = {-9'd23,-10'd224};
ram[18176] = {-9'd23,-10'd224};
ram[18177] = {-9'd20,-10'd220};
ram[18178] = {-9'd17,-10'd217};
ram[18179] = {-9'd14,-10'd214};
ram[18180] = {-9'd11,-10'd211};
ram[18181] = {-9'd8,-10'd208};
ram[18182] = {-9'd4,-10'd205};
ram[18183] = {-9'd1,-10'd202};
ram[18184] = {9'd2,-10'd198};
ram[18185] = {9'd5,-10'd195};
ram[18186] = {9'd8,-10'd192};
ram[18187] = {9'd11,-10'd189};
ram[18188] = {9'd14,-10'd186};
ram[18189] = {9'd18,-10'd183};
ram[18190] = {9'd21,-10'd180};
ram[18191] = {9'd24,-10'd176};
ram[18192] = {9'd27,-10'd173};
ram[18193] = {9'd30,-10'd170};
ram[18194] = {9'd33,-10'd167};
ram[18195] = {9'd36,-10'd164};
ram[18196] = {9'd40,-10'd161};
ram[18197] = {9'd43,-10'd158};
ram[18198] = {9'd46,-10'd154};
ram[18199] = {9'd49,-10'd151};
ram[18200] = {9'd52,-10'd148};
ram[18201] = {9'd55,-10'd145};
ram[18202] = {9'd58,-10'd142};
ram[18203] = {9'd62,-10'd139};
ram[18204] = {9'd65,-10'd136};
ram[18205] = {9'd68,-10'd132};
ram[18206] = {9'd71,-10'd129};
ram[18207] = {9'd74,-10'd126};
ram[18208] = {9'd77,-10'd123};
ram[18209] = {9'd80,-10'd120};
ram[18210] = {9'd84,-10'd117};
ram[18211] = {9'd87,-10'd114};
ram[18212] = {9'd90,-10'd110};
ram[18213] = {9'd93,-10'd107};
ram[18214] = {9'd96,-10'd104};
ram[18215] = {9'd99,-10'd101};
ram[18216] = {-9'd98,-10'd98};
ram[18217] = {-9'd95,-10'd95};
ram[18218] = {-9'd92,-10'd92};
ram[18219] = {-9'd88,-10'd88};
ram[18220] = {-9'd85,-10'd85};
ram[18221] = {-9'd82,-10'd82};
ram[18222] = {-9'd79,-10'd79};
ram[18223] = {-9'd76,-10'd76};
ram[18224] = {-9'd73,-10'd73};
ram[18225] = {-9'd70,-10'd70};
ram[18226] = {-9'd66,-10'd66};
ram[18227] = {-9'd63,-10'd63};
ram[18228] = {-9'd60,-10'd60};
ram[18229] = {-9'd57,-10'd57};
ram[18230] = {-9'd54,-10'd54};
ram[18231] = {-9'd51,-10'd51};
ram[18232] = {-9'd48,-10'd48};
ram[18233] = {-9'd44,-10'd44};
ram[18234] = {-9'd41,-10'd41};
ram[18235] = {-9'd38,-10'd38};
ram[18236] = {-9'd35,-10'd35};
ram[18237] = {-9'd32,-10'd32};
ram[18238] = {-9'd29,-10'd29};
ram[18239] = {-9'd26,-10'd26};
ram[18240] = {-9'd22,-10'd22};
ram[18241] = {-9'd19,-10'd19};
ram[18242] = {-9'd16,-10'd16};
ram[18243] = {-9'd13,-10'd13};
ram[18244] = {-9'd10,-10'd10};
ram[18245] = {-9'd7,-10'd7};
ram[18246] = {-9'd4,-10'd4};
ram[18247] = {9'd0,10'd0};
ram[18248] = {9'd3,10'd3};
ram[18249] = {9'd6,10'd6};
ram[18250] = {9'd9,10'd9};
ram[18251] = {9'd12,10'd12};
ram[18252] = {9'd15,10'd15};
ram[18253] = {9'd18,10'd18};
ram[18254] = {9'd21,10'd21};
ram[18255] = {9'd25,10'd25};
ram[18256] = {9'd28,10'd28};
ram[18257] = {9'd31,10'd31};
ram[18258] = {9'd34,10'd34};
ram[18259] = {9'd37,10'd37};
ram[18260] = {9'd40,10'd40};
ram[18261] = {9'd43,10'd43};
ram[18262] = {9'd47,10'd47};
ram[18263] = {9'd50,10'd50};
ram[18264] = {9'd53,10'd53};
ram[18265] = {9'd56,10'd56};
ram[18266] = {9'd59,10'd59};
ram[18267] = {9'd62,10'd62};
ram[18268] = {9'd65,10'd65};
ram[18269] = {9'd69,10'd69};
ram[18270] = {9'd72,10'd72};
ram[18271] = {9'd75,10'd75};
ram[18272] = {9'd78,10'd78};
ram[18273] = {9'd81,10'd81};
ram[18274] = {9'd84,10'd84};
ram[18275] = {9'd87,10'd87};
ram[18276] = {9'd91,10'd91};
ram[18277] = {9'd94,10'd94};
ram[18278] = {9'd97,10'd97};
ram[18279] = {-9'd100,10'd100};
ram[18280] = {-9'd97,10'd103};
ram[18281] = {-9'd94,10'd106};
ram[18282] = {-9'd91,10'd109};
ram[18283] = {-9'd88,10'd113};
ram[18284] = {-9'd85,10'd116};
ram[18285] = {-9'd81,10'd119};
ram[18286] = {-9'd78,10'd122};
ram[18287] = {-9'd75,10'd125};
ram[18288] = {-9'd72,10'd128};
ram[18289] = {-9'd69,10'd131};
ram[18290] = {-9'd66,10'd135};
ram[18291] = {-9'd63,10'd138};
ram[18292] = {-9'd59,10'd141};
ram[18293] = {-9'd56,10'd144};
ram[18294] = {-9'd53,10'd147};
ram[18295] = {-9'd50,10'd150};
ram[18296] = {-9'd47,10'd153};
ram[18297] = {-9'd44,10'd157};
ram[18298] = {-9'd41,10'd160};
ram[18299] = {-9'd37,10'd163};
ram[18300] = {-9'd34,10'd166};
ram[18301] = {-9'd31,10'd169};
ram[18302] = {-9'd28,10'd172};
ram[18303] = {-9'd25,10'd175};
ram[18304] = {-9'd25,10'd175};
ram[18305] = {-9'd22,10'd179};
ram[18306] = {-9'd19,10'd182};
ram[18307] = {-9'd15,10'd185};
ram[18308] = {-9'd12,10'd188};
ram[18309] = {-9'd9,10'd191};
ram[18310] = {-9'd6,10'd194};
ram[18311] = {-9'd3,10'd197};
ram[18312] = {9'd0,10'd201};
ram[18313] = {9'd3,10'd204};
ram[18314] = {9'd7,10'd207};
ram[18315] = {9'd10,10'd210};
ram[18316] = {9'd13,10'd213};
ram[18317] = {9'd16,10'd216};
ram[18318] = {9'd19,10'd219};
ram[18319] = {9'd22,10'd223};
ram[18320] = {9'd25,10'd226};
ram[18321] = {9'd29,10'd229};
ram[18322] = {9'd32,10'd232};
ram[18323] = {9'd35,10'd235};
ram[18324] = {9'd38,10'd238};
ram[18325] = {9'd41,10'd241};
ram[18326] = {9'd44,10'd245};
ram[18327] = {9'd47,10'd248};
ram[18328] = {9'd51,10'd251};
ram[18329] = {9'd54,10'd254};
ram[18330] = {9'd57,10'd257};
ram[18331] = {9'd60,10'd260};
ram[18332] = {9'd63,10'd263};
ram[18333] = {9'd66,10'd267};
ram[18334] = {9'd69,10'd270};
ram[18335] = {9'd73,10'd273};
ram[18336] = {9'd76,10'd276};
ram[18337] = {9'd79,10'd279};
ram[18338] = {9'd82,10'd282};
ram[18339] = {9'd85,10'd285};
ram[18340] = {9'd88,10'd289};
ram[18341] = {9'd91,10'd292};
ram[18342] = {9'd95,10'd295};
ram[18343] = {9'd98,10'd298};
ram[18344] = {-9'd99,10'd301};
ram[18345] = {-9'd96,10'd304};
ram[18346] = {-9'd93,10'd307};
ram[18347] = {-9'd90,10'd311};
ram[18348] = {-9'd87,10'd314};
ram[18349] = {-9'd84,10'd317};
ram[18350] = {-9'd81,10'd320};
ram[18351] = {-9'd77,10'd323};
ram[18352] = {-9'd74,10'd326};
ram[18353] = {-9'd71,10'd329};
ram[18354] = {-9'd68,10'd333};
ram[18355] = {-9'd65,10'd336};
ram[18356] = {-9'd62,10'd339};
ram[18357] = {-9'd59,10'd342};
ram[18358] = {-9'd55,10'd345};
ram[18359] = {-9'd52,10'd348};
ram[18360] = {-9'd49,10'd351};
ram[18361] = {-9'd46,10'd354};
ram[18362] = {-9'd43,10'd358};
ram[18363] = {-9'd40,10'd361};
ram[18364] = {-9'd37,10'd364};
ram[18365] = {-9'd33,10'd367};
ram[18366] = {-9'd30,10'd370};
ram[18367] = {-9'd27,10'd373};
ram[18368] = {-9'd24,10'd376};
ram[18369] = {-9'd21,10'd380};
ram[18370] = {-9'd18,10'd383};
ram[18371] = {-9'd15,10'd386};
ram[18372] = {-9'd11,10'd389};
ram[18373] = {-9'd8,10'd392};
ram[18374] = {-9'd5,10'd395};
ram[18375] = {-9'd2,10'd398};
ram[18376] = {9'd1,-10'd399};
ram[18377] = {9'd4,-10'd396};
ram[18378] = {9'd7,-10'd393};
ram[18379] = {9'd10,-10'd390};
ram[18380] = {9'd14,-10'd387};
ram[18381] = {9'd17,-10'd384};
ram[18382] = {9'd20,-10'd381};
ram[18383] = {9'd23,-10'd377};
ram[18384] = {9'd26,-10'd374};
ram[18385] = {9'd29,-10'd371};
ram[18386] = {9'd32,-10'd368};
ram[18387] = {9'd36,-10'd365};
ram[18388] = {9'd39,-10'd362};
ram[18389] = {9'd42,-10'd359};
ram[18390] = {9'd45,-10'd355};
ram[18391] = {9'd48,-10'd352};
ram[18392] = {9'd51,-10'd349};
ram[18393] = {9'd54,-10'd346};
ram[18394] = {9'd58,-10'd343};
ram[18395] = {9'd61,-10'd340};
ram[18396] = {9'd64,-10'd337};
ram[18397] = {9'd67,-10'd334};
ram[18398] = {9'd70,-10'd330};
ram[18399] = {9'd73,-10'd327};
ram[18400] = {9'd76,-10'd324};
ram[18401] = {9'd80,-10'd321};
ram[18402] = {9'd83,-10'd318};
ram[18403] = {9'd86,-10'd315};
ram[18404] = {9'd89,-10'd312};
ram[18405] = {9'd92,-10'd308};
ram[18406] = {9'd95,-10'd305};
ram[18407] = {9'd98,-10'd302};
ram[18408] = {-9'd99,-10'd299};
ram[18409] = {-9'd96,-10'd296};
ram[18410] = {-9'd92,-10'd293};
ram[18411] = {-9'd89,-10'd290};
ram[18412] = {-9'd86,-10'd286};
ram[18413] = {-9'd83,-10'd283};
ram[18414] = {-9'd80,-10'd280};
ram[18415] = {-9'd77,-10'd277};
ram[18416] = {-9'd74,-10'd274};
ram[18417] = {-9'd70,-10'd271};
ram[18418] = {-9'd67,-10'd268};
ram[18419] = {-9'd64,-10'd264};
ram[18420] = {-9'd61,-10'd261};
ram[18421] = {-9'd58,-10'd258};
ram[18422] = {-9'd55,-10'd255};
ram[18423] = {-9'd52,-10'd252};
ram[18424] = {-9'd48,-10'd249};
ram[18425] = {-9'd45,-10'd246};
ram[18426] = {-9'd42,-10'd242};
ram[18427] = {-9'd39,-10'd239};
ram[18428] = {-9'd36,-10'd236};
ram[18429] = {-9'd33,-10'd233};
ram[18430] = {-9'd30,-10'd230};
ram[18431] = {-9'd26,-10'd227};
ram[18432] = {-9'd26,-10'd227};
ram[18433] = {-9'd23,-10'd224};
ram[18434] = {-9'd20,-10'd220};
ram[18435] = {-9'd17,-10'd217};
ram[18436] = {-9'd14,-10'd214};
ram[18437] = {-9'd11,-10'd211};
ram[18438] = {-9'd8,-10'd208};
ram[18439] = {-9'd4,-10'd205};
ram[18440] = {-9'd1,-10'd202};
ram[18441] = {9'd2,-10'd198};
ram[18442] = {9'd5,-10'd195};
ram[18443] = {9'd8,-10'd192};
ram[18444] = {9'd11,-10'd189};
ram[18445] = {9'd14,-10'd186};
ram[18446] = {9'd18,-10'd183};
ram[18447] = {9'd21,-10'd180};
ram[18448] = {9'd24,-10'd176};
ram[18449] = {9'd27,-10'd173};
ram[18450] = {9'd30,-10'd170};
ram[18451] = {9'd33,-10'd167};
ram[18452] = {9'd36,-10'd164};
ram[18453] = {9'd40,-10'd161};
ram[18454] = {9'd43,-10'd158};
ram[18455] = {9'd46,-10'd154};
ram[18456] = {9'd49,-10'd151};
ram[18457] = {9'd52,-10'd148};
ram[18458] = {9'd55,-10'd145};
ram[18459] = {9'd58,-10'd142};
ram[18460] = {9'd62,-10'd139};
ram[18461] = {9'd65,-10'd136};
ram[18462] = {9'd68,-10'd132};
ram[18463] = {9'd71,-10'd129};
ram[18464] = {9'd74,-10'd126};
ram[18465] = {9'd77,-10'd123};
ram[18466] = {9'd80,-10'd120};
ram[18467] = {9'd84,-10'd117};
ram[18468] = {9'd87,-10'd114};
ram[18469] = {9'd90,-10'd110};
ram[18470] = {9'd93,-10'd107};
ram[18471] = {9'd96,-10'd104};
ram[18472] = {9'd99,-10'd101};
ram[18473] = {-9'd98,-10'd98};
ram[18474] = {-9'd95,-10'd95};
ram[18475] = {-9'd92,-10'd92};
ram[18476] = {-9'd88,-10'd88};
ram[18477] = {-9'd85,-10'd85};
ram[18478] = {-9'd82,-10'd82};
ram[18479] = {-9'd79,-10'd79};
ram[18480] = {-9'd76,-10'd76};
ram[18481] = {-9'd73,-10'd73};
ram[18482] = {-9'd70,-10'd70};
ram[18483] = {-9'd66,-10'd66};
ram[18484] = {-9'd63,-10'd63};
ram[18485] = {-9'd60,-10'd60};
ram[18486] = {-9'd57,-10'd57};
ram[18487] = {-9'd54,-10'd54};
ram[18488] = {-9'd51,-10'd51};
ram[18489] = {-9'd48,-10'd48};
ram[18490] = {-9'd44,-10'd44};
ram[18491] = {-9'd41,-10'd41};
ram[18492] = {-9'd38,-10'd38};
ram[18493] = {-9'd35,-10'd35};
ram[18494] = {-9'd32,-10'd32};
ram[18495] = {-9'd29,-10'd29};
ram[18496] = {-9'd26,-10'd26};
ram[18497] = {-9'd22,-10'd22};
ram[18498] = {-9'd19,-10'd19};
ram[18499] = {-9'd16,-10'd16};
ram[18500] = {-9'd13,-10'd13};
ram[18501] = {-9'd10,-10'd10};
ram[18502] = {-9'd7,-10'd7};
ram[18503] = {-9'd4,-10'd4};
ram[18504] = {9'd0,10'd0};
ram[18505] = {9'd3,10'd3};
ram[18506] = {9'd6,10'd6};
ram[18507] = {9'd9,10'd9};
ram[18508] = {9'd12,10'd12};
ram[18509] = {9'd15,10'd15};
ram[18510] = {9'd18,10'd18};
ram[18511] = {9'd21,10'd21};
ram[18512] = {9'd25,10'd25};
ram[18513] = {9'd28,10'd28};
ram[18514] = {9'd31,10'd31};
ram[18515] = {9'd34,10'd34};
ram[18516] = {9'd37,10'd37};
ram[18517] = {9'd40,10'd40};
ram[18518] = {9'd43,10'd43};
ram[18519] = {9'd47,10'd47};
ram[18520] = {9'd50,10'd50};
ram[18521] = {9'd53,10'd53};
ram[18522] = {9'd56,10'd56};
ram[18523] = {9'd59,10'd59};
ram[18524] = {9'd62,10'd62};
ram[18525] = {9'd65,10'd65};
ram[18526] = {9'd69,10'd69};
ram[18527] = {9'd72,10'd72};
ram[18528] = {9'd75,10'd75};
ram[18529] = {9'd78,10'd78};
ram[18530] = {9'd81,10'd81};
ram[18531] = {9'd84,10'd84};
ram[18532] = {9'd87,10'd87};
ram[18533] = {9'd91,10'd91};
ram[18534] = {9'd94,10'd94};
ram[18535] = {9'd97,10'd97};
ram[18536] = {-9'd100,10'd100};
ram[18537] = {-9'd97,10'd103};
ram[18538] = {-9'd94,10'd106};
ram[18539] = {-9'd91,10'd109};
ram[18540] = {-9'd88,10'd113};
ram[18541] = {-9'd85,10'd116};
ram[18542] = {-9'd81,10'd119};
ram[18543] = {-9'd78,10'd122};
ram[18544] = {-9'd75,10'd125};
ram[18545] = {-9'd72,10'd128};
ram[18546] = {-9'd69,10'd131};
ram[18547] = {-9'd66,10'd135};
ram[18548] = {-9'd63,10'd138};
ram[18549] = {-9'd59,10'd141};
ram[18550] = {-9'd56,10'd144};
ram[18551] = {-9'd53,10'd147};
ram[18552] = {-9'd50,10'd150};
ram[18553] = {-9'd47,10'd153};
ram[18554] = {-9'd44,10'd157};
ram[18555] = {-9'd41,10'd160};
ram[18556] = {-9'd37,10'd163};
ram[18557] = {-9'd34,10'd166};
ram[18558] = {-9'd31,10'd169};
ram[18559] = {-9'd28,10'd172};
ram[18560] = {-9'd28,10'd172};
ram[18561] = {-9'd25,10'd175};
ram[18562] = {-9'd22,10'd179};
ram[18563] = {-9'd19,10'd182};
ram[18564] = {-9'd15,10'd185};
ram[18565] = {-9'd12,10'd188};
ram[18566] = {-9'd9,10'd191};
ram[18567] = {-9'd6,10'd194};
ram[18568] = {-9'd3,10'd197};
ram[18569] = {9'd0,10'd201};
ram[18570] = {9'd3,10'd204};
ram[18571] = {9'd7,10'd207};
ram[18572] = {9'd10,10'd210};
ram[18573] = {9'd13,10'd213};
ram[18574] = {9'd16,10'd216};
ram[18575] = {9'd19,10'd219};
ram[18576] = {9'd22,10'd223};
ram[18577] = {9'd25,10'd226};
ram[18578] = {9'd29,10'd229};
ram[18579] = {9'd32,10'd232};
ram[18580] = {9'd35,10'd235};
ram[18581] = {9'd38,10'd238};
ram[18582] = {9'd41,10'd241};
ram[18583] = {9'd44,10'd245};
ram[18584] = {9'd47,10'd248};
ram[18585] = {9'd51,10'd251};
ram[18586] = {9'd54,10'd254};
ram[18587] = {9'd57,10'd257};
ram[18588] = {9'd60,10'd260};
ram[18589] = {9'd63,10'd263};
ram[18590] = {9'd66,10'd267};
ram[18591] = {9'd69,10'd270};
ram[18592] = {9'd73,10'd273};
ram[18593] = {9'd76,10'd276};
ram[18594] = {9'd79,10'd279};
ram[18595] = {9'd82,10'd282};
ram[18596] = {9'd85,10'd285};
ram[18597] = {9'd88,10'd289};
ram[18598] = {9'd91,10'd292};
ram[18599] = {9'd95,10'd295};
ram[18600] = {9'd98,10'd298};
ram[18601] = {-9'd99,10'd301};
ram[18602] = {-9'd96,10'd304};
ram[18603] = {-9'd93,10'd307};
ram[18604] = {-9'd90,10'd311};
ram[18605] = {-9'd87,10'd314};
ram[18606] = {-9'd84,10'd317};
ram[18607] = {-9'd81,10'd320};
ram[18608] = {-9'd77,10'd323};
ram[18609] = {-9'd74,10'd326};
ram[18610] = {-9'd71,10'd329};
ram[18611] = {-9'd68,10'd333};
ram[18612] = {-9'd65,10'd336};
ram[18613] = {-9'd62,10'd339};
ram[18614] = {-9'd59,10'd342};
ram[18615] = {-9'd55,10'd345};
ram[18616] = {-9'd52,10'd348};
ram[18617] = {-9'd49,10'd351};
ram[18618] = {-9'd46,10'd354};
ram[18619] = {-9'd43,10'd358};
ram[18620] = {-9'd40,10'd361};
ram[18621] = {-9'd37,10'd364};
ram[18622] = {-9'd33,10'd367};
ram[18623] = {-9'd30,10'd370};
ram[18624] = {-9'd27,10'd373};
ram[18625] = {-9'd24,10'd376};
ram[18626] = {-9'd21,10'd380};
ram[18627] = {-9'd18,10'd383};
ram[18628] = {-9'd15,10'd386};
ram[18629] = {-9'd11,10'd389};
ram[18630] = {-9'd8,10'd392};
ram[18631] = {-9'd5,10'd395};
ram[18632] = {-9'd2,10'd398};
ram[18633] = {9'd1,-10'd399};
ram[18634] = {9'd4,-10'd396};
ram[18635] = {9'd7,-10'd393};
ram[18636] = {9'd10,-10'd390};
ram[18637] = {9'd14,-10'd387};
ram[18638] = {9'd17,-10'd384};
ram[18639] = {9'd20,-10'd381};
ram[18640] = {9'd23,-10'd377};
ram[18641] = {9'd26,-10'd374};
ram[18642] = {9'd29,-10'd371};
ram[18643] = {9'd32,-10'd368};
ram[18644] = {9'd36,-10'd365};
ram[18645] = {9'd39,-10'd362};
ram[18646] = {9'd42,-10'd359};
ram[18647] = {9'd45,-10'd355};
ram[18648] = {9'd48,-10'd352};
ram[18649] = {9'd51,-10'd349};
ram[18650] = {9'd54,-10'd346};
ram[18651] = {9'd58,-10'd343};
ram[18652] = {9'd61,-10'd340};
ram[18653] = {9'd64,-10'd337};
ram[18654] = {9'd67,-10'd334};
ram[18655] = {9'd70,-10'd330};
ram[18656] = {9'd73,-10'd327};
ram[18657] = {9'd76,-10'd324};
ram[18658] = {9'd80,-10'd321};
ram[18659] = {9'd83,-10'd318};
ram[18660] = {9'd86,-10'd315};
ram[18661] = {9'd89,-10'd312};
ram[18662] = {9'd92,-10'd308};
ram[18663] = {9'd95,-10'd305};
ram[18664] = {9'd98,-10'd302};
ram[18665] = {-9'd99,-10'd299};
ram[18666] = {-9'd96,-10'd296};
ram[18667] = {-9'd92,-10'd293};
ram[18668] = {-9'd89,-10'd290};
ram[18669] = {-9'd86,-10'd286};
ram[18670] = {-9'd83,-10'd283};
ram[18671] = {-9'd80,-10'd280};
ram[18672] = {-9'd77,-10'd277};
ram[18673] = {-9'd74,-10'd274};
ram[18674] = {-9'd70,-10'd271};
ram[18675] = {-9'd67,-10'd268};
ram[18676] = {-9'd64,-10'd264};
ram[18677] = {-9'd61,-10'd261};
ram[18678] = {-9'd58,-10'd258};
ram[18679] = {-9'd55,-10'd255};
ram[18680] = {-9'd52,-10'd252};
ram[18681] = {-9'd48,-10'd249};
ram[18682] = {-9'd45,-10'd246};
ram[18683] = {-9'd42,-10'd242};
ram[18684] = {-9'd39,-10'd239};
ram[18685] = {-9'd36,-10'd236};
ram[18686] = {-9'd33,-10'd233};
ram[18687] = {-9'd30,-10'd230};
ram[18688] = {-9'd30,-10'd230};
ram[18689] = {-9'd26,-10'd227};
ram[18690] = {-9'd23,-10'd224};
ram[18691] = {-9'd20,-10'd220};
ram[18692] = {-9'd17,-10'd217};
ram[18693] = {-9'd14,-10'd214};
ram[18694] = {-9'd11,-10'd211};
ram[18695] = {-9'd8,-10'd208};
ram[18696] = {-9'd4,-10'd205};
ram[18697] = {-9'd1,-10'd202};
ram[18698] = {9'd2,-10'd198};
ram[18699] = {9'd5,-10'd195};
ram[18700] = {9'd8,-10'd192};
ram[18701] = {9'd11,-10'd189};
ram[18702] = {9'd14,-10'd186};
ram[18703] = {9'd18,-10'd183};
ram[18704] = {9'd21,-10'd180};
ram[18705] = {9'd24,-10'd176};
ram[18706] = {9'd27,-10'd173};
ram[18707] = {9'd30,-10'd170};
ram[18708] = {9'd33,-10'd167};
ram[18709] = {9'd36,-10'd164};
ram[18710] = {9'd40,-10'd161};
ram[18711] = {9'd43,-10'd158};
ram[18712] = {9'd46,-10'd154};
ram[18713] = {9'd49,-10'd151};
ram[18714] = {9'd52,-10'd148};
ram[18715] = {9'd55,-10'd145};
ram[18716] = {9'd58,-10'd142};
ram[18717] = {9'd62,-10'd139};
ram[18718] = {9'd65,-10'd136};
ram[18719] = {9'd68,-10'd132};
ram[18720] = {9'd71,-10'd129};
ram[18721] = {9'd74,-10'd126};
ram[18722] = {9'd77,-10'd123};
ram[18723] = {9'd80,-10'd120};
ram[18724] = {9'd84,-10'd117};
ram[18725] = {9'd87,-10'd114};
ram[18726] = {9'd90,-10'd110};
ram[18727] = {9'd93,-10'd107};
ram[18728] = {9'd96,-10'd104};
ram[18729] = {9'd99,-10'd101};
ram[18730] = {-9'd98,-10'd98};
ram[18731] = {-9'd95,-10'd95};
ram[18732] = {-9'd92,-10'd92};
ram[18733] = {-9'd88,-10'd88};
ram[18734] = {-9'd85,-10'd85};
ram[18735] = {-9'd82,-10'd82};
ram[18736] = {-9'd79,-10'd79};
ram[18737] = {-9'd76,-10'd76};
ram[18738] = {-9'd73,-10'd73};
ram[18739] = {-9'd70,-10'd70};
ram[18740] = {-9'd66,-10'd66};
ram[18741] = {-9'd63,-10'd63};
ram[18742] = {-9'd60,-10'd60};
ram[18743] = {-9'd57,-10'd57};
ram[18744] = {-9'd54,-10'd54};
ram[18745] = {-9'd51,-10'd51};
ram[18746] = {-9'd48,-10'd48};
ram[18747] = {-9'd44,-10'd44};
ram[18748] = {-9'd41,-10'd41};
ram[18749] = {-9'd38,-10'd38};
ram[18750] = {-9'd35,-10'd35};
ram[18751] = {-9'd32,-10'd32};
ram[18752] = {-9'd29,-10'd29};
ram[18753] = {-9'd26,-10'd26};
ram[18754] = {-9'd22,-10'd22};
ram[18755] = {-9'd19,-10'd19};
ram[18756] = {-9'd16,-10'd16};
ram[18757] = {-9'd13,-10'd13};
ram[18758] = {-9'd10,-10'd10};
ram[18759] = {-9'd7,-10'd7};
ram[18760] = {-9'd4,-10'd4};
ram[18761] = {9'd0,10'd0};
ram[18762] = {9'd3,10'd3};
ram[18763] = {9'd6,10'd6};
ram[18764] = {9'd9,10'd9};
ram[18765] = {9'd12,10'd12};
ram[18766] = {9'd15,10'd15};
ram[18767] = {9'd18,10'd18};
ram[18768] = {9'd21,10'd21};
ram[18769] = {9'd25,10'd25};
ram[18770] = {9'd28,10'd28};
ram[18771] = {9'd31,10'd31};
ram[18772] = {9'd34,10'd34};
ram[18773] = {9'd37,10'd37};
ram[18774] = {9'd40,10'd40};
ram[18775] = {9'd43,10'd43};
ram[18776] = {9'd47,10'd47};
ram[18777] = {9'd50,10'd50};
ram[18778] = {9'd53,10'd53};
ram[18779] = {9'd56,10'd56};
ram[18780] = {9'd59,10'd59};
ram[18781] = {9'd62,10'd62};
ram[18782] = {9'd65,10'd65};
ram[18783] = {9'd69,10'd69};
ram[18784] = {9'd72,10'd72};
ram[18785] = {9'd75,10'd75};
ram[18786] = {9'd78,10'd78};
ram[18787] = {9'd81,10'd81};
ram[18788] = {9'd84,10'd84};
ram[18789] = {9'd87,10'd87};
ram[18790] = {9'd91,10'd91};
ram[18791] = {9'd94,10'd94};
ram[18792] = {9'd97,10'd97};
ram[18793] = {-9'd100,10'd100};
ram[18794] = {-9'd97,10'd103};
ram[18795] = {-9'd94,10'd106};
ram[18796] = {-9'd91,10'd109};
ram[18797] = {-9'd88,10'd113};
ram[18798] = {-9'd85,10'd116};
ram[18799] = {-9'd81,10'd119};
ram[18800] = {-9'd78,10'd122};
ram[18801] = {-9'd75,10'd125};
ram[18802] = {-9'd72,10'd128};
ram[18803] = {-9'd69,10'd131};
ram[18804] = {-9'd66,10'd135};
ram[18805] = {-9'd63,10'd138};
ram[18806] = {-9'd59,10'd141};
ram[18807] = {-9'd56,10'd144};
ram[18808] = {-9'd53,10'd147};
ram[18809] = {-9'd50,10'd150};
ram[18810] = {-9'd47,10'd153};
ram[18811] = {-9'd44,10'd157};
ram[18812] = {-9'd41,10'd160};
ram[18813] = {-9'd37,10'd163};
ram[18814] = {-9'd34,10'd166};
ram[18815] = {-9'd31,10'd169};
ram[18816] = {-9'd31,10'd169};
ram[18817] = {-9'd28,10'd172};
ram[18818] = {-9'd25,10'd175};
ram[18819] = {-9'd22,10'd179};
ram[18820] = {-9'd19,10'd182};
ram[18821] = {-9'd15,10'd185};
ram[18822] = {-9'd12,10'd188};
ram[18823] = {-9'd9,10'd191};
ram[18824] = {-9'd6,10'd194};
ram[18825] = {-9'd3,10'd197};
ram[18826] = {9'd0,10'd201};
ram[18827] = {9'd3,10'd204};
ram[18828] = {9'd7,10'd207};
ram[18829] = {9'd10,10'd210};
ram[18830] = {9'd13,10'd213};
ram[18831] = {9'd16,10'd216};
ram[18832] = {9'd19,10'd219};
ram[18833] = {9'd22,10'd223};
ram[18834] = {9'd25,10'd226};
ram[18835] = {9'd29,10'd229};
ram[18836] = {9'd32,10'd232};
ram[18837] = {9'd35,10'd235};
ram[18838] = {9'd38,10'd238};
ram[18839] = {9'd41,10'd241};
ram[18840] = {9'd44,10'd245};
ram[18841] = {9'd47,10'd248};
ram[18842] = {9'd51,10'd251};
ram[18843] = {9'd54,10'd254};
ram[18844] = {9'd57,10'd257};
ram[18845] = {9'd60,10'd260};
ram[18846] = {9'd63,10'd263};
ram[18847] = {9'd66,10'd267};
ram[18848] = {9'd69,10'd270};
ram[18849] = {9'd73,10'd273};
ram[18850] = {9'd76,10'd276};
ram[18851] = {9'd79,10'd279};
ram[18852] = {9'd82,10'd282};
ram[18853] = {9'd85,10'd285};
ram[18854] = {9'd88,10'd289};
ram[18855] = {9'd91,10'd292};
ram[18856] = {9'd95,10'd295};
ram[18857] = {9'd98,10'd298};
ram[18858] = {-9'd99,10'd301};
ram[18859] = {-9'd96,10'd304};
ram[18860] = {-9'd93,10'd307};
ram[18861] = {-9'd90,10'd311};
ram[18862] = {-9'd87,10'd314};
ram[18863] = {-9'd84,10'd317};
ram[18864] = {-9'd81,10'd320};
ram[18865] = {-9'd77,10'd323};
ram[18866] = {-9'd74,10'd326};
ram[18867] = {-9'd71,10'd329};
ram[18868] = {-9'd68,10'd333};
ram[18869] = {-9'd65,10'd336};
ram[18870] = {-9'd62,10'd339};
ram[18871] = {-9'd59,10'd342};
ram[18872] = {-9'd55,10'd345};
ram[18873] = {-9'd52,10'd348};
ram[18874] = {-9'd49,10'd351};
ram[18875] = {-9'd46,10'd354};
ram[18876] = {-9'd43,10'd358};
ram[18877] = {-9'd40,10'd361};
ram[18878] = {-9'd37,10'd364};
ram[18879] = {-9'd33,10'd367};
ram[18880] = {-9'd30,10'd370};
ram[18881] = {-9'd27,10'd373};
ram[18882] = {-9'd24,10'd376};
ram[18883] = {-9'd21,10'd380};
ram[18884] = {-9'd18,10'd383};
ram[18885] = {-9'd15,10'd386};
ram[18886] = {-9'd11,10'd389};
ram[18887] = {-9'd8,10'd392};
ram[18888] = {-9'd5,10'd395};
ram[18889] = {-9'd2,10'd398};
ram[18890] = {9'd1,-10'd399};
ram[18891] = {9'd4,-10'd396};
ram[18892] = {9'd7,-10'd393};
ram[18893] = {9'd10,-10'd390};
ram[18894] = {9'd14,-10'd387};
ram[18895] = {9'd17,-10'd384};
ram[18896] = {9'd20,-10'd381};
ram[18897] = {9'd23,-10'd377};
ram[18898] = {9'd26,-10'd374};
ram[18899] = {9'd29,-10'd371};
ram[18900] = {9'd32,-10'd368};
ram[18901] = {9'd36,-10'd365};
ram[18902] = {9'd39,-10'd362};
ram[18903] = {9'd42,-10'd359};
ram[18904] = {9'd45,-10'd355};
ram[18905] = {9'd48,-10'd352};
ram[18906] = {9'd51,-10'd349};
ram[18907] = {9'd54,-10'd346};
ram[18908] = {9'd58,-10'd343};
ram[18909] = {9'd61,-10'd340};
ram[18910] = {9'd64,-10'd337};
ram[18911] = {9'd67,-10'd334};
ram[18912] = {9'd70,-10'd330};
ram[18913] = {9'd73,-10'd327};
ram[18914] = {9'd76,-10'd324};
ram[18915] = {9'd80,-10'd321};
ram[18916] = {9'd83,-10'd318};
ram[18917] = {9'd86,-10'd315};
ram[18918] = {9'd89,-10'd312};
ram[18919] = {9'd92,-10'd308};
ram[18920] = {9'd95,-10'd305};
ram[18921] = {9'd98,-10'd302};
ram[18922] = {-9'd99,-10'd299};
ram[18923] = {-9'd96,-10'd296};
ram[18924] = {-9'd92,-10'd293};
ram[18925] = {-9'd89,-10'd290};
ram[18926] = {-9'd86,-10'd286};
ram[18927] = {-9'd83,-10'd283};
ram[18928] = {-9'd80,-10'd280};
ram[18929] = {-9'd77,-10'd277};
ram[18930] = {-9'd74,-10'd274};
ram[18931] = {-9'd70,-10'd271};
ram[18932] = {-9'd67,-10'd268};
ram[18933] = {-9'd64,-10'd264};
ram[18934] = {-9'd61,-10'd261};
ram[18935] = {-9'd58,-10'd258};
ram[18936] = {-9'd55,-10'd255};
ram[18937] = {-9'd52,-10'd252};
ram[18938] = {-9'd48,-10'd249};
ram[18939] = {-9'd45,-10'd246};
ram[18940] = {-9'd42,-10'd242};
ram[18941] = {-9'd39,-10'd239};
ram[18942] = {-9'd36,-10'd236};
ram[18943] = {-9'd33,-10'd233};
ram[18944] = {-9'd33,-10'd233};
ram[18945] = {-9'd30,-10'd230};
ram[18946] = {-9'd26,-10'd227};
ram[18947] = {-9'd23,-10'd224};
ram[18948] = {-9'd20,-10'd220};
ram[18949] = {-9'd17,-10'd217};
ram[18950] = {-9'd14,-10'd214};
ram[18951] = {-9'd11,-10'd211};
ram[18952] = {-9'd8,-10'd208};
ram[18953] = {-9'd4,-10'd205};
ram[18954] = {-9'd1,-10'd202};
ram[18955] = {9'd2,-10'd198};
ram[18956] = {9'd5,-10'd195};
ram[18957] = {9'd8,-10'd192};
ram[18958] = {9'd11,-10'd189};
ram[18959] = {9'd14,-10'd186};
ram[18960] = {9'd18,-10'd183};
ram[18961] = {9'd21,-10'd180};
ram[18962] = {9'd24,-10'd176};
ram[18963] = {9'd27,-10'd173};
ram[18964] = {9'd30,-10'd170};
ram[18965] = {9'd33,-10'd167};
ram[18966] = {9'd36,-10'd164};
ram[18967] = {9'd40,-10'd161};
ram[18968] = {9'd43,-10'd158};
ram[18969] = {9'd46,-10'd154};
ram[18970] = {9'd49,-10'd151};
ram[18971] = {9'd52,-10'd148};
ram[18972] = {9'd55,-10'd145};
ram[18973] = {9'd58,-10'd142};
ram[18974] = {9'd62,-10'd139};
ram[18975] = {9'd65,-10'd136};
ram[18976] = {9'd68,-10'd132};
ram[18977] = {9'd71,-10'd129};
ram[18978] = {9'd74,-10'd126};
ram[18979] = {9'd77,-10'd123};
ram[18980] = {9'd80,-10'd120};
ram[18981] = {9'd84,-10'd117};
ram[18982] = {9'd87,-10'd114};
ram[18983] = {9'd90,-10'd110};
ram[18984] = {9'd93,-10'd107};
ram[18985] = {9'd96,-10'd104};
ram[18986] = {9'd99,-10'd101};
ram[18987] = {-9'd98,-10'd98};
ram[18988] = {-9'd95,-10'd95};
ram[18989] = {-9'd92,-10'd92};
ram[18990] = {-9'd88,-10'd88};
ram[18991] = {-9'd85,-10'd85};
ram[18992] = {-9'd82,-10'd82};
ram[18993] = {-9'd79,-10'd79};
ram[18994] = {-9'd76,-10'd76};
ram[18995] = {-9'd73,-10'd73};
ram[18996] = {-9'd70,-10'd70};
ram[18997] = {-9'd66,-10'd66};
ram[18998] = {-9'd63,-10'd63};
ram[18999] = {-9'd60,-10'd60};
ram[19000] = {-9'd57,-10'd57};
ram[19001] = {-9'd54,-10'd54};
ram[19002] = {-9'd51,-10'd51};
ram[19003] = {-9'd48,-10'd48};
ram[19004] = {-9'd44,-10'd44};
ram[19005] = {-9'd41,-10'd41};
ram[19006] = {-9'd38,-10'd38};
ram[19007] = {-9'd35,-10'd35};
ram[19008] = {-9'd32,-10'd32};
ram[19009] = {-9'd29,-10'd29};
ram[19010] = {-9'd26,-10'd26};
ram[19011] = {-9'd22,-10'd22};
ram[19012] = {-9'd19,-10'd19};
ram[19013] = {-9'd16,-10'd16};
ram[19014] = {-9'd13,-10'd13};
ram[19015] = {-9'd10,-10'd10};
ram[19016] = {-9'd7,-10'd7};
ram[19017] = {-9'd4,-10'd4};
ram[19018] = {9'd0,10'd0};
ram[19019] = {9'd3,10'd3};
ram[19020] = {9'd6,10'd6};
ram[19021] = {9'd9,10'd9};
ram[19022] = {9'd12,10'd12};
ram[19023] = {9'd15,10'd15};
ram[19024] = {9'd18,10'd18};
ram[19025] = {9'd21,10'd21};
ram[19026] = {9'd25,10'd25};
ram[19027] = {9'd28,10'd28};
ram[19028] = {9'd31,10'd31};
ram[19029] = {9'd34,10'd34};
ram[19030] = {9'd37,10'd37};
ram[19031] = {9'd40,10'd40};
ram[19032] = {9'd43,10'd43};
ram[19033] = {9'd47,10'd47};
ram[19034] = {9'd50,10'd50};
ram[19035] = {9'd53,10'd53};
ram[19036] = {9'd56,10'd56};
ram[19037] = {9'd59,10'd59};
ram[19038] = {9'd62,10'd62};
ram[19039] = {9'd65,10'd65};
ram[19040] = {9'd69,10'd69};
ram[19041] = {9'd72,10'd72};
ram[19042] = {9'd75,10'd75};
ram[19043] = {9'd78,10'd78};
ram[19044] = {9'd81,10'd81};
ram[19045] = {9'd84,10'd84};
ram[19046] = {9'd87,10'd87};
ram[19047] = {9'd91,10'd91};
ram[19048] = {9'd94,10'd94};
ram[19049] = {9'd97,10'd97};
ram[19050] = {-9'd100,10'd100};
ram[19051] = {-9'd97,10'd103};
ram[19052] = {-9'd94,10'd106};
ram[19053] = {-9'd91,10'd109};
ram[19054] = {-9'd88,10'd113};
ram[19055] = {-9'd85,10'd116};
ram[19056] = {-9'd81,10'd119};
ram[19057] = {-9'd78,10'd122};
ram[19058] = {-9'd75,10'd125};
ram[19059] = {-9'd72,10'd128};
ram[19060] = {-9'd69,10'd131};
ram[19061] = {-9'd66,10'd135};
ram[19062] = {-9'd63,10'd138};
ram[19063] = {-9'd59,10'd141};
ram[19064] = {-9'd56,10'd144};
ram[19065] = {-9'd53,10'd147};
ram[19066] = {-9'd50,10'd150};
ram[19067] = {-9'd47,10'd153};
ram[19068] = {-9'd44,10'd157};
ram[19069] = {-9'd41,10'd160};
ram[19070] = {-9'd37,10'd163};
ram[19071] = {-9'd34,10'd166};
ram[19072] = {-9'd34,10'd166};
ram[19073] = {-9'd31,10'd169};
ram[19074] = {-9'd28,10'd172};
ram[19075] = {-9'd25,10'd175};
ram[19076] = {-9'd22,10'd179};
ram[19077] = {-9'd19,10'd182};
ram[19078] = {-9'd15,10'd185};
ram[19079] = {-9'd12,10'd188};
ram[19080] = {-9'd9,10'd191};
ram[19081] = {-9'd6,10'd194};
ram[19082] = {-9'd3,10'd197};
ram[19083] = {9'd0,10'd201};
ram[19084] = {9'd3,10'd204};
ram[19085] = {9'd7,10'd207};
ram[19086] = {9'd10,10'd210};
ram[19087] = {9'd13,10'd213};
ram[19088] = {9'd16,10'd216};
ram[19089] = {9'd19,10'd219};
ram[19090] = {9'd22,10'd223};
ram[19091] = {9'd25,10'd226};
ram[19092] = {9'd29,10'd229};
ram[19093] = {9'd32,10'd232};
ram[19094] = {9'd35,10'd235};
ram[19095] = {9'd38,10'd238};
ram[19096] = {9'd41,10'd241};
ram[19097] = {9'd44,10'd245};
ram[19098] = {9'd47,10'd248};
ram[19099] = {9'd51,10'd251};
ram[19100] = {9'd54,10'd254};
ram[19101] = {9'd57,10'd257};
ram[19102] = {9'd60,10'd260};
ram[19103] = {9'd63,10'd263};
ram[19104] = {9'd66,10'd267};
ram[19105] = {9'd69,10'd270};
ram[19106] = {9'd73,10'd273};
ram[19107] = {9'd76,10'd276};
ram[19108] = {9'd79,10'd279};
ram[19109] = {9'd82,10'd282};
ram[19110] = {9'd85,10'd285};
ram[19111] = {9'd88,10'd289};
ram[19112] = {9'd91,10'd292};
ram[19113] = {9'd95,10'd295};
ram[19114] = {9'd98,10'd298};
ram[19115] = {-9'd99,10'd301};
ram[19116] = {-9'd96,10'd304};
ram[19117] = {-9'd93,10'd307};
ram[19118] = {-9'd90,10'd311};
ram[19119] = {-9'd87,10'd314};
ram[19120] = {-9'd84,10'd317};
ram[19121] = {-9'd81,10'd320};
ram[19122] = {-9'd77,10'd323};
ram[19123] = {-9'd74,10'd326};
ram[19124] = {-9'd71,10'd329};
ram[19125] = {-9'd68,10'd333};
ram[19126] = {-9'd65,10'd336};
ram[19127] = {-9'd62,10'd339};
ram[19128] = {-9'd59,10'd342};
ram[19129] = {-9'd55,10'd345};
ram[19130] = {-9'd52,10'd348};
ram[19131] = {-9'd49,10'd351};
ram[19132] = {-9'd46,10'd354};
ram[19133] = {-9'd43,10'd358};
ram[19134] = {-9'd40,10'd361};
ram[19135] = {-9'd37,10'd364};
ram[19136] = {-9'd33,10'd367};
ram[19137] = {-9'd30,10'd370};
ram[19138] = {-9'd27,10'd373};
ram[19139] = {-9'd24,10'd376};
ram[19140] = {-9'd21,10'd380};
ram[19141] = {-9'd18,10'd383};
ram[19142] = {-9'd15,10'd386};
ram[19143] = {-9'd11,10'd389};
ram[19144] = {-9'd8,10'd392};
ram[19145] = {-9'd5,10'd395};
ram[19146] = {-9'd2,10'd398};
ram[19147] = {9'd1,-10'd399};
ram[19148] = {9'd4,-10'd396};
ram[19149] = {9'd7,-10'd393};
ram[19150] = {9'd10,-10'd390};
ram[19151] = {9'd14,-10'd387};
ram[19152] = {9'd17,-10'd384};
ram[19153] = {9'd20,-10'd381};
ram[19154] = {9'd23,-10'd377};
ram[19155] = {9'd26,-10'd374};
ram[19156] = {9'd29,-10'd371};
ram[19157] = {9'd32,-10'd368};
ram[19158] = {9'd36,-10'd365};
ram[19159] = {9'd39,-10'd362};
ram[19160] = {9'd42,-10'd359};
ram[19161] = {9'd45,-10'd355};
ram[19162] = {9'd48,-10'd352};
ram[19163] = {9'd51,-10'd349};
ram[19164] = {9'd54,-10'd346};
ram[19165] = {9'd58,-10'd343};
ram[19166] = {9'd61,-10'd340};
ram[19167] = {9'd64,-10'd337};
ram[19168] = {9'd67,-10'd334};
ram[19169] = {9'd70,-10'd330};
ram[19170] = {9'd73,-10'd327};
ram[19171] = {9'd76,-10'd324};
ram[19172] = {9'd80,-10'd321};
ram[19173] = {9'd83,-10'd318};
ram[19174] = {9'd86,-10'd315};
ram[19175] = {9'd89,-10'd312};
ram[19176] = {9'd92,-10'd308};
ram[19177] = {9'd95,-10'd305};
ram[19178] = {9'd98,-10'd302};
ram[19179] = {-9'd99,-10'd299};
ram[19180] = {-9'd96,-10'd296};
ram[19181] = {-9'd92,-10'd293};
ram[19182] = {-9'd89,-10'd290};
ram[19183] = {-9'd86,-10'd286};
ram[19184] = {-9'd83,-10'd283};
ram[19185] = {-9'd80,-10'd280};
ram[19186] = {-9'd77,-10'd277};
ram[19187] = {-9'd74,-10'd274};
ram[19188] = {-9'd70,-10'd271};
ram[19189] = {-9'd67,-10'd268};
ram[19190] = {-9'd64,-10'd264};
ram[19191] = {-9'd61,-10'd261};
ram[19192] = {-9'd58,-10'd258};
ram[19193] = {-9'd55,-10'd255};
ram[19194] = {-9'd52,-10'd252};
ram[19195] = {-9'd48,-10'd249};
ram[19196] = {-9'd45,-10'd246};
ram[19197] = {-9'd42,-10'd242};
ram[19198] = {-9'd39,-10'd239};
ram[19199] = {-9'd36,-10'd236};
ram[19200] = {-9'd36,-10'd236};
ram[19201] = {-9'd33,-10'd233};
ram[19202] = {-9'd30,-10'd230};
ram[19203] = {-9'd26,-10'd227};
ram[19204] = {-9'd23,-10'd224};
ram[19205] = {-9'd20,-10'd220};
ram[19206] = {-9'd17,-10'd217};
ram[19207] = {-9'd14,-10'd214};
ram[19208] = {-9'd11,-10'd211};
ram[19209] = {-9'd8,-10'd208};
ram[19210] = {-9'd4,-10'd205};
ram[19211] = {-9'd1,-10'd202};
ram[19212] = {9'd2,-10'd198};
ram[19213] = {9'd5,-10'd195};
ram[19214] = {9'd8,-10'd192};
ram[19215] = {9'd11,-10'd189};
ram[19216] = {9'd14,-10'd186};
ram[19217] = {9'd18,-10'd183};
ram[19218] = {9'd21,-10'd180};
ram[19219] = {9'd24,-10'd176};
ram[19220] = {9'd27,-10'd173};
ram[19221] = {9'd30,-10'd170};
ram[19222] = {9'd33,-10'd167};
ram[19223] = {9'd36,-10'd164};
ram[19224] = {9'd40,-10'd161};
ram[19225] = {9'd43,-10'd158};
ram[19226] = {9'd46,-10'd154};
ram[19227] = {9'd49,-10'd151};
ram[19228] = {9'd52,-10'd148};
ram[19229] = {9'd55,-10'd145};
ram[19230] = {9'd58,-10'd142};
ram[19231] = {9'd62,-10'd139};
ram[19232] = {9'd65,-10'd136};
ram[19233] = {9'd68,-10'd132};
ram[19234] = {9'd71,-10'd129};
ram[19235] = {9'd74,-10'd126};
ram[19236] = {9'd77,-10'd123};
ram[19237] = {9'd80,-10'd120};
ram[19238] = {9'd84,-10'd117};
ram[19239] = {9'd87,-10'd114};
ram[19240] = {9'd90,-10'd110};
ram[19241] = {9'd93,-10'd107};
ram[19242] = {9'd96,-10'd104};
ram[19243] = {9'd99,-10'd101};
ram[19244] = {-9'd98,-10'd98};
ram[19245] = {-9'd95,-10'd95};
ram[19246] = {-9'd92,-10'd92};
ram[19247] = {-9'd88,-10'd88};
ram[19248] = {-9'd85,-10'd85};
ram[19249] = {-9'd82,-10'd82};
ram[19250] = {-9'd79,-10'd79};
ram[19251] = {-9'd76,-10'd76};
ram[19252] = {-9'd73,-10'd73};
ram[19253] = {-9'd70,-10'd70};
ram[19254] = {-9'd66,-10'd66};
ram[19255] = {-9'd63,-10'd63};
ram[19256] = {-9'd60,-10'd60};
ram[19257] = {-9'd57,-10'd57};
ram[19258] = {-9'd54,-10'd54};
ram[19259] = {-9'd51,-10'd51};
ram[19260] = {-9'd48,-10'd48};
ram[19261] = {-9'd44,-10'd44};
ram[19262] = {-9'd41,-10'd41};
ram[19263] = {-9'd38,-10'd38};
ram[19264] = {-9'd35,-10'd35};
ram[19265] = {-9'd32,-10'd32};
ram[19266] = {-9'd29,-10'd29};
ram[19267] = {-9'd26,-10'd26};
ram[19268] = {-9'd22,-10'd22};
ram[19269] = {-9'd19,-10'd19};
ram[19270] = {-9'd16,-10'd16};
ram[19271] = {-9'd13,-10'd13};
ram[19272] = {-9'd10,-10'd10};
ram[19273] = {-9'd7,-10'd7};
ram[19274] = {-9'd4,-10'd4};
ram[19275] = {9'd0,10'd0};
ram[19276] = {9'd3,10'd3};
ram[19277] = {9'd6,10'd6};
ram[19278] = {9'd9,10'd9};
ram[19279] = {9'd12,10'd12};
ram[19280] = {9'd15,10'd15};
ram[19281] = {9'd18,10'd18};
ram[19282] = {9'd21,10'd21};
ram[19283] = {9'd25,10'd25};
ram[19284] = {9'd28,10'd28};
ram[19285] = {9'd31,10'd31};
ram[19286] = {9'd34,10'd34};
ram[19287] = {9'd37,10'd37};
ram[19288] = {9'd40,10'd40};
ram[19289] = {9'd43,10'd43};
ram[19290] = {9'd47,10'd47};
ram[19291] = {9'd50,10'd50};
ram[19292] = {9'd53,10'd53};
ram[19293] = {9'd56,10'd56};
ram[19294] = {9'd59,10'd59};
ram[19295] = {9'd62,10'd62};
ram[19296] = {9'd65,10'd65};
ram[19297] = {9'd69,10'd69};
ram[19298] = {9'd72,10'd72};
ram[19299] = {9'd75,10'd75};
ram[19300] = {9'd78,10'd78};
ram[19301] = {9'd81,10'd81};
ram[19302] = {9'd84,10'd84};
ram[19303] = {9'd87,10'd87};
ram[19304] = {9'd91,10'd91};
ram[19305] = {9'd94,10'd94};
ram[19306] = {9'd97,10'd97};
ram[19307] = {-9'd100,10'd100};
ram[19308] = {-9'd97,10'd103};
ram[19309] = {-9'd94,10'd106};
ram[19310] = {-9'd91,10'd109};
ram[19311] = {-9'd88,10'd113};
ram[19312] = {-9'd85,10'd116};
ram[19313] = {-9'd81,10'd119};
ram[19314] = {-9'd78,10'd122};
ram[19315] = {-9'd75,10'd125};
ram[19316] = {-9'd72,10'd128};
ram[19317] = {-9'd69,10'd131};
ram[19318] = {-9'd66,10'd135};
ram[19319] = {-9'd63,10'd138};
ram[19320] = {-9'd59,10'd141};
ram[19321] = {-9'd56,10'd144};
ram[19322] = {-9'd53,10'd147};
ram[19323] = {-9'd50,10'd150};
ram[19324] = {-9'd47,10'd153};
ram[19325] = {-9'd44,10'd157};
ram[19326] = {-9'd41,10'd160};
ram[19327] = {-9'd37,10'd163};
ram[19328] = {-9'd37,10'd163};
ram[19329] = {-9'd34,10'd166};
ram[19330] = {-9'd31,10'd169};
ram[19331] = {-9'd28,10'd172};
ram[19332] = {-9'd25,10'd175};
ram[19333] = {-9'd22,10'd179};
ram[19334] = {-9'd19,10'd182};
ram[19335] = {-9'd15,10'd185};
ram[19336] = {-9'd12,10'd188};
ram[19337] = {-9'd9,10'd191};
ram[19338] = {-9'd6,10'd194};
ram[19339] = {-9'd3,10'd197};
ram[19340] = {9'd0,10'd201};
ram[19341] = {9'd3,10'd204};
ram[19342] = {9'd7,10'd207};
ram[19343] = {9'd10,10'd210};
ram[19344] = {9'd13,10'd213};
ram[19345] = {9'd16,10'd216};
ram[19346] = {9'd19,10'd219};
ram[19347] = {9'd22,10'd223};
ram[19348] = {9'd25,10'd226};
ram[19349] = {9'd29,10'd229};
ram[19350] = {9'd32,10'd232};
ram[19351] = {9'd35,10'd235};
ram[19352] = {9'd38,10'd238};
ram[19353] = {9'd41,10'd241};
ram[19354] = {9'd44,10'd245};
ram[19355] = {9'd47,10'd248};
ram[19356] = {9'd51,10'd251};
ram[19357] = {9'd54,10'd254};
ram[19358] = {9'd57,10'd257};
ram[19359] = {9'd60,10'd260};
ram[19360] = {9'd63,10'd263};
ram[19361] = {9'd66,10'd267};
ram[19362] = {9'd69,10'd270};
ram[19363] = {9'd73,10'd273};
ram[19364] = {9'd76,10'd276};
ram[19365] = {9'd79,10'd279};
ram[19366] = {9'd82,10'd282};
ram[19367] = {9'd85,10'd285};
ram[19368] = {9'd88,10'd289};
ram[19369] = {9'd91,10'd292};
ram[19370] = {9'd95,10'd295};
ram[19371] = {9'd98,10'd298};
ram[19372] = {-9'd99,10'd301};
ram[19373] = {-9'd96,10'd304};
ram[19374] = {-9'd93,10'd307};
ram[19375] = {-9'd90,10'd311};
ram[19376] = {-9'd87,10'd314};
ram[19377] = {-9'd84,10'd317};
ram[19378] = {-9'd81,10'd320};
ram[19379] = {-9'd77,10'd323};
ram[19380] = {-9'd74,10'd326};
ram[19381] = {-9'd71,10'd329};
ram[19382] = {-9'd68,10'd333};
ram[19383] = {-9'd65,10'd336};
ram[19384] = {-9'd62,10'd339};
ram[19385] = {-9'd59,10'd342};
ram[19386] = {-9'd55,10'd345};
ram[19387] = {-9'd52,10'd348};
ram[19388] = {-9'd49,10'd351};
ram[19389] = {-9'd46,10'd354};
ram[19390] = {-9'd43,10'd358};
ram[19391] = {-9'd40,10'd361};
ram[19392] = {-9'd37,10'd364};
ram[19393] = {-9'd33,10'd367};
ram[19394] = {-9'd30,10'd370};
ram[19395] = {-9'd27,10'd373};
ram[19396] = {-9'd24,10'd376};
ram[19397] = {-9'd21,10'd380};
ram[19398] = {-9'd18,10'd383};
ram[19399] = {-9'd15,10'd386};
ram[19400] = {-9'd11,10'd389};
ram[19401] = {-9'd8,10'd392};
ram[19402] = {-9'd5,10'd395};
ram[19403] = {-9'd2,10'd398};
ram[19404] = {9'd1,-10'd399};
ram[19405] = {9'd4,-10'd396};
ram[19406] = {9'd7,-10'd393};
ram[19407] = {9'd10,-10'd390};
ram[19408] = {9'd14,-10'd387};
ram[19409] = {9'd17,-10'd384};
ram[19410] = {9'd20,-10'd381};
ram[19411] = {9'd23,-10'd377};
ram[19412] = {9'd26,-10'd374};
ram[19413] = {9'd29,-10'd371};
ram[19414] = {9'd32,-10'd368};
ram[19415] = {9'd36,-10'd365};
ram[19416] = {9'd39,-10'd362};
ram[19417] = {9'd42,-10'd359};
ram[19418] = {9'd45,-10'd355};
ram[19419] = {9'd48,-10'd352};
ram[19420] = {9'd51,-10'd349};
ram[19421] = {9'd54,-10'd346};
ram[19422] = {9'd58,-10'd343};
ram[19423] = {9'd61,-10'd340};
ram[19424] = {9'd64,-10'd337};
ram[19425] = {9'd67,-10'd334};
ram[19426] = {9'd70,-10'd330};
ram[19427] = {9'd73,-10'd327};
ram[19428] = {9'd76,-10'd324};
ram[19429] = {9'd80,-10'd321};
ram[19430] = {9'd83,-10'd318};
ram[19431] = {9'd86,-10'd315};
ram[19432] = {9'd89,-10'd312};
ram[19433] = {9'd92,-10'd308};
ram[19434] = {9'd95,-10'd305};
ram[19435] = {9'd98,-10'd302};
ram[19436] = {-9'd99,-10'd299};
ram[19437] = {-9'd96,-10'd296};
ram[19438] = {-9'd92,-10'd293};
ram[19439] = {-9'd89,-10'd290};
ram[19440] = {-9'd86,-10'd286};
ram[19441] = {-9'd83,-10'd283};
ram[19442] = {-9'd80,-10'd280};
ram[19443] = {-9'd77,-10'd277};
ram[19444] = {-9'd74,-10'd274};
ram[19445] = {-9'd70,-10'd271};
ram[19446] = {-9'd67,-10'd268};
ram[19447] = {-9'd64,-10'd264};
ram[19448] = {-9'd61,-10'd261};
ram[19449] = {-9'd58,-10'd258};
ram[19450] = {-9'd55,-10'd255};
ram[19451] = {-9'd52,-10'd252};
ram[19452] = {-9'd48,-10'd249};
ram[19453] = {-9'd45,-10'd246};
ram[19454] = {-9'd42,-10'd242};
ram[19455] = {-9'd39,-10'd239};
ram[19456] = {-9'd39,-10'd239};
ram[19457] = {-9'd36,-10'd236};
ram[19458] = {-9'd33,-10'd233};
ram[19459] = {-9'd30,-10'd230};
ram[19460] = {-9'd26,-10'd227};
ram[19461] = {-9'd23,-10'd224};
ram[19462] = {-9'd20,-10'd220};
ram[19463] = {-9'd17,-10'd217};
ram[19464] = {-9'd14,-10'd214};
ram[19465] = {-9'd11,-10'd211};
ram[19466] = {-9'd8,-10'd208};
ram[19467] = {-9'd4,-10'd205};
ram[19468] = {-9'd1,-10'd202};
ram[19469] = {9'd2,-10'd198};
ram[19470] = {9'd5,-10'd195};
ram[19471] = {9'd8,-10'd192};
ram[19472] = {9'd11,-10'd189};
ram[19473] = {9'd14,-10'd186};
ram[19474] = {9'd18,-10'd183};
ram[19475] = {9'd21,-10'd180};
ram[19476] = {9'd24,-10'd176};
ram[19477] = {9'd27,-10'd173};
ram[19478] = {9'd30,-10'd170};
ram[19479] = {9'd33,-10'd167};
ram[19480] = {9'd36,-10'd164};
ram[19481] = {9'd40,-10'd161};
ram[19482] = {9'd43,-10'd158};
ram[19483] = {9'd46,-10'd154};
ram[19484] = {9'd49,-10'd151};
ram[19485] = {9'd52,-10'd148};
ram[19486] = {9'd55,-10'd145};
ram[19487] = {9'd58,-10'd142};
ram[19488] = {9'd62,-10'd139};
ram[19489] = {9'd65,-10'd136};
ram[19490] = {9'd68,-10'd132};
ram[19491] = {9'd71,-10'd129};
ram[19492] = {9'd74,-10'd126};
ram[19493] = {9'd77,-10'd123};
ram[19494] = {9'd80,-10'd120};
ram[19495] = {9'd84,-10'd117};
ram[19496] = {9'd87,-10'd114};
ram[19497] = {9'd90,-10'd110};
ram[19498] = {9'd93,-10'd107};
ram[19499] = {9'd96,-10'd104};
ram[19500] = {9'd99,-10'd101};
ram[19501] = {-9'd98,-10'd98};
ram[19502] = {-9'd95,-10'd95};
ram[19503] = {-9'd92,-10'd92};
ram[19504] = {-9'd88,-10'd88};
ram[19505] = {-9'd85,-10'd85};
ram[19506] = {-9'd82,-10'd82};
ram[19507] = {-9'd79,-10'd79};
ram[19508] = {-9'd76,-10'd76};
ram[19509] = {-9'd73,-10'd73};
ram[19510] = {-9'd70,-10'd70};
ram[19511] = {-9'd66,-10'd66};
ram[19512] = {-9'd63,-10'd63};
ram[19513] = {-9'd60,-10'd60};
ram[19514] = {-9'd57,-10'd57};
ram[19515] = {-9'd54,-10'd54};
ram[19516] = {-9'd51,-10'd51};
ram[19517] = {-9'd48,-10'd48};
ram[19518] = {-9'd44,-10'd44};
ram[19519] = {-9'd41,-10'd41};
ram[19520] = {-9'd38,-10'd38};
ram[19521] = {-9'd35,-10'd35};
ram[19522] = {-9'd32,-10'd32};
ram[19523] = {-9'd29,-10'd29};
ram[19524] = {-9'd26,-10'd26};
ram[19525] = {-9'd22,-10'd22};
ram[19526] = {-9'd19,-10'd19};
ram[19527] = {-9'd16,-10'd16};
ram[19528] = {-9'd13,-10'd13};
ram[19529] = {-9'd10,-10'd10};
ram[19530] = {-9'd7,-10'd7};
ram[19531] = {-9'd4,-10'd4};
ram[19532] = {9'd0,10'd0};
ram[19533] = {9'd3,10'd3};
ram[19534] = {9'd6,10'd6};
ram[19535] = {9'd9,10'd9};
ram[19536] = {9'd12,10'd12};
ram[19537] = {9'd15,10'd15};
ram[19538] = {9'd18,10'd18};
ram[19539] = {9'd21,10'd21};
ram[19540] = {9'd25,10'd25};
ram[19541] = {9'd28,10'd28};
ram[19542] = {9'd31,10'd31};
ram[19543] = {9'd34,10'd34};
ram[19544] = {9'd37,10'd37};
ram[19545] = {9'd40,10'd40};
ram[19546] = {9'd43,10'd43};
ram[19547] = {9'd47,10'd47};
ram[19548] = {9'd50,10'd50};
ram[19549] = {9'd53,10'd53};
ram[19550] = {9'd56,10'd56};
ram[19551] = {9'd59,10'd59};
ram[19552] = {9'd62,10'd62};
ram[19553] = {9'd65,10'd65};
ram[19554] = {9'd69,10'd69};
ram[19555] = {9'd72,10'd72};
ram[19556] = {9'd75,10'd75};
ram[19557] = {9'd78,10'd78};
ram[19558] = {9'd81,10'd81};
ram[19559] = {9'd84,10'd84};
ram[19560] = {9'd87,10'd87};
ram[19561] = {9'd91,10'd91};
ram[19562] = {9'd94,10'd94};
ram[19563] = {9'd97,10'd97};
ram[19564] = {-9'd100,10'd100};
ram[19565] = {-9'd97,10'd103};
ram[19566] = {-9'd94,10'd106};
ram[19567] = {-9'd91,10'd109};
ram[19568] = {-9'd88,10'd113};
ram[19569] = {-9'd85,10'd116};
ram[19570] = {-9'd81,10'd119};
ram[19571] = {-9'd78,10'd122};
ram[19572] = {-9'd75,10'd125};
ram[19573] = {-9'd72,10'd128};
ram[19574] = {-9'd69,10'd131};
ram[19575] = {-9'd66,10'd135};
ram[19576] = {-9'd63,10'd138};
ram[19577] = {-9'd59,10'd141};
ram[19578] = {-9'd56,10'd144};
ram[19579] = {-9'd53,10'd147};
ram[19580] = {-9'd50,10'd150};
ram[19581] = {-9'd47,10'd153};
ram[19582] = {-9'd44,10'd157};
ram[19583] = {-9'd41,10'd160};
ram[19584] = {-9'd41,10'd160};
ram[19585] = {-9'd37,10'd163};
ram[19586] = {-9'd34,10'd166};
ram[19587] = {-9'd31,10'd169};
ram[19588] = {-9'd28,10'd172};
ram[19589] = {-9'd25,10'd175};
ram[19590] = {-9'd22,10'd179};
ram[19591] = {-9'd19,10'd182};
ram[19592] = {-9'd15,10'd185};
ram[19593] = {-9'd12,10'd188};
ram[19594] = {-9'd9,10'd191};
ram[19595] = {-9'd6,10'd194};
ram[19596] = {-9'd3,10'd197};
ram[19597] = {9'd0,10'd201};
ram[19598] = {9'd3,10'd204};
ram[19599] = {9'd7,10'd207};
ram[19600] = {9'd10,10'd210};
ram[19601] = {9'd13,10'd213};
ram[19602] = {9'd16,10'd216};
ram[19603] = {9'd19,10'd219};
ram[19604] = {9'd22,10'd223};
ram[19605] = {9'd25,10'd226};
ram[19606] = {9'd29,10'd229};
ram[19607] = {9'd32,10'd232};
ram[19608] = {9'd35,10'd235};
ram[19609] = {9'd38,10'd238};
ram[19610] = {9'd41,10'd241};
ram[19611] = {9'd44,10'd245};
ram[19612] = {9'd47,10'd248};
ram[19613] = {9'd51,10'd251};
ram[19614] = {9'd54,10'd254};
ram[19615] = {9'd57,10'd257};
ram[19616] = {9'd60,10'd260};
ram[19617] = {9'd63,10'd263};
ram[19618] = {9'd66,10'd267};
ram[19619] = {9'd69,10'd270};
ram[19620] = {9'd73,10'd273};
ram[19621] = {9'd76,10'd276};
ram[19622] = {9'd79,10'd279};
ram[19623] = {9'd82,10'd282};
ram[19624] = {9'd85,10'd285};
ram[19625] = {9'd88,10'd289};
ram[19626] = {9'd91,10'd292};
ram[19627] = {9'd95,10'd295};
ram[19628] = {9'd98,10'd298};
ram[19629] = {-9'd99,10'd301};
ram[19630] = {-9'd96,10'd304};
ram[19631] = {-9'd93,10'd307};
ram[19632] = {-9'd90,10'd311};
ram[19633] = {-9'd87,10'd314};
ram[19634] = {-9'd84,10'd317};
ram[19635] = {-9'd81,10'd320};
ram[19636] = {-9'd77,10'd323};
ram[19637] = {-9'd74,10'd326};
ram[19638] = {-9'd71,10'd329};
ram[19639] = {-9'd68,10'd333};
ram[19640] = {-9'd65,10'd336};
ram[19641] = {-9'd62,10'd339};
ram[19642] = {-9'd59,10'd342};
ram[19643] = {-9'd55,10'd345};
ram[19644] = {-9'd52,10'd348};
ram[19645] = {-9'd49,10'd351};
ram[19646] = {-9'd46,10'd354};
ram[19647] = {-9'd43,10'd358};
ram[19648] = {-9'd40,10'd361};
ram[19649] = {-9'd37,10'd364};
ram[19650] = {-9'd33,10'd367};
ram[19651] = {-9'd30,10'd370};
ram[19652] = {-9'd27,10'd373};
ram[19653] = {-9'd24,10'd376};
ram[19654] = {-9'd21,10'd380};
ram[19655] = {-9'd18,10'd383};
ram[19656] = {-9'd15,10'd386};
ram[19657] = {-9'd11,10'd389};
ram[19658] = {-9'd8,10'd392};
ram[19659] = {-9'd5,10'd395};
ram[19660] = {-9'd2,10'd398};
ram[19661] = {9'd1,-10'd399};
ram[19662] = {9'd4,-10'd396};
ram[19663] = {9'd7,-10'd393};
ram[19664] = {9'd10,-10'd390};
ram[19665] = {9'd14,-10'd387};
ram[19666] = {9'd17,-10'd384};
ram[19667] = {9'd20,-10'd381};
ram[19668] = {9'd23,-10'd377};
ram[19669] = {9'd26,-10'd374};
ram[19670] = {9'd29,-10'd371};
ram[19671] = {9'd32,-10'd368};
ram[19672] = {9'd36,-10'd365};
ram[19673] = {9'd39,-10'd362};
ram[19674] = {9'd42,-10'd359};
ram[19675] = {9'd45,-10'd355};
ram[19676] = {9'd48,-10'd352};
ram[19677] = {9'd51,-10'd349};
ram[19678] = {9'd54,-10'd346};
ram[19679] = {9'd58,-10'd343};
ram[19680] = {9'd61,-10'd340};
ram[19681] = {9'd64,-10'd337};
ram[19682] = {9'd67,-10'd334};
ram[19683] = {9'd70,-10'd330};
ram[19684] = {9'd73,-10'd327};
ram[19685] = {9'd76,-10'd324};
ram[19686] = {9'd80,-10'd321};
ram[19687] = {9'd83,-10'd318};
ram[19688] = {9'd86,-10'd315};
ram[19689] = {9'd89,-10'd312};
ram[19690] = {9'd92,-10'd308};
ram[19691] = {9'd95,-10'd305};
ram[19692] = {9'd98,-10'd302};
ram[19693] = {-9'd99,-10'd299};
ram[19694] = {-9'd96,-10'd296};
ram[19695] = {-9'd92,-10'd293};
ram[19696] = {-9'd89,-10'd290};
ram[19697] = {-9'd86,-10'd286};
ram[19698] = {-9'd83,-10'd283};
ram[19699] = {-9'd80,-10'd280};
ram[19700] = {-9'd77,-10'd277};
ram[19701] = {-9'd74,-10'd274};
ram[19702] = {-9'd70,-10'd271};
ram[19703] = {-9'd67,-10'd268};
ram[19704] = {-9'd64,-10'd264};
ram[19705] = {-9'd61,-10'd261};
ram[19706] = {-9'd58,-10'd258};
ram[19707] = {-9'd55,-10'd255};
ram[19708] = {-9'd52,-10'd252};
ram[19709] = {-9'd48,-10'd249};
ram[19710] = {-9'd45,-10'd246};
ram[19711] = {-9'd42,-10'd242};
ram[19712] = {-9'd42,-10'd242};
ram[19713] = {-9'd39,-10'd239};
ram[19714] = {-9'd36,-10'd236};
ram[19715] = {-9'd33,-10'd233};
ram[19716] = {-9'd30,-10'd230};
ram[19717] = {-9'd26,-10'd227};
ram[19718] = {-9'd23,-10'd224};
ram[19719] = {-9'd20,-10'd220};
ram[19720] = {-9'd17,-10'd217};
ram[19721] = {-9'd14,-10'd214};
ram[19722] = {-9'd11,-10'd211};
ram[19723] = {-9'd8,-10'd208};
ram[19724] = {-9'd4,-10'd205};
ram[19725] = {-9'd1,-10'd202};
ram[19726] = {9'd2,-10'd198};
ram[19727] = {9'd5,-10'd195};
ram[19728] = {9'd8,-10'd192};
ram[19729] = {9'd11,-10'd189};
ram[19730] = {9'd14,-10'd186};
ram[19731] = {9'd18,-10'd183};
ram[19732] = {9'd21,-10'd180};
ram[19733] = {9'd24,-10'd176};
ram[19734] = {9'd27,-10'd173};
ram[19735] = {9'd30,-10'd170};
ram[19736] = {9'd33,-10'd167};
ram[19737] = {9'd36,-10'd164};
ram[19738] = {9'd40,-10'd161};
ram[19739] = {9'd43,-10'd158};
ram[19740] = {9'd46,-10'd154};
ram[19741] = {9'd49,-10'd151};
ram[19742] = {9'd52,-10'd148};
ram[19743] = {9'd55,-10'd145};
ram[19744] = {9'd58,-10'd142};
ram[19745] = {9'd62,-10'd139};
ram[19746] = {9'd65,-10'd136};
ram[19747] = {9'd68,-10'd132};
ram[19748] = {9'd71,-10'd129};
ram[19749] = {9'd74,-10'd126};
ram[19750] = {9'd77,-10'd123};
ram[19751] = {9'd80,-10'd120};
ram[19752] = {9'd84,-10'd117};
ram[19753] = {9'd87,-10'd114};
ram[19754] = {9'd90,-10'd110};
ram[19755] = {9'd93,-10'd107};
ram[19756] = {9'd96,-10'd104};
ram[19757] = {9'd99,-10'd101};
ram[19758] = {-9'd98,-10'd98};
ram[19759] = {-9'd95,-10'd95};
ram[19760] = {-9'd92,-10'd92};
ram[19761] = {-9'd88,-10'd88};
ram[19762] = {-9'd85,-10'd85};
ram[19763] = {-9'd82,-10'd82};
ram[19764] = {-9'd79,-10'd79};
ram[19765] = {-9'd76,-10'd76};
ram[19766] = {-9'd73,-10'd73};
ram[19767] = {-9'd70,-10'd70};
ram[19768] = {-9'd66,-10'd66};
ram[19769] = {-9'd63,-10'd63};
ram[19770] = {-9'd60,-10'd60};
ram[19771] = {-9'd57,-10'd57};
ram[19772] = {-9'd54,-10'd54};
ram[19773] = {-9'd51,-10'd51};
ram[19774] = {-9'd48,-10'd48};
ram[19775] = {-9'd44,-10'd44};
ram[19776] = {-9'd41,-10'd41};
ram[19777] = {-9'd38,-10'd38};
ram[19778] = {-9'd35,-10'd35};
ram[19779] = {-9'd32,-10'd32};
ram[19780] = {-9'd29,-10'd29};
ram[19781] = {-9'd26,-10'd26};
ram[19782] = {-9'd22,-10'd22};
ram[19783] = {-9'd19,-10'd19};
ram[19784] = {-9'd16,-10'd16};
ram[19785] = {-9'd13,-10'd13};
ram[19786] = {-9'd10,-10'd10};
ram[19787] = {-9'd7,-10'd7};
ram[19788] = {-9'd4,-10'd4};
ram[19789] = {9'd0,10'd0};
ram[19790] = {9'd3,10'd3};
ram[19791] = {9'd6,10'd6};
ram[19792] = {9'd9,10'd9};
ram[19793] = {9'd12,10'd12};
ram[19794] = {9'd15,10'd15};
ram[19795] = {9'd18,10'd18};
ram[19796] = {9'd21,10'd21};
ram[19797] = {9'd25,10'd25};
ram[19798] = {9'd28,10'd28};
ram[19799] = {9'd31,10'd31};
ram[19800] = {9'd34,10'd34};
ram[19801] = {9'd37,10'd37};
ram[19802] = {9'd40,10'd40};
ram[19803] = {9'd43,10'd43};
ram[19804] = {9'd47,10'd47};
ram[19805] = {9'd50,10'd50};
ram[19806] = {9'd53,10'd53};
ram[19807] = {9'd56,10'd56};
ram[19808] = {9'd59,10'd59};
ram[19809] = {9'd62,10'd62};
ram[19810] = {9'd65,10'd65};
ram[19811] = {9'd69,10'd69};
ram[19812] = {9'd72,10'd72};
ram[19813] = {9'd75,10'd75};
ram[19814] = {9'd78,10'd78};
ram[19815] = {9'd81,10'd81};
ram[19816] = {9'd84,10'd84};
ram[19817] = {9'd87,10'd87};
ram[19818] = {9'd91,10'd91};
ram[19819] = {9'd94,10'd94};
ram[19820] = {9'd97,10'd97};
ram[19821] = {-9'd100,10'd100};
ram[19822] = {-9'd97,10'd103};
ram[19823] = {-9'd94,10'd106};
ram[19824] = {-9'd91,10'd109};
ram[19825] = {-9'd88,10'd113};
ram[19826] = {-9'd85,10'd116};
ram[19827] = {-9'd81,10'd119};
ram[19828] = {-9'd78,10'd122};
ram[19829] = {-9'd75,10'd125};
ram[19830] = {-9'd72,10'd128};
ram[19831] = {-9'd69,10'd131};
ram[19832] = {-9'd66,10'd135};
ram[19833] = {-9'd63,10'd138};
ram[19834] = {-9'd59,10'd141};
ram[19835] = {-9'd56,10'd144};
ram[19836] = {-9'd53,10'd147};
ram[19837] = {-9'd50,10'd150};
ram[19838] = {-9'd47,10'd153};
ram[19839] = {-9'd44,10'd157};
ram[19840] = {-9'd44,10'd157};
ram[19841] = {-9'd41,10'd160};
ram[19842] = {-9'd37,10'd163};
ram[19843] = {-9'd34,10'd166};
ram[19844] = {-9'd31,10'd169};
ram[19845] = {-9'd28,10'd172};
ram[19846] = {-9'd25,10'd175};
ram[19847] = {-9'd22,10'd179};
ram[19848] = {-9'd19,10'd182};
ram[19849] = {-9'd15,10'd185};
ram[19850] = {-9'd12,10'd188};
ram[19851] = {-9'd9,10'd191};
ram[19852] = {-9'd6,10'd194};
ram[19853] = {-9'd3,10'd197};
ram[19854] = {9'd0,10'd201};
ram[19855] = {9'd3,10'd204};
ram[19856] = {9'd7,10'd207};
ram[19857] = {9'd10,10'd210};
ram[19858] = {9'd13,10'd213};
ram[19859] = {9'd16,10'd216};
ram[19860] = {9'd19,10'd219};
ram[19861] = {9'd22,10'd223};
ram[19862] = {9'd25,10'd226};
ram[19863] = {9'd29,10'd229};
ram[19864] = {9'd32,10'd232};
ram[19865] = {9'd35,10'd235};
ram[19866] = {9'd38,10'd238};
ram[19867] = {9'd41,10'd241};
ram[19868] = {9'd44,10'd245};
ram[19869] = {9'd47,10'd248};
ram[19870] = {9'd51,10'd251};
ram[19871] = {9'd54,10'd254};
ram[19872] = {9'd57,10'd257};
ram[19873] = {9'd60,10'd260};
ram[19874] = {9'd63,10'd263};
ram[19875] = {9'd66,10'd267};
ram[19876] = {9'd69,10'd270};
ram[19877] = {9'd73,10'd273};
ram[19878] = {9'd76,10'd276};
ram[19879] = {9'd79,10'd279};
ram[19880] = {9'd82,10'd282};
ram[19881] = {9'd85,10'd285};
ram[19882] = {9'd88,10'd289};
ram[19883] = {9'd91,10'd292};
ram[19884] = {9'd95,10'd295};
ram[19885] = {9'd98,10'd298};
ram[19886] = {-9'd99,10'd301};
ram[19887] = {-9'd96,10'd304};
ram[19888] = {-9'd93,10'd307};
ram[19889] = {-9'd90,10'd311};
ram[19890] = {-9'd87,10'd314};
ram[19891] = {-9'd84,10'd317};
ram[19892] = {-9'd81,10'd320};
ram[19893] = {-9'd77,10'd323};
ram[19894] = {-9'd74,10'd326};
ram[19895] = {-9'd71,10'd329};
ram[19896] = {-9'd68,10'd333};
ram[19897] = {-9'd65,10'd336};
ram[19898] = {-9'd62,10'd339};
ram[19899] = {-9'd59,10'd342};
ram[19900] = {-9'd55,10'd345};
ram[19901] = {-9'd52,10'd348};
ram[19902] = {-9'd49,10'd351};
ram[19903] = {-9'd46,10'd354};
ram[19904] = {-9'd43,10'd358};
ram[19905] = {-9'd40,10'd361};
ram[19906] = {-9'd37,10'd364};
ram[19907] = {-9'd33,10'd367};
ram[19908] = {-9'd30,10'd370};
ram[19909] = {-9'd27,10'd373};
ram[19910] = {-9'd24,10'd376};
ram[19911] = {-9'd21,10'd380};
ram[19912] = {-9'd18,10'd383};
ram[19913] = {-9'd15,10'd386};
ram[19914] = {-9'd11,10'd389};
ram[19915] = {-9'd8,10'd392};
ram[19916] = {-9'd5,10'd395};
ram[19917] = {-9'd2,10'd398};
ram[19918] = {9'd1,-10'd399};
ram[19919] = {9'd4,-10'd396};
ram[19920] = {9'd7,-10'd393};
ram[19921] = {9'd10,-10'd390};
ram[19922] = {9'd14,-10'd387};
ram[19923] = {9'd17,-10'd384};
ram[19924] = {9'd20,-10'd381};
ram[19925] = {9'd23,-10'd377};
ram[19926] = {9'd26,-10'd374};
ram[19927] = {9'd29,-10'd371};
ram[19928] = {9'd32,-10'd368};
ram[19929] = {9'd36,-10'd365};
ram[19930] = {9'd39,-10'd362};
ram[19931] = {9'd42,-10'd359};
ram[19932] = {9'd45,-10'd355};
ram[19933] = {9'd48,-10'd352};
ram[19934] = {9'd51,-10'd349};
ram[19935] = {9'd54,-10'd346};
ram[19936] = {9'd58,-10'd343};
ram[19937] = {9'd61,-10'd340};
ram[19938] = {9'd64,-10'd337};
ram[19939] = {9'd67,-10'd334};
ram[19940] = {9'd70,-10'd330};
ram[19941] = {9'd73,-10'd327};
ram[19942] = {9'd76,-10'd324};
ram[19943] = {9'd80,-10'd321};
ram[19944] = {9'd83,-10'd318};
ram[19945] = {9'd86,-10'd315};
ram[19946] = {9'd89,-10'd312};
ram[19947] = {9'd92,-10'd308};
ram[19948] = {9'd95,-10'd305};
ram[19949] = {9'd98,-10'd302};
ram[19950] = {-9'd99,-10'd299};
ram[19951] = {-9'd96,-10'd296};
ram[19952] = {-9'd92,-10'd293};
ram[19953] = {-9'd89,-10'd290};
ram[19954] = {-9'd86,-10'd286};
ram[19955] = {-9'd83,-10'd283};
ram[19956] = {-9'd80,-10'd280};
ram[19957] = {-9'd77,-10'd277};
ram[19958] = {-9'd74,-10'd274};
ram[19959] = {-9'd70,-10'd271};
ram[19960] = {-9'd67,-10'd268};
ram[19961] = {-9'd64,-10'd264};
ram[19962] = {-9'd61,-10'd261};
ram[19963] = {-9'd58,-10'd258};
ram[19964] = {-9'd55,-10'd255};
ram[19965] = {-9'd52,-10'd252};
ram[19966] = {-9'd48,-10'd249};
ram[19967] = {-9'd45,-10'd246};
ram[19968] = {-9'd45,-10'd246};
ram[19969] = {-9'd42,-10'd242};
ram[19970] = {-9'd39,-10'd239};
ram[19971] = {-9'd36,-10'd236};
ram[19972] = {-9'd33,-10'd233};
ram[19973] = {-9'd30,-10'd230};
ram[19974] = {-9'd26,-10'd227};
ram[19975] = {-9'd23,-10'd224};
ram[19976] = {-9'd20,-10'd220};
ram[19977] = {-9'd17,-10'd217};
ram[19978] = {-9'd14,-10'd214};
ram[19979] = {-9'd11,-10'd211};
ram[19980] = {-9'd8,-10'd208};
ram[19981] = {-9'd4,-10'd205};
ram[19982] = {-9'd1,-10'd202};
ram[19983] = {9'd2,-10'd198};
ram[19984] = {9'd5,-10'd195};
ram[19985] = {9'd8,-10'd192};
ram[19986] = {9'd11,-10'd189};
ram[19987] = {9'd14,-10'd186};
ram[19988] = {9'd18,-10'd183};
ram[19989] = {9'd21,-10'd180};
ram[19990] = {9'd24,-10'd176};
ram[19991] = {9'd27,-10'd173};
ram[19992] = {9'd30,-10'd170};
ram[19993] = {9'd33,-10'd167};
ram[19994] = {9'd36,-10'd164};
ram[19995] = {9'd40,-10'd161};
ram[19996] = {9'd43,-10'd158};
ram[19997] = {9'd46,-10'd154};
ram[19998] = {9'd49,-10'd151};
ram[19999] = {9'd52,-10'd148};
ram[20000] = {9'd55,-10'd145};
ram[20001] = {9'd58,-10'd142};
ram[20002] = {9'd62,-10'd139};
ram[20003] = {9'd65,-10'd136};
ram[20004] = {9'd68,-10'd132};
ram[20005] = {9'd71,-10'd129};
ram[20006] = {9'd74,-10'd126};
ram[20007] = {9'd77,-10'd123};
ram[20008] = {9'd80,-10'd120};
ram[20009] = {9'd84,-10'd117};
ram[20010] = {9'd87,-10'd114};
ram[20011] = {9'd90,-10'd110};
ram[20012] = {9'd93,-10'd107};
ram[20013] = {9'd96,-10'd104};
ram[20014] = {9'd99,-10'd101};
ram[20015] = {-9'd98,-10'd98};
ram[20016] = {-9'd95,-10'd95};
ram[20017] = {-9'd92,-10'd92};
ram[20018] = {-9'd88,-10'd88};
ram[20019] = {-9'd85,-10'd85};
ram[20020] = {-9'd82,-10'd82};
ram[20021] = {-9'd79,-10'd79};
ram[20022] = {-9'd76,-10'd76};
ram[20023] = {-9'd73,-10'd73};
ram[20024] = {-9'd70,-10'd70};
ram[20025] = {-9'd66,-10'd66};
ram[20026] = {-9'd63,-10'd63};
ram[20027] = {-9'd60,-10'd60};
ram[20028] = {-9'd57,-10'd57};
ram[20029] = {-9'd54,-10'd54};
ram[20030] = {-9'd51,-10'd51};
ram[20031] = {-9'd48,-10'd48};
ram[20032] = {-9'd44,-10'd44};
ram[20033] = {-9'd41,-10'd41};
ram[20034] = {-9'd38,-10'd38};
ram[20035] = {-9'd35,-10'd35};
ram[20036] = {-9'd32,-10'd32};
ram[20037] = {-9'd29,-10'd29};
ram[20038] = {-9'd26,-10'd26};
ram[20039] = {-9'd22,-10'd22};
ram[20040] = {-9'd19,-10'd19};
ram[20041] = {-9'd16,-10'd16};
ram[20042] = {-9'd13,-10'd13};
ram[20043] = {-9'd10,-10'd10};
ram[20044] = {-9'd7,-10'd7};
ram[20045] = {-9'd4,-10'd4};
ram[20046] = {9'd0,10'd0};
ram[20047] = {9'd3,10'd3};
ram[20048] = {9'd6,10'd6};
ram[20049] = {9'd9,10'd9};
ram[20050] = {9'd12,10'd12};
ram[20051] = {9'd15,10'd15};
ram[20052] = {9'd18,10'd18};
ram[20053] = {9'd21,10'd21};
ram[20054] = {9'd25,10'd25};
ram[20055] = {9'd28,10'd28};
ram[20056] = {9'd31,10'd31};
ram[20057] = {9'd34,10'd34};
ram[20058] = {9'd37,10'd37};
ram[20059] = {9'd40,10'd40};
ram[20060] = {9'd43,10'd43};
ram[20061] = {9'd47,10'd47};
ram[20062] = {9'd50,10'd50};
ram[20063] = {9'd53,10'd53};
ram[20064] = {9'd56,10'd56};
ram[20065] = {9'd59,10'd59};
ram[20066] = {9'd62,10'd62};
ram[20067] = {9'd65,10'd65};
ram[20068] = {9'd69,10'd69};
ram[20069] = {9'd72,10'd72};
ram[20070] = {9'd75,10'd75};
ram[20071] = {9'd78,10'd78};
ram[20072] = {9'd81,10'd81};
ram[20073] = {9'd84,10'd84};
ram[20074] = {9'd87,10'd87};
ram[20075] = {9'd91,10'd91};
ram[20076] = {9'd94,10'd94};
ram[20077] = {9'd97,10'd97};
ram[20078] = {-9'd100,10'd100};
ram[20079] = {-9'd97,10'd103};
ram[20080] = {-9'd94,10'd106};
ram[20081] = {-9'd91,10'd109};
ram[20082] = {-9'd88,10'd113};
ram[20083] = {-9'd85,10'd116};
ram[20084] = {-9'd81,10'd119};
ram[20085] = {-9'd78,10'd122};
ram[20086] = {-9'd75,10'd125};
ram[20087] = {-9'd72,10'd128};
ram[20088] = {-9'd69,10'd131};
ram[20089] = {-9'd66,10'd135};
ram[20090] = {-9'd63,10'd138};
ram[20091] = {-9'd59,10'd141};
ram[20092] = {-9'd56,10'd144};
ram[20093] = {-9'd53,10'd147};
ram[20094] = {-9'd50,10'd150};
ram[20095] = {-9'd47,10'd153};
ram[20096] = {-9'd47,10'd153};
ram[20097] = {-9'd44,10'd157};
ram[20098] = {-9'd41,10'd160};
ram[20099] = {-9'd37,10'd163};
ram[20100] = {-9'd34,10'd166};
ram[20101] = {-9'd31,10'd169};
ram[20102] = {-9'd28,10'd172};
ram[20103] = {-9'd25,10'd175};
ram[20104] = {-9'd22,10'd179};
ram[20105] = {-9'd19,10'd182};
ram[20106] = {-9'd15,10'd185};
ram[20107] = {-9'd12,10'd188};
ram[20108] = {-9'd9,10'd191};
ram[20109] = {-9'd6,10'd194};
ram[20110] = {-9'd3,10'd197};
ram[20111] = {9'd0,10'd201};
ram[20112] = {9'd3,10'd204};
ram[20113] = {9'd7,10'd207};
ram[20114] = {9'd10,10'd210};
ram[20115] = {9'd13,10'd213};
ram[20116] = {9'd16,10'd216};
ram[20117] = {9'd19,10'd219};
ram[20118] = {9'd22,10'd223};
ram[20119] = {9'd25,10'd226};
ram[20120] = {9'd29,10'd229};
ram[20121] = {9'd32,10'd232};
ram[20122] = {9'd35,10'd235};
ram[20123] = {9'd38,10'd238};
ram[20124] = {9'd41,10'd241};
ram[20125] = {9'd44,10'd245};
ram[20126] = {9'd47,10'd248};
ram[20127] = {9'd51,10'd251};
ram[20128] = {9'd54,10'd254};
ram[20129] = {9'd57,10'd257};
ram[20130] = {9'd60,10'd260};
ram[20131] = {9'd63,10'd263};
ram[20132] = {9'd66,10'd267};
ram[20133] = {9'd69,10'd270};
ram[20134] = {9'd73,10'd273};
ram[20135] = {9'd76,10'd276};
ram[20136] = {9'd79,10'd279};
ram[20137] = {9'd82,10'd282};
ram[20138] = {9'd85,10'd285};
ram[20139] = {9'd88,10'd289};
ram[20140] = {9'd91,10'd292};
ram[20141] = {9'd95,10'd295};
ram[20142] = {9'd98,10'd298};
ram[20143] = {-9'd99,10'd301};
ram[20144] = {-9'd96,10'd304};
ram[20145] = {-9'd93,10'd307};
ram[20146] = {-9'd90,10'd311};
ram[20147] = {-9'd87,10'd314};
ram[20148] = {-9'd84,10'd317};
ram[20149] = {-9'd81,10'd320};
ram[20150] = {-9'd77,10'd323};
ram[20151] = {-9'd74,10'd326};
ram[20152] = {-9'd71,10'd329};
ram[20153] = {-9'd68,10'd333};
ram[20154] = {-9'd65,10'd336};
ram[20155] = {-9'd62,10'd339};
ram[20156] = {-9'd59,10'd342};
ram[20157] = {-9'd55,10'd345};
ram[20158] = {-9'd52,10'd348};
ram[20159] = {-9'd49,10'd351};
ram[20160] = {-9'd46,10'd354};
ram[20161] = {-9'd43,10'd358};
ram[20162] = {-9'd40,10'd361};
ram[20163] = {-9'd37,10'd364};
ram[20164] = {-9'd33,10'd367};
ram[20165] = {-9'd30,10'd370};
ram[20166] = {-9'd27,10'd373};
ram[20167] = {-9'd24,10'd376};
ram[20168] = {-9'd21,10'd380};
ram[20169] = {-9'd18,10'd383};
ram[20170] = {-9'd15,10'd386};
ram[20171] = {-9'd11,10'd389};
ram[20172] = {-9'd8,10'd392};
ram[20173] = {-9'd5,10'd395};
ram[20174] = {-9'd2,10'd398};
ram[20175] = {9'd1,-10'd399};
ram[20176] = {9'd4,-10'd396};
ram[20177] = {9'd7,-10'd393};
ram[20178] = {9'd10,-10'd390};
ram[20179] = {9'd14,-10'd387};
ram[20180] = {9'd17,-10'd384};
ram[20181] = {9'd20,-10'd381};
ram[20182] = {9'd23,-10'd377};
ram[20183] = {9'd26,-10'd374};
ram[20184] = {9'd29,-10'd371};
ram[20185] = {9'd32,-10'd368};
ram[20186] = {9'd36,-10'd365};
ram[20187] = {9'd39,-10'd362};
ram[20188] = {9'd42,-10'd359};
ram[20189] = {9'd45,-10'd355};
ram[20190] = {9'd48,-10'd352};
ram[20191] = {9'd51,-10'd349};
ram[20192] = {9'd54,-10'd346};
ram[20193] = {9'd58,-10'd343};
ram[20194] = {9'd61,-10'd340};
ram[20195] = {9'd64,-10'd337};
ram[20196] = {9'd67,-10'd334};
ram[20197] = {9'd70,-10'd330};
ram[20198] = {9'd73,-10'd327};
ram[20199] = {9'd76,-10'd324};
ram[20200] = {9'd80,-10'd321};
ram[20201] = {9'd83,-10'd318};
ram[20202] = {9'd86,-10'd315};
ram[20203] = {9'd89,-10'd312};
ram[20204] = {9'd92,-10'd308};
ram[20205] = {9'd95,-10'd305};
ram[20206] = {9'd98,-10'd302};
ram[20207] = {-9'd99,-10'd299};
ram[20208] = {-9'd96,-10'd296};
ram[20209] = {-9'd92,-10'd293};
ram[20210] = {-9'd89,-10'd290};
ram[20211] = {-9'd86,-10'd286};
ram[20212] = {-9'd83,-10'd283};
ram[20213] = {-9'd80,-10'd280};
ram[20214] = {-9'd77,-10'd277};
ram[20215] = {-9'd74,-10'd274};
ram[20216] = {-9'd70,-10'd271};
ram[20217] = {-9'd67,-10'd268};
ram[20218] = {-9'd64,-10'd264};
ram[20219] = {-9'd61,-10'd261};
ram[20220] = {-9'd58,-10'd258};
ram[20221] = {-9'd55,-10'd255};
ram[20222] = {-9'd52,-10'd252};
ram[20223] = {-9'd48,-10'd249};
ram[20224] = {-9'd48,-10'd249};
ram[20225] = {-9'd45,-10'd246};
ram[20226] = {-9'd42,-10'd242};
ram[20227] = {-9'd39,-10'd239};
ram[20228] = {-9'd36,-10'd236};
ram[20229] = {-9'd33,-10'd233};
ram[20230] = {-9'd30,-10'd230};
ram[20231] = {-9'd26,-10'd227};
ram[20232] = {-9'd23,-10'd224};
ram[20233] = {-9'd20,-10'd220};
ram[20234] = {-9'd17,-10'd217};
ram[20235] = {-9'd14,-10'd214};
ram[20236] = {-9'd11,-10'd211};
ram[20237] = {-9'd8,-10'd208};
ram[20238] = {-9'd4,-10'd205};
ram[20239] = {-9'd1,-10'd202};
ram[20240] = {9'd2,-10'd198};
ram[20241] = {9'd5,-10'd195};
ram[20242] = {9'd8,-10'd192};
ram[20243] = {9'd11,-10'd189};
ram[20244] = {9'd14,-10'd186};
ram[20245] = {9'd18,-10'd183};
ram[20246] = {9'd21,-10'd180};
ram[20247] = {9'd24,-10'd176};
ram[20248] = {9'd27,-10'd173};
ram[20249] = {9'd30,-10'd170};
ram[20250] = {9'd33,-10'd167};
ram[20251] = {9'd36,-10'd164};
ram[20252] = {9'd40,-10'd161};
ram[20253] = {9'd43,-10'd158};
ram[20254] = {9'd46,-10'd154};
ram[20255] = {9'd49,-10'd151};
ram[20256] = {9'd52,-10'd148};
ram[20257] = {9'd55,-10'd145};
ram[20258] = {9'd58,-10'd142};
ram[20259] = {9'd62,-10'd139};
ram[20260] = {9'd65,-10'd136};
ram[20261] = {9'd68,-10'd132};
ram[20262] = {9'd71,-10'd129};
ram[20263] = {9'd74,-10'd126};
ram[20264] = {9'd77,-10'd123};
ram[20265] = {9'd80,-10'd120};
ram[20266] = {9'd84,-10'd117};
ram[20267] = {9'd87,-10'd114};
ram[20268] = {9'd90,-10'd110};
ram[20269] = {9'd93,-10'd107};
ram[20270] = {9'd96,-10'd104};
ram[20271] = {9'd99,-10'd101};
ram[20272] = {-9'd98,-10'd98};
ram[20273] = {-9'd95,-10'd95};
ram[20274] = {-9'd92,-10'd92};
ram[20275] = {-9'd88,-10'd88};
ram[20276] = {-9'd85,-10'd85};
ram[20277] = {-9'd82,-10'd82};
ram[20278] = {-9'd79,-10'd79};
ram[20279] = {-9'd76,-10'd76};
ram[20280] = {-9'd73,-10'd73};
ram[20281] = {-9'd70,-10'd70};
ram[20282] = {-9'd66,-10'd66};
ram[20283] = {-9'd63,-10'd63};
ram[20284] = {-9'd60,-10'd60};
ram[20285] = {-9'd57,-10'd57};
ram[20286] = {-9'd54,-10'd54};
ram[20287] = {-9'd51,-10'd51};
ram[20288] = {-9'd48,-10'd48};
ram[20289] = {-9'd44,-10'd44};
ram[20290] = {-9'd41,-10'd41};
ram[20291] = {-9'd38,-10'd38};
ram[20292] = {-9'd35,-10'd35};
ram[20293] = {-9'd32,-10'd32};
ram[20294] = {-9'd29,-10'd29};
ram[20295] = {-9'd26,-10'd26};
ram[20296] = {-9'd22,-10'd22};
ram[20297] = {-9'd19,-10'd19};
ram[20298] = {-9'd16,-10'd16};
ram[20299] = {-9'd13,-10'd13};
ram[20300] = {-9'd10,-10'd10};
ram[20301] = {-9'd7,-10'd7};
ram[20302] = {-9'd4,-10'd4};
ram[20303] = {9'd0,10'd0};
ram[20304] = {9'd3,10'd3};
ram[20305] = {9'd6,10'd6};
ram[20306] = {9'd9,10'd9};
ram[20307] = {9'd12,10'd12};
ram[20308] = {9'd15,10'd15};
ram[20309] = {9'd18,10'd18};
ram[20310] = {9'd21,10'd21};
ram[20311] = {9'd25,10'd25};
ram[20312] = {9'd28,10'd28};
ram[20313] = {9'd31,10'd31};
ram[20314] = {9'd34,10'd34};
ram[20315] = {9'd37,10'd37};
ram[20316] = {9'd40,10'd40};
ram[20317] = {9'd43,10'd43};
ram[20318] = {9'd47,10'd47};
ram[20319] = {9'd50,10'd50};
ram[20320] = {9'd53,10'd53};
ram[20321] = {9'd56,10'd56};
ram[20322] = {9'd59,10'd59};
ram[20323] = {9'd62,10'd62};
ram[20324] = {9'd65,10'd65};
ram[20325] = {9'd69,10'd69};
ram[20326] = {9'd72,10'd72};
ram[20327] = {9'd75,10'd75};
ram[20328] = {9'd78,10'd78};
ram[20329] = {9'd81,10'd81};
ram[20330] = {9'd84,10'd84};
ram[20331] = {9'd87,10'd87};
ram[20332] = {9'd91,10'd91};
ram[20333] = {9'd94,10'd94};
ram[20334] = {9'd97,10'd97};
ram[20335] = {-9'd100,10'd100};
ram[20336] = {-9'd97,10'd103};
ram[20337] = {-9'd94,10'd106};
ram[20338] = {-9'd91,10'd109};
ram[20339] = {-9'd88,10'd113};
ram[20340] = {-9'd85,10'd116};
ram[20341] = {-9'd81,10'd119};
ram[20342] = {-9'd78,10'd122};
ram[20343] = {-9'd75,10'd125};
ram[20344] = {-9'd72,10'd128};
ram[20345] = {-9'd69,10'd131};
ram[20346] = {-9'd66,10'd135};
ram[20347] = {-9'd63,10'd138};
ram[20348] = {-9'd59,10'd141};
ram[20349] = {-9'd56,10'd144};
ram[20350] = {-9'd53,10'd147};
ram[20351] = {-9'd50,10'd150};
ram[20352] = {-9'd50,10'd150};
ram[20353] = {-9'd47,10'd153};
ram[20354] = {-9'd44,10'd157};
ram[20355] = {-9'd41,10'd160};
ram[20356] = {-9'd37,10'd163};
ram[20357] = {-9'd34,10'd166};
ram[20358] = {-9'd31,10'd169};
ram[20359] = {-9'd28,10'd172};
ram[20360] = {-9'd25,10'd175};
ram[20361] = {-9'd22,10'd179};
ram[20362] = {-9'd19,10'd182};
ram[20363] = {-9'd15,10'd185};
ram[20364] = {-9'd12,10'd188};
ram[20365] = {-9'd9,10'd191};
ram[20366] = {-9'd6,10'd194};
ram[20367] = {-9'd3,10'd197};
ram[20368] = {9'd0,10'd201};
ram[20369] = {9'd3,10'd204};
ram[20370] = {9'd7,10'd207};
ram[20371] = {9'd10,10'd210};
ram[20372] = {9'd13,10'd213};
ram[20373] = {9'd16,10'd216};
ram[20374] = {9'd19,10'd219};
ram[20375] = {9'd22,10'd223};
ram[20376] = {9'd25,10'd226};
ram[20377] = {9'd29,10'd229};
ram[20378] = {9'd32,10'd232};
ram[20379] = {9'd35,10'd235};
ram[20380] = {9'd38,10'd238};
ram[20381] = {9'd41,10'd241};
ram[20382] = {9'd44,10'd245};
ram[20383] = {9'd47,10'd248};
ram[20384] = {9'd51,10'd251};
ram[20385] = {9'd54,10'd254};
ram[20386] = {9'd57,10'd257};
ram[20387] = {9'd60,10'd260};
ram[20388] = {9'd63,10'd263};
ram[20389] = {9'd66,10'd267};
ram[20390] = {9'd69,10'd270};
ram[20391] = {9'd73,10'd273};
ram[20392] = {9'd76,10'd276};
ram[20393] = {9'd79,10'd279};
ram[20394] = {9'd82,10'd282};
ram[20395] = {9'd85,10'd285};
ram[20396] = {9'd88,10'd289};
ram[20397] = {9'd91,10'd292};
ram[20398] = {9'd95,10'd295};
ram[20399] = {9'd98,10'd298};
ram[20400] = {-9'd99,10'd301};
ram[20401] = {-9'd96,10'd304};
ram[20402] = {-9'd93,10'd307};
ram[20403] = {-9'd90,10'd311};
ram[20404] = {-9'd87,10'd314};
ram[20405] = {-9'd84,10'd317};
ram[20406] = {-9'd81,10'd320};
ram[20407] = {-9'd77,10'd323};
ram[20408] = {-9'd74,10'd326};
ram[20409] = {-9'd71,10'd329};
ram[20410] = {-9'd68,10'd333};
ram[20411] = {-9'd65,10'd336};
ram[20412] = {-9'd62,10'd339};
ram[20413] = {-9'd59,10'd342};
ram[20414] = {-9'd55,10'd345};
ram[20415] = {-9'd52,10'd348};
ram[20416] = {-9'd49,10'd351};
ram[20417] = {-9'd46,10'd354};
ram[20418] = {-9'd43,10'd358};
ram[20419] = {-9'd40,10'd361};
ram[20420] = {-9'd37,10'd364};
ram[20421] = {-9'd33,10'd367};
ram[20422] = {-9'd30,10'd370};
ram[20423] = {-9'd27,10'd373};
ram[20424] = {-9'd24,10'd376};
ram[20425] = {-9'd21,10'd380};
ram[20426] = {-9'd18,10'd383};
ram[20427] = {-9'd15,10'd386};
ram[20428] = {-9'd11,10'd389};
ram[20429] = {-9'd8,10'd392};
ram[20430] = {-9'd5,10'd395};
ram[20431] = {-9'd2,10'd398};
ram[20432] = {9'd1,-10'd399};
ram[20433] = {9'd4,-10'd396};
ram[20434] = {9'd7,-10'd393};
ram[20435] = {9'd10,-10'd390};
ram[20436] = {9'd14,-10'd387};
ram[20437] = {9'd17,-10'd384};
ram[20438] = {9'd20,-10'd381};
ram[20439] = {9'd23,-10'd377};
ram[20440] = {9'd26,-10'd374};
ram[20441] = {9'd29,-10'd371};
ram[20442] = {9'd32,-10'd368};
ram[20443] = {9'd36,-10'd365};
ram[20444] = {9'd39,-10'd362};
ram[20445] = {9'd42,-10'd359};
ram[20446] = {9'd45,-10'd355};
ram[20447] = {9'd48,-10'd352};
ram[20448] = {9'd51,-10'd349};
ram[20449] = {9'd54,-10'd346};
ram[20450] = {9'd58,-10'd343};
ram[20451] = {9'd61,-10'd340};
ram[20452] = {9'd64,-10'd337};
ram[20453] = {9'd67,-10'd334};
ram[20454] = {9'd70,-10'd330};
ram[20455] = {9'd73,-10'd327};
ram[20456] = {9'd76,-10'd324};
ram[20457] = {9'd80,-10'd321};
ram[20458] = {9'd83,-10'd318};
ram[20459] = {9'd86,-10'd315};
ram[20460] = {9'd89,-10'd312};
ram[20461] = {9'd92,-10'd308};
ram[20462] = {9'd95,-10'd305};
ram[20463] = {9'd98,-10'd302};
ram[20464] = {-9'd99,-10'd299};
ram[20465] = {-9'd96,-10'd296};
ram[20466] = {-9'd92,-10'd293};
ram[20467] = {-9'd89,-10'd290};
ram[20468] = {-9'd86,-10'd286};
ram[20469] = {-9'd83,-10'd283};
ram[20470] = {-9'd80,-10'd280};
ram[20471] = {-9'd77,-10'd277};
ram[20472] = {-9'd74,-10'd274};
ram[20473] = {-9'd70,-10'd271};
ram[20474] = {-9'd67,-10'd268};
ram[20475] = {-9'd64,-10'd264};
ram[20476] = {-9'd61,-10'd261};
ram[20477] = {-9'd58,-10'd258};
ram[20478] = {-9'd55,-10'd255};
ram[20479] = {-9'd52,-10'd252};
ram[20480] = {-9'd52,-10'd252};
ram[20481] = {-9'd48,-10'd249};
ram[20482] = {-9'd45,-10'd246};
ram[20483] = {-9'd42,-10'd242};
ram[20484] = {-9'd39,-10'd239};
ram[20485] = {-9'd36,-10'd236};
ram[20486] = {-9'd33,-10'd233};
ram[20487] = {-9'd30,-10'd230};
ram[20488] = {-9'd26,-10'd227};
ram[20489] = {-9'd23,-10'd224};
ram[20490] = {-9'd20,-10'd220};
ram[20491] = {-9'd17,-10'd217};
ram[20492] = {-9'd14,-10'd214};
ram[20493] = {-9'd11,-10'd211};
ram[20494] = {-9'd8,-10'd208};
ram[20495] = {-9'd4,-10'd205};
ram[20496] = {-9'd1,-10'd202};
ram[20497] = {9'd2,-10'd198};
ram[20498] = {9'd5,-10'd195};
ram[20499] = {9'd8,-10'd192};
ram[20500] = {9'd11,-10'd189};
ram[20501] = {9'd14,-10'd186};
ram[20502] = {9'd18,-10'd183};
ram[20503] = {9'd21,-10'd180};
ram[20504] = {9'd24,-10'd176};
ram[20505] = {9'd27,-10'd173};
ram[20506] = {9'd30,-10'd170};
ram[20507] = {9'd33,-10'd167};
ram[20508] = {9'd36,-10'd164};
ram[20509] = {9'd40,-10'd161};
ram[20510] = {9'd43,-10'd158};
ram[20511] = {9'd46,-10'd154};
ram[20512] = {9'd49,-10'd151};
ram[20513] = {9'd52,-10'd148};
ram[20514] = {9'd55,-10'd145};
ram[20515] = {9'd58,-10'd142};
ram[20516] = {9'd62,-10'd139};
ram[20517] = {9'd65,-10'd136};
ram[20518] = {9'd68,-10'd132};
ram[20519] = {9'd71,-10'd129};
ram[20520] = {9'd74,-10'd126};
ram[20521] = {9'd77,-10'd123};
ram[20522] = {9'd80,-10'd120};
ram[20523] = {9'd84,-10'd117};
ram[20524] = {9'd87,-10'd114};
ram[20525] = {9'd90,-10'd110};
ram[20526] = {9'd93,-10'd107};
ram[20527] = {9'd96,-10'd104};
ram[20528] = {9'd99,-10'd101};
ram[20529] = {-9'd98,-10'd98};
ram[20530] = {-9'd95,-10'd95};
ram[20531] = {-9'd92,-10'd92};
ram[20532] = {-9'd88,-10'd88};
ram[20533] = {-9'd85,-10'd85};
ram[20534] = {-9'd82,-10'd82};
ram[20535] = {-9'd79,-10'd79};
ram[20536] = {-9'd76,-10'd76};
ram[20537] = {-9'd73,-10'd73};
ram[20538] = {-9'd70,-10'd70};
ram[20539] = {-9'd66,-10'd66};
ram[20540] = {-9'd63,-10'd63};
ram[20541] = {-9'd60,-10'd60};
ram[20542] = {-9'd57,-10'd57};
ram[20543] = {-9'd54,-10'd54};
ram[20544] = {-9'd51,-10'd51};
ram[20545] = {-9'd48,-10'd48};
ram[20546] = {-9'd44,-10'd44};
ram[20547] = {-9'd41,-10'd41};
ram[20548] = {-9'd38,-10'd38};
ram[20549] = {-9'd35,-10'd35};
ram[20550] = {-9'd32,-10'd32};
ram[20551] = {-9'd29,-10'd29};
ram[20552] = {-9'd26,-10'd26};
ram[20553] = {-9'd22,-10'd22};
ram[20554] = {-9'd19,-10'd19};
ram[20555] = {-9'd16,-10'd16};
ram[20556] = {-9'd13,-10'd13};
ram[20557] = {-9'd10,-10'd10};
ram[20558] = {-9'd7,-10'd7};
ram[20559] = {-9'd4,-10'd4};
ram[20560] = {9'd0,10'd0};
ram[20561] = {9'd3,10'd3};
ram[20562] = {9'd6,10'd6};
ram[20563] = {9'd9,10'd9};
ram[20564] = {9'd12,10'd12};
ram[20565] = {9'd15,10'd15};
ram[20566] = {9'd18,10'd18};
ram[20567] = {9'd21,10'd21};
ram[20568] = {9'd25,10'd25};
ram[20569] = {9'd28,10'd28};
ram[20570] = {9'd31,10'd31};
ram[20571] = {9'd34,10'd34};
ram[20572] = {9'd37,10'd37};
ram[20573] = {9'd40,10'd40};
ram[20574] = {9'd43,10'd43};
ram[20575] = {9'd47,10'd47};
ram[20576] = {9'd50,10'd50};
ram[20577] = {9'd53,10'd53};
ram[20578] = {9'd56,10'd56};
ram[20579] = {9'd59,10'd59};
ram[20580] = {9'd62,10'd62};
ram[20581] = {9'd65,10'd65};
ram[20582] = {9'd69,10'd69};
ram[20583] = {9'd72,10'd72};
ram[20584] = {9'd75,10'd75};
ram[20585] = {9'd78,10'd78};
ram[20586] = {9'd81,10'd81};
ram[20587] = {9'd84,10'd84};
ram[20588] = {9'd87,10'd87};
ram[20589] = {9'd91,10'd91};
ram[20590] = {9'd94,10'd94};
ram[20591] = {9'd97,10'd97};
ram[20592] = {-9'd100,10'd100};
ram[20593] = {-9'd97,10'd103};
ram[20594] = {-9'd94,10'd106};
ram[20595] = {-9'd91,10'd109};
ram[20596] = {-9'd88,10'd113};
ram[20597] = {-9'd85,10'd116};
ram[20598] = {-9'd81,10'd119};
ram[20599] = {-9'd78,10'd122};
ram[20600] = {-9'd75,10'd125};
ram[20601] = {-9'd72,10'd128};
ram[20602] = {-9'd69,10'd131};
ram[20603] = {-9'd66,10'd135};
ram[20604] = {-9'd63,10'd138};
ram[20605] = {-9'd59,10'd141};
ram[20606] = {-9'd56,10'd144};
ram[20607] = {-9'd53,10'd147};
ram[20608] = {-9'd53,10'd147};
ram[20609] = {-9'd50,10'd150};
ram[20610] = {-9'd47,10'd153};
ram[20611] = {-9'd44,10'd157};
ram[20612] = {-9'd41,10'd160};
ram[20613] = {-9'd37,10'd163};
ram[20614] = {-9'd34,10'd166};
ram[20615] = {-9'd31,10'd169};
ram[20616] = {-9'd28,10'd172};
ram[20617] = {-9'd25,10'd175};
ram[20618] = {-9'd22,10'd179};
ram[20619] = {-9'd19,10'd182};
ram[20620] = {-9'd15,10'd185};
ram[20621] = {-9'd12,10'd188};
ram[20622] = {-9'd9,10'd191};
ram[20623] = {-9'd6,10'd194};
ram[20624] = {-9'd3,10'd197};
ram[20625] = {9'd0,10'd201};
ram[20626] = {9'd3,10'd204};
ram[20627] = {9'd7,10'd207};
ram[20628] = {9'd10,10'd210};
ram[20629] = {9'd13,10'd213};
ram[20630] = {9'd16,10'd216};
ram[20631] = {9'd19,10'd219};
ram[20632] = {9'd22,10'd223};
ram[20633] = {9'd25,10'd226};
ram[20634] = {9'd29,10'd229};
ram[20635] = {9'd32,10'd232};
ram[20636] = {9'd35,10'd235};
ram[20637] = {9'd38,10'd238};
ram[20638] = {9'd41,10'd241};
ram[20639] = {9'd44,10'd245};
ram[20640] = {9'd47,10'd248};
ram[20641] = {9'd51,10'd251};
ram[20642] = {9'd54,10'd254};
ram[20643] = {9'd57,10'd257};
ram[20644] = {9'd60,10'd260};
ram[20645] = {9'd63,10'd263};
ram[20646] = {9'd66,10'd267};
ram[20647] = {9'd69,10'd270};
ram[20648] = {9'd73,10'd273};
ram[20649] = {9'd76,10'd276};
ram[20650] = {9'd79,10'd279};
ram[20651] = {9'd82,10'd282};
ram[20652] = {9'd85,10'd285};
ram[20653] = {9'd88,10'd289};
ram[20654] = {9'd91,10'd292};
ram[20655] = {9'd95,10'd295};
ram[20656] = {9'd98,10'd298};
ram[20657] = {-9'd99,10'd301};
ram[20658] = {-9'd96,10'd304};
ram[20659] = {-9'd93,10'd307};
ram[20660] = {-9'd90,10'd311};
ram[20661] = {-9'd87,10'd314};
ram[20662] = {-9'd84,10'd317};
ram[20663] = {-9'd81,10'd320};
ram[20664] = {-9'd77,10'd323};
ram[20665] = {-9'd74,10'd326};
ram[20666] = {-9'd71,10'd329};
ram[20667] = {-9'd68,10'd333};
ram[20668] = {-9'd65,10'd336};
ram[20669] = {-9'd62,10'd339};
ram[20670] = {-9'd59,10'd342};
ram[20671] = {-9'd55,10'd345};
ram[20672] = {-9'd52,10'd348};
ram[20673] = {-9'd49,10'd351};
ram[20674] = {-9'd46,10'd354};
ram[20675] = {-9'd43,10'd358};
ram[20676] = {-9'd40,10'd361};
ram[20677] = {-9'd37,10'd364};
ram[20678] = {-9'd33,10'd367};
ram[20679] = {-9'd30,10'd370};
ram[20680] = {-9'd27,10'd373};
ram[20681] = {-9'd24,10'd376};
ram[20682] = {-9'd21,10'd380};
ram[20683] = {-9'd18,10'd383};
ram[20684] = {-9'd15,10'd386};
ram[20685] = {-9'd11,10'd389};
ram[20686] = {-9'd8,10'd392};
ram[20687] = {-9'd5,10'd395};
ram[20688] = {-9'd2,10'd398};
ram[20689] = {9'd1,-10'd399};
ram[20690] = {9'd4,-10'd396};
ram[20691] = {9'd7,-10'd393};
ram[20692] = {9'd10,-10'd390};
ram[20693] = {9'd14,-10'd387};
ram[20694] = {9'd17,-10'd384};
ram[20695] = {9'd20,-10'd381};
ram[20696] = {9'd23,-10'd377};
ram[20697] = {9'd26,-10'd374};
ram[20698] = {9'd29,-10'd371};
ram[20699] = {9'd32,-10'd368};
ram[20700] = {9'd36,-10'd365};
ram[20701] = {9'd39,-10'd362};
ram[20702] = {9'd42,-10'd359};
ram[20703] = {9'd45,-10'd355};
ram[20704] = {9'd48,-10'd352};
ram[20705] = {9'd51,-10'd349};
ram[20706] = {9'd54,-10'd346};
ram[20707] = {9'd58,-10'd343};
ram[20708] = {9'd61,-10'd340};
ram[20709] = {9'd64,-10'd337};
ram[20710] = {9'd67,-10'd334};
ram[20711] = {9'd70,-10'd330};
ram[20712] = {9'd73,-10'd327};
ram[20713] = {9'd76,-10'd324};
ram[20714] = {9'd80,-10'd321};
ram[20715] = {9'd83,-10'd318};
ram[20716] = {9'd86,-10'd315};
ram[20717] = {9'd89,-10'd312};
ram[20718] = {9'd92,-10'd308};
ram[20719] = {9'd95,-10'd305};
ram[20720] = {9'd98,-10'd302};
ram[20721] = {-9'd99,-10'd299};
ram[20722] = {-9'd96,-10'd296};
ram[20723] = {-9'd92,-10'd293};
ram[20724] = {-9'd89,-10'd290};
ram[20725] = {-9'd86,-10'd286};
ram[20726] = {-9'd83,-10'd283};
ram[20727] = {-9'd80,-10'd280};
ram[20728] = {-9'd77,-10'd277};
ram[20729] = {-9'd74,-10'd274};
ram[20730] = {-9'd70,-10'd271};
ram[20731] = {-9'd67,-10'd268};
ram[20732] = {-9'd64,-10'd264};
ram[20733] = {-9'd61,-10'd261};
ram[20734] = {-9'd58,-10'd258};
ram[20735] = {-9'd55,-10'd255};
ram[20736] = {-9'd55,-10'd255};
ram[20737] = {-9'd52,-10'd252};
ram[20738] = {-9'd48,-10'd249};
ram[20739] = {-9'd45,-10'd246};
ram[20740] = {-9'd42,-10'd242};
ram[20741] = {-9'd39,-10'd239};
ram[20742] = {-9'd36,-10'd236};
ram[20743] = {-9'd33,-10'd233};
ram[20744] = {-9'd30,-10'd230};
ram[20745] = {-9'd26,-10'd227};
ram[20746] = {-9'd23,-10'd224};
ram[20747] = {-9'd20,-10'd220};
ram[20748] = {-9'd17,-10'd217};
ram[20749] = {-9'd14,-10'd214};
ram[20750] = {-9'd11,-10'd211};
ram[20751] = {-9'd8,-10'd208};
ram[20752] = {-9'd4,-10'd205};
ram[20753] = {-9'd1,-10'd202};
ram[20754] = {9'd2,-10'd198};
ram[20755] = {9'd5,-10'd195};
ram[20756] = {9'd8,-10'd192};
ram[20757] = {9'd11,-10'd189};
ram[20758] = {9'd14,-10'd186};
ram[20759] = {9'd18,-10'd183};
ram[20760] = {9'd21,-10'd180};
ram[20761] = {9'd24,-10'd176};
ram[20762] = {9'd27,-10'd173};
ram[20763] = {9'd30,-10'd170};
ram[20764] = {9'd33,-10'd167};
ram[20765] = {9'd36,-10'd164};
ram[20766] = {9'd40,-10'd161};
ram[20767] = {9'd43,-10'd158};
ram[20768] = {9'd46,-10'd154};
ram[20769] = {9'd49,-10'd151};
ram[20770] = {9'd52,-10'd148};
ram[20771] = {9'd55,-10'd145};
ram[20772] = {9'd58,-10'd142};
ram[20773] = {9'd62,-10'd139};
ram[20774] = {9'd65,-10'd136};
ram[20775] = {9'd68,-10'd132};
ram[20776] = {9'd71,-10'd129};
ram[20777] = {9'd74,-10'd126};
ram[20778] = {9'd77,-10'd123};
ram[20779] = {9'd80,-10'd120};
ram[20780] = {9'd84,-10'd117};
ram[20781] = {9'd87,-10'd114};
ram[20782] = {9'd90,-10'd110};
ram[20783] = {9'd93,-10'd107};
ram[20784] = {9'd96,-10'd104};
ram[20785] = {9'd99,-10'd101};
ram[20786] = {-9'd98,-10'd98};
ram[20787] = {-9'd95,-10'd95};
ram[20788] = {-9'd92,-10'd92};
ram[20789] = {-9'd88,-10'd88};
ram[20790] = {-9'd85,-10'd85};
ram[20791] = {-9'd82,-10'd82};
ram[20792] = {-9'd79,-10'd79};
ram[20793] = {-9'd76,-10'd76};
ram[20794] = {-9'd73,-10'd73};
ram[20795] = {-9'd70,-10'd70};
ram[20796] = {-9'd66,-10'd66};
ram[20797] = {-9'd63,-10'd63};
ram[20798] = {-9'd60,-10'd60};
ram[20799] = {-9'd57,-10'd57};
ram[20800] = {-9'd54,-10'd54};
ram[20801] = {-9'd51,-10'd51};
ram[20802] = {-9'd48,-10'd48};
ram[20803] = {-9'd44,-10'd44};
ram[20804] = {-9'd41,-10'd41};
ram[20805] = {-9'd38,-10'd38};
ram[20806] = {-9'd35,-10'd35};
ram[20807] = {-9'd32,-10'd32};
ram[20808] = {-9'd29,-10'd29};
ram[20809] = {-9'd26,-10'd26};
ram[20810] = {-9'd22,-10'd22};
ram[20811] = {-9'd19,-10'd19};
ram[20812] = {-9'd16,-10'd16};
ram[20813] = {-9'd13,-10'd13};
ram[20814] = {-9'd10,-10'd10};
ram[20815] = {-9'd7,-10'd7};
ram[20816] = {-9'd4,-10'd4};
ram[20817] = {9'd0,10'd0};
ram[20818] = {9'd3,10'd3};
ram[20819] = {9'd6,10'd6};
ram[20820] = {9'd9,10'd9};
ram[20821] = {9'd12,10'd12};
ram[20822] = {9'd15,10'd15};
ram[20823] = {9'd18,10'd18};
ram[20824] = {9'd21,10'd21};
ram[20825] = {9'd25,10'd25};
ram[20826] = {9'd28,10'd28};
ram[20827] = {9'd31,10'd31};
ram[20828] = {9'd34,10'd34};
ram[20829] = {9'd37,10'd37};
ram[20830] = {9'd40,10'd40};
ram[20831] = {9'd43,10'd43};
ram[20832] = {9'd47,10'd47};
ram[20833] = {9'd50,10'd50};
ram[20834] = {9'd53,10'd53};
ram[20835] = {9'd56,10'd56};
ram[20836] = {9'd59,10'd59};
ram[20837] = {9'd62,10'd62};
ram[20838] = {9'd65,10'd65};
ram[20839] = {9'd69,10'd69};
ram[20840] = {9'd72,10'd72};
ram[20841] = {9'd75,10'd75};
ram[20842] = {9'd78,10'd78};
ram[20843] = {9'd81,10'd81};
ram[20844] = {9'd84,10'd84};
ram[20845] = {9'd87,10'd87};
ram[20846] = {9'd91,10'd91};
ram[20847] = {9'd94,10'd94};
ram[20848] = {9'd97,10'd97};
ram[20849] = {-9'd100,10'd100};
ram[20850] = {-9'd97,10'd103};
ram[20851] = {-9'd94,10'd106};
ram[20852] = {-9'd91,10'd109};
ram[20853] = {-9'd88,10'd113};
ram[20854] = {-9'd85,10'd116};
ram[20855] = {-9'd81,10'd119};
ram[20856] = {-9'd78,10'd122};
ram[20857] = {-9'd75,10'd125};
ram[20858] = {-9'd72,10'd128};
ram[20859] = {-9'd69,10'd131};
ram[20860] = {-9'd66,10'd135};
ram[20861] = {-9'd63,10'd138};
ram[20862] = {-9'd59,10'd141};
ram[20863] = {-9'd56,10'd144};
ram[20864] = {-9'd56,10'd144};
ram[20865] = {-9'd53,10'd147};
ram[20866] = {-9'd50,10'd150};
ram[20867] = {-9'd47,10'd153};
ram[20868] = {-9'd44,10'd157};
ram[20869] = {-9'd41,10'd160};
ram[20870] = {-9'd37,10'd163};
ram[20871] = {-9'd34,10'd166};
ram[20872] = {-9'd31,10'd169};
ram[20873] = {-9'd28,10'd172};
ram[20874] = {-9'd25,10'd175};
ram[20875] = {-9'd22,10'd179};
ram[20876] = {-9'd19,10'd182};
ram[20877] = {-9'd15,10'd185};
ram[20878] = {-9'd12,10'd188};
ram[20879] = {-9'd9,10'd191};
ram[20880] = {-9'd6,10'd194};
ram[20881] = {-9'd3,10'd197};
ram[20882] = {9'd0,10'd201};
ram[20883] = {9'd3,10'd204};
ram[20884] = {9'd7,10'd207};
ram[20885] = {9'd10,10'd210};
ram[20886] = {9'd13,10'd213};
ram[20887] = {9'd16,10'd216};
ram[20888] = {9'd19,10'd219};
ram[20889] = {9'd22,10'd223};
ram[20890] = {9'd25,10'd226};
ram[20891] = {9'd29,10'd229};
ram[20892] = {9'd32,10'd232};
ram[20893] = {9'd35,10'd235};
ram[20894] = {9'd38,10'd238};
ram[20895] = {9'd41,10'd241};
ram[20896] = {9'd44,10'd245};
ram[20897] = {9'd47,10'd248};
ram[20898] = {9'd51,10'd251};
ram[20899] = {9'd54,10'd254};
ram[20900] = {9'd57,10'd257};
ram[20901] = {9'd60,10'd260};
ram[20902] = {9'd63,10'd263};
ram[20903] = {9'd66,10'd267};
ram[20904] = {9'd69,10'd270};
ram[20905] = {9'd73,10'd273};
ram[20906] = {9'd76,10'd276};
ram[20907] = {9'd79,10'd279};
ram[20908] = {9'd82,10'd282};
ram[20909] = {9'd85,10'd285};
ram[20910] = {9'd88,10'd289};
ram[20911] = {9'd91,10'd292};
ram[20912] = {9'd95,10'd295};
ram[20913] = {9'd98,10'd298};
ram[20914] = {-9'd99,10'd301};
ram[20915] = {-9'd96,10'd304};
ram[20916] = {-9'd93,10'd307};
ram[20917] = {-9'd90,10'd311};
ram[20918] = {-9'd87,10'd314};
ram[20919] = {-9'd84,10'd317};
ram[20920] = {-9'd81,10'd320};
ram[20921] = {-9'd77,10'd323};
ram[20922] = {-9'd74,10'd326};
ram[20923] = {-9'd71,10'd329};
ram[20924] = {-9'd68,10'd333};
ram[20925] = {-9'd65,10'd336};
ram[20926] = {-9'd62,10'd339};
ram[20927] = {-9'd59,10'd342};
ram[20928] = {-9'd55,10'd345};
ram[20929] = {-9'd52,10'd348};
ram[20930] = {-9'd49,10'd351};
ram[20931] = {-9'd46,10'd354};
ram[20932] = {-9'd43,10'd358};
ram[20933] = {-9'd40,10'd361};
ram[20934] = {-9'd37,10'd364};
ram[20935] = {-9'd33,10'd367};
ram[20936] = {-9'd30,10'd370};
ram[20937] = {-9'd27,10'd373};
ram[20938] = {-9'd24,10'd376};
ram[20939] = {-9'd21,10'd380};
ram[20940] = {-9'd18,10'd383};
ram[20941] = {-9'd15,10'd386};
ram[20942] = {-9'd11,10'd389};
ram[20943] = {-9'd8,10'd392};
ram[20944] = {-9'd5,10'd395};
ram[20945] = {-9'd2,10'd398};
ram[20946] = {9'd1,-10'd399};
ram[20947] = {9'd4,-10'd396};
ram[20948] = {9'd7,-10'd393};
ram[20949] = {9'd10,-10'd390};
ram[20950] = {9'd14,-10'd387};
ram[20951] = {9'd17,-10'd384};
ram[20952] = {9'd20,-10'd381};
ram[20953] = {9'd23,-10'd377};
ram[20954] = {9'd26,-10'd374};
ram[20955] = {9'd29,-10'd371};
ram[20956] = {9'd32,-10'd368};
ram[20957] = {9'd36,-10'd365};
ram[20958] = {9'd39,-10'd362};
ram[20959] = {9'd42,-10'd359};
ram[20960] = {9'd45,-10'd355};
ram[20961] = {9'd48,-10'd352};
ram[20962] = {9'd51,-10'd349};
ram[20963] = {9'd54,-10'd346};
ram[20964] = {9'd58,-10'd343};
ram[20965] = {9'd61,-10'd340};
ram[20966] = {9'd64,-10'd337};
ram[20967] = {9'd67,-10'd334};
ram[20968] = {9'd70,-10'd330};
ram[20969] = {9'd73,-10'd327};
ram[20970] = {9'd76,-10'd324};
ram[20971] = {9'd80,-10'd321};
ram[20972] = {9'd83,-10'd318};
ram[20973] = {9'd86,-10'd315};
ram[20974] = {9'd89,-10'd312};
ram[20975] = {9'd92,-10'd308};
ram[20976] = {9'd95,-10'd305};
ram[20977] = {9'd98,-10'd302};
ram[20978] = {-9'd99,-10'd299};
ram[20979] = {-9'd96,-10'd296};
ram[20980] = {-9'd92,-10'd293};
ram[20981] = {-9'd89,-10'd290};
ram[20982] = {-9'd86,-10'd286};
ram[20983] = {-9'd83,-10'd283};
ram[20984] = {-9'd80,-10'd280};
ram[20985] = {-9'd77,-10'd277};
ram[20986] = {-9'd74,-10'd274};
ram[20987] = {-9'd70,-10'd271};
ram[20988] = {-9'd67,-10'd268};
ram[20989] = {-9'd64,-10'd264};
ram[20990] = {-9'd61,-10'd261};
ram[20991] = {-9'd58,-10'd258};
ram[20992] = {-9'd58,-10'd258};
ram[20993] = {-9'd55,-10'd255};
ram[20994] = {-9'd52,-10'd252};
ram[20995] = {-9'd48,-10'd249};
ram[20996] = {-9'd45,-10'd246};
ram[20997] = {-9'd42,-10'd242};
ram[20998] = {-9'd39,-10'd239};
ram[20999] = {-9'd36,-10'd236};
ram[21000] = {-9'd33,-10'd233};
ram[21001] = {-9'd30,-10'd230};
ram[21002] = {-9'd26,-10'd227};
ram[21003] = {-9'd23,-10'd224};
ram[21004] = {-9'd20,-10'd220};
ram[21005] = {-9'd17,-10'd217};
ram[21006] = {-9'd14,-10'd214};
ram[21007] = {-9'd11,-10'd211};
ram[21008] = {-9'd8,-10'd208};
ram[21009] = {-9'd4,-10'd205};
ram[21010] = {-9'd1,-10'd202};
ram[21011] = {9'd2,-10'd198};
ram[21012] = {9'd5,-10'd195};
ram[21013] = {9'd8,-10'd192};
ram[21014] = {9'd11,-10'd189};
ram[21015] = {9'd14,-10'd186};
ram[21016] = {9'd18,-10'd183};
ram[21017] = {9'd21,-10'd180};
ram[21018] = {9'd24,-10'd176};
ram[21019] = {9'd27,-10'd173};
ram[21020] = {9'd30,-10'd170};
ram[21021] = {9'd33,-10'd167};
ram[21022] = {9'd36,-10'd164};
ram[21023] = {9'd40,-10'd161};
ram[21024] = {9'd43,-10'd158};
ram[21025] = {9'd46,-10'd154};
ram[21026] = {9'd49,-10'd151};
ram[21027] = {9'd52,-10'd148};
ram[21028] = {9'd55,-10'd145};
ram[21029] = {9'd58,-10'd142};
ram[21030] = {9'd62,-10'd139};
ram[21031] = {9'd65,-10'd136};
ram[21032] = {9'd68,-10'd132};
ram[21033] = {9'd71,-10'd129};
ram[21034] = {9'd74,-10'd126};
ram[21035] = {9'd77,-10'd123};
ram[21036] = {9'd80,-10'd120};
ram[21037] = {9'd84,-10'd117};
ram[21038] = {9'd87,-10'd114};
ram[21039] = {9'd90,-10'd110};
ram[21040] = {9'd93,-10'd107};
ram[21041] = {9'd96,-10'd104};
ram[21042] = {9'd99,-10'd101};
ram[21043] = {-9'd98,-10'd98};
ram[21044] = {-9'd95,-10'd95};
ram[21045] = {-9'd92,-10'd92};
ram[21046] = {-9'd88,-10'd88};
ram[21047] = {-9'd85,-10'd85};
ram[21048] = {-9'd82,-10'd82};
ram[21049] = {-9'd79,-10'd79};
ram[21050] = {-9'd76,-10'd76};
ram[21051] = {-9'd73,-10'd73};
ram[21052] = {-9'd70,-10'd70};
ram[21053] = {-9'd66,-10'd66};
ram[21054] = {-9'd63,-10'd63};
ram[21055] = {-9'd60,-10'd60};
ram[21056] = {-9'd57,-10'd57};
ram[21057] = {-9'd54,-10'd54};
ram[21058] = {-9'd51,-10'd51};
ram[21059] = {-9'd48,-10'd48};
ram[21060] = {-9'd44,-10'd44};
ram[21061] = {-9'd41,-10'd41};
ram[21062] = {-9'd38,-10'd38};
ram[21063] = {-9'd35,-10'd35};
ram[21064] = {-9'd32,-10'd32};
ram[21065] = {-9'd29,-10'd29};
ram[21066] = {-9'd26,-10'd26};
ram[21067] = {-9'd22,-10'd22};
ram[21068] = {-9'd19,-10'd19};
ram[21069] = {-9'd16,-10'd16};
ram[21070] = {-9'd13,-10'd13};
ram[21071] = {-9'd10,-10'd10};
ram[21072] = {-9'd7,-10'd7};
ram[21073] = {-9'd4,-10'd4};
ram[21074] = {9'd0,10'd0};
ram[21075] = {9'd3,10'd3};
ram[21076] = {9'd6,10'd6};
ram[21077] = {9'd9,10'd9};
ram[21078] = {9'd12,10'd12};
ram[21079] = {9'd15,10'd15};
ram[21080] = {9'd18,10'd18};
ram[21081] = {9'd21,10'd21};
ram[21082] = {9'd25,10'd25};
ram[21083] = {9'd28,10'd28};
ram[21084] = {9'd31,10'd31};
ram[21085] = {9'd34,10'd34};
ram[21086] = {9'd37,10'd37};
ram[21087] = {9'd40,10'd40};
ram[21088] = {9'd43,10'd43};
ram[21089] = {9'd47,10'd47};
ram[21090] = {9'd50,10'd50};
ram[21091] = {9'd53,10'd53};
ram[21092] = {9'd56,10'd56};
ram[21093] = {9'd59,10'd59};
ram[21094] = {9'd62,10'd62};
ram[21095] = {9'd65,10'd65};
ram[21096] = {9'd69,10'd69};
ram[21097] = {9'd72,10'd72};
ram[21098] = {9'd75,10'd75};
ram[21099] = {9'd78,10'd78};
ram[21100] = {9'd81,10'd81};
ram[21101] = {9'd84,10'd84};
ram[21102] = {9'd87,10'd87};
ram[21103] = {9'd91,10'd91};
ram[21104] = {9'd94,10'd94};
ram[21105] = {9'd97,10'd97};
ram[21106] = {-9'd100,10'd100};
ram[21107] = {-9'd97,10'd103};
ram[21108] = {-9'd94,10'd106};
ram[21109] = {-9'd91,10'd109};
ram[21110] = {-9'd88,10'd113};
ram[21111] = {-9'd85,10'd116};
ram[21112] = {-9'd81,10'd119};
ram[21113] = {-9'd78,10'd122};
ram[21114] = {-9'd75,10'd125};
ram[21115] = {-9'd72,10'd128};
ram[21116] = {-9'd69,10'd131};
ram[21117] = {-9'd66,10'd135};
ram[21118] = {-9'd63,10'd138};
ram[21119] = {-9'd59,10'd141};
ram[21120] = {-9'd59,10'd141};
ram[21121] = {-9'd56,10'd144};
ram[21122] = {-9'd53,10'd147};
ram[21123] = {-9'd50,10'd150};
ram[21124] = {-9'd47,10'd153};
ram[21125] = {-9'd44,10'd157};
ram[21126] = {-9'd41,10'd160};
ram[21127] = {-9'd37,10'd163};
ram[21128] = {-9'd34,10'd166};
ram[21129] = {-9'd31,10'd169};
ram[21130] = {-9'd28,10'd172};
ram[21131] = {-9'd25,10'd175};
ram[21132] = {-9'd22,10'd179};
ram[21133] = {-9'd19,10'd182};
ram[21134] = {-9'd15,10'd185};
ram[21135] = {-9'd12,10'd188};
ram[21136] = {-9'd9,10'd191};
ram[21137] = {-9'd6,10'd194};
ram[21138] = {-9'd3,10'd197};
ram[21139] = {9'd0,10'd201};
ram[21140] = {9'd3,10'd204};
ram[21141] = {9'd7,10'd207};
ram[21142] = {9'd10,10'd210};
ram[21143] = {9'd13,10'd213};
ram[21144] = {9'd16,10'd216};
ram[21145] = {9'd19,10'd219};
ram[21146] = {9'd22,10'd223};
ram[21147] = {9'd25,10'd226};
ram[21148] = {9'd29,10'd229};
ram[21149] = {9'd32,10'd232};
ram[21150] = {9'd35,10'd235};
ram[21151] = {9'd38,10'd238};
ram[21152] = {9'd41,10'd241};
ram[21153] = {9'd44,10'd245};
ram[21154] = {9'd47,10'd248};
ram[21155] = {9'd51,10'd251};
ram[21156] = {9'd54,10'd254};
ram[21157] = {9'd57,10'd257};
ram[21158] = {9'd60,10'd260};
ram[21159] = {9'd63,10'd263};
ram[21160] = {9'd66,10'd267};
ram[21161] = {9'd69,10'd270};
ram[21162] = {9'd73,10'd273};
ram[21163] = {9'd76,10'd276};
ram[21164] = {9'd79,10'd279};
ram[21165] = {9'd82,10'd282};
ram[21166] = {9'd85,10'd285};
ram[21167] = {9'd88,10'd289};
ram[21168] = {9'd91,10'd292};
ram[21169] = {9'd95,10'd295};
ram[21170] = {9'd98,10'd298};
ram[21171] = {-9'd99,10'd301};
ram[21172] = {-9'd96,10'd304};
ram[21173] = {-9'd93,10'd307};
ram[21174] = {-9'd90,10'd311};
ram[21175] = {-9'd87,10'd314};
ram[21176] = {-9'd84,10'd317};
ram[21177] = {-9'd81,10'd320};
ram[21178] = {-9'd77,10'd323};
ram[21179] = {-9'd74,10'd326};
ram[21180] = {-9'd71,10'd329};
ram[21181] = {-9'd68,10'd333};
ram[21182] = {-9'd65,10'd336};
ram[21183] = {-9'd62,10'd339};
ram[21184] = {-9'd59,10'd342};
ram[21185] = {-9'd55,10'd345};
ram[21186] = {-9'd52,10'd348};
ram[21187] = {-9'd49,10'd351};
ram[21188] = {-9'd46,10'd354};
ram[21189] = {-9'd43,10'd358};
ram[21190] = {-9'd40,10'd361};
ram[21191] = {-9'd37,10'd364};
ram[21192] = {-9'd33,10'd367};
ram[21193] = {-9'd30,10'd370};
ram[21194] = {-9'd27,10'd373};
ram[21195] = {-9'd24,10'd376};
ram[21196] = {-9'd21,10'd380};
ram[21197] = {-9'd18,10'd383};
ram[21198] = {-9'd15,10'd386};
ram[21199] = {-9'd11,10'd389};
ram[21200] = {-9'd8,10'd392};
ram[21201] = {-9'd5,10'd395};
ram[21202] = {-9'd2,10'd398};
ram[21203] = {9'd1,-10'd399};
ram[21204] = {9'd4,-10'd396};
ram[21205] = {9'd7,-10'd393};
ram[21206] = {9'd10,-10'd390};
ram[21207] = {9'd14,-10'd387};
ram[21208] = {9'd17,-10'd384};
ram[21209] = {9'd20,-10'd381};
ram[21210] = {9'd23,-10'd377};
ram[21211] = {9'd26,-10'd374};
ram[21212] = {9'd29,-10'd371};
ram[21213] = {9'd32,-10'd368};
ram[21214] = {9'd36,-10'd365};
ram[21215] = {9'd39,-10'd362};
ram[21216] = {9'd42,-10'd359};
ram[21217] = {9'd45,-10'd355};
ram[21218] = {9'd48,-10'd352};
ram[21219] = {9'd51,-10'd349};
ram[21220] = {9'd54,-10'd346};
ram[21221] = {9'd58,-10'd343};
ram[21222] = {9'd61,-10'd340};
ram[21223] = {9'd64,-10'd337};
ram[21224] = {9'd67,-10'd334};
ram[21225] = {9'd70,-10'd330};
ram[21226] = {9'd73,-10'd327};
ram[21227] = {9'd76,-10'd324};
ram[21228] = {9'd80,-10'd321};
ram[21229] = {9'd83,-10'd318};
ram[21230] = {9'd86,-10'd315};
ram[21231] = {9'd89,-10'd312};
ram[21232] = {9'd92,-10'd308};
ram[21233] = {9'd95,-10'd305};
ram[21234] = {9'd98,-10'd302};
ram[21235] = {-9'd99,-10'd299};
ram[21236] = {-9'd96,-10'd296};
ram[21237] = {-9'd92,-10'd293};
ram[21238] = {-9'd89,-10'd290};
ram[21239] = {-9'd86,-10'd286};
ram[21240] = {-9'd83,-10'd283};
ram[21241] = {-9'd80,-10'd280};
ram[21242] = {-9'd77,-10'd277};
ram[21243] = {-9'd74,-10'd274};
ram[21244] = {-9'd70,-10'd271};
ram[21245] = {-9'd67,-10'd268};
ram[21246] = {-9'd64,-10'd264};
ram[21247] = {-9'd61,-10'd261};
ram[21248] = {-9'd61,-10'd261};
ram[21249] = {-9'd58,-10'd258};
ram[21250] = {-9'd55,-10'd255};
ram[21251] = {-9'd52,-10'd252};
ram[21252] = {-9'd48,-10'd249};
ram[21253] = {-9'd45,-10'd246};
ram[21254] = {-9'd42,-10'd242};
ram[21255] = {-9'd39,-10'd239};
ram[21256] = {-9'd36,-10'd236};
ram[21257] = {-9'd33,-10'd233};
ram[21258] = {-9'd30,-10'd230};
ram[21259] = {-9'd26,-10'd227};
ram[21260] = {-9'd23,-10'd224};
ram[21261] = {-9'd20,-10'd220};
ram[21262] = {-9'd17,-10'd217};
ram[21263] = {-9'd14,-10'd214};
ram[21264] = {-9'd11,-10'd211};
ram[21265] = {-9'd8,-10'd208};
ram[21266] = {-9'd4,-10'd205};
ram[21267] = {-9'd1,-10'd202};
ram[21268] = {9'd2,-10'd198};
ram[21269] = {9'd5,-10'd195};
ram[21270] = {9'd8,-10'd192};
ram[21271] = {9'd11,-10'd189};
ram[21272] = {9'd14,-10'd186};
ram[21273] = {9'd18,-10'd183};
ram[21274] = {9'd21,-10'd180};
ram[21275] = {9'd24,-10'd176};
ram[21276] = {9'd27,-10'd173};
ram[21277] = {9'd30,-10'd170};
ram[21278] = {9'd33,-10'd167};
ram[21279] = {9'd36,-10'd164};
ram[21280] = {9'd40,-10'd161};
ram[21281] = {9'd43,-10'd158};
ram[21282] = {9'd46,-10'd154};
ram[21283] = {9'd49,-10'd151};
ram[21284] = {9'd52,-10'd148};
ram[21285] = {9'd55,-10'd145};
ram[21286] = {9'd58,-10'd142};
ram[21287] = {9'd62,-10'd139};
ram[21288] = {9'd65,-10'd136};
ram[21289] = {9'd68,-10'd132};
ram[21290] = {9'd71,-10'd129};
ram[21291] = {9'd74,-10'd126};
ram[21292] = {9'd77,-10'd123};
ram[21293] = {9'd80,-10'd120};
ram[21294] = {9'd84,-10'd117};
ram[21295] = {9'd87,-10'd114};
ram[21296] = {9'd90,-10'd110};
ram[21297] = {9'd93,-10'd107};
ram[21298] = {9'd96,-10'd104};
ram[21299] = {9'd99,-10'd101};
ram[21300] = {-9'd98,-10'd98};
ram[21301] = {-9'd95,-10'd95};
ram[21302] = {-9'd92,-10'd92};
ram[21303] = {-9'd88,-10'd88};
ram[21304] = {-9'd85,-10'd85};
ram[21305] = {-9'd82,-10'd82};
ram[21306] = {-9'd79,-10'd79};
ram[21307] = {-9'd76,-10'd76};
ram[21308] = {-9'd73,-10'd73};
ram[21309] = {-9'd70,-10'd70};
ram[21310] = {-9'd66,-10'd66};
ram[21311] = {-9'd63,-10'd63};
ram[21312] = {-9'd60,-10'd60};
ram[21313] = {-9'd57,-10'd57};
ram[21314] = {-9'd54,-10'd54};
ram[21315] = {-9'd51,-10'd51};
ram[21316] = {-9'd48,-10'd48};
ram[21317] = {-9'd44,-10'd44};
ram[21318] = {-9'd41,-10'd41};
ram[21319] = {-9'd38,-10'd38};
ram[21320] = {-9'd35,-10'd35};
ram[21321] = {-9'd32,-10'd32};
ram[21322] = {-9'd29,-10'd29};
ram[21323] = {-9'd26,-10'd26};
ram[21324] = {-9'd22,-10'd22};
ram[21325] = {-9'd19,-10'd19};
ram[21326] = {-9'd16,-10'd16};
ram[21327] = {-9'd13,-10'd13};
ram[21328] = {-9'd10,-10'd10};
ram[21329] = {-9'd7,-10'd7};
ram[21330] = {-9'd4,-10'd4};
ram[21331] = {9'd0,10'd0};
ram[21332] = {9'd3,10'd3};
ram[21333] = {9'd6,10'd6};
ram[21334] = {9'd9,10'd9};
ram[21335] = {9'd12,10'd12};
ram[21336] = {9'd15,10'd15};
ram[21337] = {9'd18,10'd18};
ram[21338] = {9'd21,10'd21};
ram[21339] = {9'd25,10'd25};
ram[21340] = {9'd28,10'd28};
ram[21341] = {9'd31,10'd31};
ram[21342] = {9'd34,10'd34};
ram[21343] = {9'd37,10'd37};
ram[21344] = {9'd40,10'd40};
ram[21345] = {9'd43,10'd43};
ram[21346] = {9'd47,10'd47};
ram[21347] = {9'd50,10'd50};
ram[21348] = {9'd53,10'd53};
ram[21349] = {9'd56,10'd56};
ram[21350] = {9'd59,10'd59};
ram[21351] = {9'd62,10'd62};
ram[21352] = {9'd65,10'd65};
ram[21353] = {9'd69,10'd69};
ram[21354] = {9'd72,10'd72};
ram[21355] = {9'd75,10'd75};
ram[21356] = {9'd78,10'd78};
ram[21357] = {9'd81,10'd81};
ram[21358] = {9'd84,10'd84};
ram[21359] = {9'd87,10'd87};
ram[21360] = {9'd91,10'd91};
ram[21361] = {9'd94,10'd94};
ram[21362] = {9'd97,10'd97};
ram[21363] = {-9'd100,10'd100};
ram[21364] = {-9'd97,10'd103};
ram[21365] = {-9'd94,10'd106};
ram[21366] = {-9'd91,10'd109};
ram[21367] = {-9'd88,10'd113};
ram[21368] = {-9'd85,10'd116};
ram[21369] = {-9'd81,10'd119};
ram[21370] = {-9'd78,10'd122};
ram[21371] = {-9'd75,10'd125};
ram[21372] = {-9'd72,10'd128};
ram[21373] = {-9'd69,10'd131};
ram[21374] = {-9'd66,10'd135};
ram[21375] = {-9'd63,10'd138};
ram[21376] = {-9'd63,10'd138};
ram[21377] = {-9'd59,10'd141};
ram[21378] = {-9'd56,10'd144};
ram[21379] = {-9'd53,10'd147};
ram[21380] = {-9'd50,10'd150};
ram[21381] = {-9'd47,10'd153};
ram[21382] = {-9'd44,10'd157};
ram[21383] = {-9'd41,10'd160};
ram[21384] = {-9'd37,10'd163};
ram[21385] = {-9'd34,10'd166};
ram[21386] = {-9'd31,10'd169};
ram[21387] = {-9'd28,10'd172};
ram[21388] = {-9'd25,10'd175};
ram[21389] = {-9'd22,10'd179};
ram[21390] = {-9'd19,10'd182};
ram[21391] = {-9'd15,10'd185};
ram[21392] = {-9'd12,10'd188};
ram[21393] = {-9'd9,10'd191};
ram[21394] = {-9'd6,10'd194};
ram[21395] = {-9'd3,10'd197};
ram[21396] = {9'd0,10'd201};
ram[21397] = {9'd3,10'd204};
ram[21398] = {9'd7,10'd207};
ram[21399] = {9'd10,10'd210};
ram[21400] = {9'd13,10'd213};
ram[21401] = {9'd16,10'd216};
ram[21402] = {9'd19,10'd219};
ram[21403] = {9'd22,10'd223};
ram[21404] = {9'd25,10'd226};
ram[21405] = {9'd29,10'd229};
ram[21406] = {9'd32,10'd232};
ram[21407] = {9'd35,10'd235};
ram[21408] = {9'd38,10'd238};
ram[21409] = {9'd41,10'd241};
ram[21410] = {9'd44,10'd245};
ram[21411] = {9'd47,10'd248};
ram[21412] = {9'd51,10'd251};
ram[21413] = {9'd54,10'd254};
ram[21414] = {9'd57,10'd257};
ram[21415] = {9'd60,10'd260};
ram[21416] = {9'd63,10'd263};
ram[21417] = {9'd66,10'd267};
ram[21418] = {9'd69,10'd270};
ram[21419] = {9'd73,10'd273};
ram[21420] = {9'd76,10'd276};
ram[21421] = {9'd79,10'd279};
ram[21422] = {9'd82,10'd282};
ram[21423] = {9'd85,10'd285};
ram[21424] = {9'd88,10'd289};
ram[21425] = {9'd91,10'd292};
ram[21426] = {9'd95,10'd295};
ram[21427] = {9'd98,10'd298};
ram[21428] = {-9'd99,10'd301};
ram[21429] = {-9'd96,10'd304};
ram[21430] = {-9'd93,10'd307};
ram[21431] = {-9'd90,10'd311};
ram[21432] = {-9'd87,10'd314};
ram[21433] = {-9'd84,10'd317};
ram[21434] = {-9'd81,10'd320};
ram[21435] = {-9'd77,10'd323};
ram[21436] = {-9'd74,10'd326};
ram[21437] = {-9'd71,10'd329};
ram[21438] = {-9'd68,10'd333};
ram[21439] = {-9'd65,10'd336};
ram[21440] = {-9'd62,10'd339};
ram[21441] = {-9'd59,10'd342};
ram[21442] = {-9'd55,10'd345};
ram[21443] = {-9'd52,10'd348};
ram[21444] = {-9'd49,10'd351};
ram[21445] = {-9'd46,10'd354};
ram[21446] = {-9'd43,10'd358};
ram[21447] = {-9'd40,10'd361};
ram[21448] = {-9'd37,10'd364};
ram[21449] = {-9'd33,10'd367};
ram[21450] = {-9'd30,10'd370};
ram[21451] = {-9'd27,10'd373};
ram[21452] = {-9'd24,10'd376};
ram[21453] = {-9'd21,10'd380};
ram[21454] = {-9'd18,10'd383};
ram[21455] = {-9'd15,10'd386};
ram[21456] = {-9'd11,10'd389};
ram[21457] = {-9'd8,10'd392};
ram[21458] = {-9'd5,10'd395};
ram[21459] = {-9'd2,10'd398};
ram[21460] = {9'd1,-10'd399};
ram[21461] = {9'd4,-10'd396};
ram[21462] = {9'd7,-10'd393};
ram[21463] = {9'd10,-10'd390};
ram[21464] = {9'd14,-10'd387};
ram[21465] = {9'd17,-10'd384};
ram[21466] = {9'd20,-10'd381};
ram[21467] = {9'd23,-10'd377};
ram[21468] = {9'd26,-10'd374};
ram[21469] = {9'd29,-10'd371};
ram[21470] = {9'd32,-10'd368};
ram[21471] = {9'd36,-10'd365};
ram[21472] = {9'd39,-10'd362};
ram[21473] = {9'd42,-10'd359};
ram[21474] = {9'd45,-10'd355};
ram[21475] = {9'd48,-10'd352};
ram[21476] = {9'd51,-10'd349};
ram[21477] = {9'd54,-10'd346};
ram[21478] = {9'd58,-10'd343};
ram[21479] = {9'd61,-10'd340};
ram[21480] = {9'd64,-10'd337};
ram[21481] = {9'd67,-10'd334};
ram[21482] = {9'd70,-10'd330};
ram[21483] = {9'd73,-10'd327};
ram[21484] = {9'd76,-10'd324};
ram[21485] = {9'd80,-10'd321};
ram[21486] = {9'd83,-10'd318};
ram[21487] = {9'd86,-10'd315};
ram[21488] = {9'd89,-10'd312};
ram[21489] = {9'd92,-10'd308};
ram[21490] = {9'd95,-10'd305};
ram[21491] = {9'd98,-10'd302};
ram[21492] = {-9'd99,-10'd299};
ram[21493] = {-9'd96,-10'd296};
ram[21494] = {-9'd92,-10'd293};
ram[21495] = {-9'd89,-10'd290};
ram[21496] = {-9'd86,-10'd286};
ram[21497] = {-9'd83,-10'd283};
ram[21498] = {-9'd80,-10'd280};
ram[21499] = {-9'd77,-10'd277};
ram[21500] = {-9'd74,-10'd274};
ram[21501] = {-9'd70,-10'd271};
ram[21502] = {-9'd67,-10'd268};
ram[21503] = {-9'd64,-10'd264};
ram[21504] = {-9'd64,-10'd264};
ram[21505] = {-9'd61,-10'd261};
ram[21506] = {-9'd58,-10'd258};
ram[21507] = {-9'd55,-10'd255};
ram[21508] = {-9'd52,-10'd252};
ram[21509] = {-9'd48,-10'd249};
ram[21510] = {-9'd45,-10'd246};
ram[21511] = {-9'd42,-10'd242};
ram[21512] = {-9'd39,-10'd239};
ram[21513] = {-9'd36,-10'd236};
ram[21514] = {-9'd33,-10'd233};
ram[21515] = {-9'd30,-10'd230};
ram[21516] = {-9'd26,-10'd227};
ram[21517] = {-9'd23,-10'd224};
ram[21518] = {-9'd20,-10'd220};
ram[21519] = {-9'd17,-10'd217};
ram[21520] = {-9'd14,-10'd214};
ram[21521] = {-9'd11,-10'd211};
ram[21522] = {-9'd8,-10'd208};
ram[21523] = {-9'd4,-10'd205};
ram[21524] = {-9'd1,-10'd202};
ram[21525] = {9'd2,-10'd198};
ram[21526] = {9'd5,-10'd195};
ram[21527] = {9'd8,-10'd192};
ram[21528] = {9'd11,-10'd189};
ram[21529] = {9'd14,-10'd186};
ram[21530] = {9'd18,-10'd183};
ram[21531] = {9'd21,-10'd180};
ram[21532] = {9'd24,-10'd176};
ram[21533] = {9'd27,-10'd173};
ram[21534] = {9'd30,-10'd170};
ram[21535] = {9'd33,-10'd167};
ram[21536] = {9'd36,-10'd164};
ram[21537] = {9'd40,-10'd161};
ram[21538] = {9'd43,-10'd158};
ram[21539] = {9'd46,-10'd154};
ram[21540] = {9'd49,-10'd151};
ram[21541] = {9'd52,-10'd148};
ram[21542] = {9'd55,-10'd145};
ram[21543] = {9'd58,-10'd142};
ram[21544] = {9'd62,-10'd139};
ram[21545] = {9'd65,-10'd136};
ram[21546] = {9'd68,-10'd132};
ram[21547] = {9'd71,-10'd129};
ram[21548] = {9'd74,-10'd126};
ram[21549] = {9'd77,-10'd123};
ram[21550] = {9'd80,-10'd120};
ram[21551] = {9'd84,-10'd117};
ram[21552] = {9'd87,-10'd114};
ram[21553] = {9'd90,-10'd110};
ram[21554] = {9'd93,-10'd107};
ram[21555] = {9'd96,-10'd104};
ram[21556] = {9'd99,-10'd101};
ram[21557] = {-9'd98,-10'd98};
ram[21558] = {-9'd95,-10'd95};
ram[21559] = {-9'd92,-10'd92};
ram[21560] = {-9'd88,-10'd88};
ram[21561] = {-9'd85,-10'd85};
ram[21562] = {-9'd82,-10'd82};
ram[21563] = {-9'd79,-10'd79};
ram[21564] = {-9'd76,-10'd76};
ram[21565] = {-9'd73,-10'd73};
ram[21566] = {-9'd70,-10'd70};
ram[21567] = {-9'd66,-10'd66};
ram[21568] = {-9'd63,-10'd63};
ram[21569] = {-9'd60,-10'd60};
ram[21570] = {-9'd57,-10'd57};
ram[21571] = {-9'd54,-10'd54};
ram[21572] = {-9'd51,-10'd51};
ram[21573] = {-9'd48,-10'd48};
ram[21574] = {-9'd44,-10'd44};
ram[21575] = {-9'd41,-10'd41};
ram[21576] = {-9'd38,-10'd38};
ram[21577] = {-9'd35,-10'd35};
ram[21578] = {-9'd32,-10'd32};
ram[21579] = {-9'd29,-10'd29};
ram[21580] = {-9'd26,-10'd26};
ram[21581] = {-9'd22,-10'd22};
ram[21582] = {-9'd19,-10'd19};
ram[21583] = {-9'd16,-10'd16};
ram[21584] = {-9'd13,-10'd13};
ram[21585] = {-9'd10,-10'd10};
ram[21586] = {-9'd7,-10'd7};
ram[21587] = {-9'd4,-10'd4};
ram[21588] = {9'd0,10'd0};
ram[21589] = {9'd3,10'd3};
ram[21590] = {9'd6,10'd6};
ram[21591] = {9'd9,10'd9};
ram[21592] = {9'd12,10'd12};
ram[21593] = {9'd15,10'd15};
ram[21594] = {9'd18,10'd18};
ram[21595] = {9'd21,10'd21};
ram[21596] = {9'd25,10'd25};
ram[21597] = {9'd28,10'd28};
ram[21598] = {9'd31,10'd31};
ram[21599] = {9'd34,10'd34};
ram[21600] = {9'd37,10'd37};
ram[21601] = {9'd40,10'd40};
ram[21602] = {9'd43,10'd43};
ram[21603] = {9'd47,10'd47};
ram[21604] = {9'd50,10'd50};
ram[21605] = {9'd53,10'd53};
ram[21606] = {9'd56,10'd56};
ram[21607] = {9'd59,10'd59};
ram[21608] = {9'd62,10'd62};
ram[21609] = {9'd65,10'd65};
ram[21610] = {9'd69,10'd69};
ram[21611] = {9'd72,10'd72};
ram[21612] = {9'd75,10'd75};
ram[21613] = {9'd78,10'd78};
ram[21614] = {9'd81,10'd81};
ram[21615] = {9'd84,10'd84};
ram[21616] = {9'd87,10'd87};
ram[21617] = {9'd91,10'd91};
ram[21618] = {9'd94,10'd94};
ram[21619] = {9'd97,10'd97};
ram[21620] = {-9'd100,10'd100};
ram[21621] = {-9'd97,10'd103};
ram[21622] = {-9'd94,10'd106};
ram[21623] = {-9'd91,10'd109};
ram[21624] = {-9'd88,10'd113};
ram[21625] = {-9'd85,10'd116};
ram[21626] = {-9'd81,10'd119};
ram[21627] = {-9'd78,10'd122};
ram[21628] = {-9'd75,10'd125};
ram[21629] = {-9'd72,10'd128};
ram[21630] = {-9'd69,10'd131};
ram[21631] = {-9'd66,10'd135};
ram[21632] = {-9'd66,10'd135};
ram[21633] = {-9'd63,10'd138};
ram[21634] = {-9'd59,10'd141};
ram[21635] = {-9'd56,10'd144};
ram[21636] = {-9'd53,10'd147};
ram[21637] = {-9'd50,10'd150};
ram[21638] = {-9'd47,10'd153};
ram[21639] = {-9'd44,10'd157};
ram[21640] = {-9'd41,10'd160};
ram[21641] = {-9'd37,10'd163};
ram[21642] = {-9'd34,10'd166};
ram[21643] = {-9'd31,10'd169};
ram[21644] = {-9'd28,10'd172};
ram[21645] = {-9'd25,10'd175};
ram[21646] = {-9'd22,10'd179};
ram[21647] = {-9'd19,10'd182};
ram[21648] = {-9'd15,10'd185};
ram[21649] = {-9'd12,10'd188};
ram[21650] = {-9'd9,10'd191};
ram[21651] = {-9'd6,10'd194};
ram[21652] = {-9'd3,10'd197};
ram[21653] = {9'd0,10'd201};
ram[21654] = {9'd3,10'd204};
ram[21655] = {9'd7,10'd207};
ram[21656] = {9'd10,10'd210};
ram[21657] = {9'd13,10'd213};
ram[21658] = {9'd16,10'd216};
ram[21659] = {9'd19,10'd219};
ram[21660] = {9'd22,10'd223};
ram[21661] = {9'd25,10'd226};
ram[21662] = {9'd29,10'd229};
ram[21663] = {9'd32,10'd232};
ram[21664] = {9'd35,10'd235};
ram[21665] = {9'd38,10'd238};
ram[21666] = {9'd41,10'd241};
ram[21667] = {9'd44,10'd245};
ram[21668] = {9'd47,10'd248};
ram[21669] = {9'd51,10'd251};
ram[21670] = {9'd54,10'd254};
ram[21671] = {9'd57,10'd257};
ram[21672] = {9'd60,10'd260};
ram[21673] = {9'd63,10'd263};
ram[21674] = {9'd66,10'd267};
ram[21675] = {9'd69,10'd270};
ram[21676] = {9'd73,10'd273};
ram[21677] = {9'd76,10'd276};
ram[21678] = {9'd79,10'd279};
ram[21679] = {9'd82,10'd282};
ram[21680] = {9'd85,10'd285};
ram[21681] = {9'd88,10'd289};
ram[21682] = {9'd91,10'd292};
ram[21683] = {9'd95,10'd295};
ram[21684] = {9'd98,10'd298};
ram[21685] = {-9'd99,10'd301};
ram[21686] = {-9'd96,10'd304};
ram[21687] = {-9'd93,10'd307};
ram[21688] = {-9'd90,10'd311};
ram[21689] = {-9'd87,10'd314};
ram[21690] = {-9'd84,10'd317};
ram[21691] = {-9'd81,10'd320};
ram[21692] = {-9'd77,10'd323};
ram[21693] = {-9'd74,10'd326};
ram[21694] = {-9'd71,10'd329};
ram[21695] = {-9'd68,10'd333};
ram[21696] = {-9'd65,10'd336};
ram[21697] = {-9'd62,10'd339};
ram[21698] = {-9'd59,10'd342};
ram[21699] = {-9'd55,10'd345};
ram[21700] = {-9'd52,10'd348};
ram[21701] = {-9'd49,10'd351};
ram[21702] = {-9'd46,10'd354};
ram[21703] = {-9'd43,10'd358};
ram[21704] = {-9'd40,10'd361};
ram[21705] = {-9'd37,10'd364};
ram[21706] = {-9'd33,10'd367};
ram[21707] = {-9'd30,10'd370};
ram[21708] = {-9'd27,10'd373};
ram[21709] = {-9'd24,10'd376};
ram[21710] = {-9'd21,10'd380};
ram[21711] = {-9'd18,10'd383};
ram[21712] = {-9'd15,10'd386};
ram[21713] = {-9'd11,10'd389};
ram[21714] = {-9'd8,10'd392};
ram[21715] = {-9'd5,10'd395};
ram[21716] = {-9'd2,10'd398};
ram[21717] = {9'd1,-10'd399};
ram[21718] = {9'd4,-10'd396};
ram[21719] = {9'd7,-10'd393};
ram[21720] = {9'd10,-10'd390};
ram[21721] = {9'd14,-10'd387};
ram[21722] = {9'd17,-10'd384};
ram[21723] = {9'd20,-10'd381};
ram[21724] = {9'd23,-10'd377};
ram[21725] = {9'd26,-10'd374};
ram[21726] = {9'd29,-10'd371};
ram[21727] = {9'd32,-10'd368};
ram[21728] = {9'd36,-10'd365};
ram[21729] = {9'd39,-10'd362};
ram[21730] = {9'd42,-10'd359};
ram[21731] = {9'd45,-10'd355};
ram[21732] = {9'd48,-10'd352};
ram[21733] = {9'd51,-10'd349};
ram[21734] = {9'd54,-10'd346};
ram[21735] = {9'd58,-10'd343};
ram[21736] = {9'd61,-10'd340};
ram[21737] = {9'd64,-10'd337};
ram[21738] = {9'd67,-10'd334};
ram[21739] = {9'd70,-10'd330};
ram[21740] = {9'd73,-10'd327};
ram[21741] = {9'd76,-10'd324};
ram[21742] = {9'd80,-10'd321};
ram[21743] = {9'd83,-10'd318};
ram[21744] = {9'd86,-10'd315};
ram[21745] = {9'd89,-10'd312};
ram[21746] = {9'd92,-10'd308};
ram[21747] = {9'd95,-10'd305};
ram[21748] = {9'd98,-10'd302};
ram[21749] = {-9'd99,-10'd299};
ram[21750] = {-9'd96,-10'd296};
ram[21751] = {-9'd92,-10'd293};
ram[21752] = {-9'd89,-10'd290};
ram[21753] = {-9'd86,-10'd286};
ram[21754] = {-9'd83,-10'd283};
ram[21755] = {-9'd80,-10'd280};
ram[21756] = {-9'd77,-10'd277};
ram[21757] = {-9'd74,-10'd274};
ram[21758] = {-9'd70,-10'd271};
ram[21759] = {-9'd67,-10'd268};
ram[21760] = {-9'd67,-10'd268};
ram[21761] = {-9'd64,-10'd264};
ram[21762] = {-9'd61,-10'd261};
ram[21763] = {-9'd58,-10'd258};
ram[21764] = {-9'd55,-10'd255};
ram[21765] = {-9'd52,-10'd252};
ram[21766] = {-9'd48,-10'd249};
ram[21767] = {-9'd45,-10'd246};
ram[21768] = {-9'd42,-10'd242};
ram[21769] = {-9'd39,-10'd239};
ram[21770] = {-9'd36,-10'd236};
ram[21771] = {-9'd33,-10'd233};
ram[21772] = {-9'd30,-10'd230};
ram[21773] = {-9'd26,-10'd227};
ram[21774] = {-9'd23,-10'd224};
ram[21775] = {-9'd20,-10'd220};
ram[21776] = {-9'd17,-10'd217};
ram[21777] = {-9'd14,-10'd214};
ram[21778] = {-9'd11,-10'd211};
ram[21779] = {-9'd8,-10'd208};
ram[21780] = {-9'd4,-10'd205};
ram[21781] = {-9'd1,-10'd202};
ram[21782] = {9'd2,-10'd198};
ram[21783] = {9'd5,-10'd195};
ram[21784] = {9'd8,-10'd192};
ram[21785] = {9'd11,-10'd189};
ram[21786] = {9'd14,-10'd186};
ram[21787] = {9'd18,-10'd183};
ram[21788] = {9'd21,-10'd180};
ram[21789] = {9'd24,-10'd176};
ram[21790] = {9'd27,-10'd173};
ram[21791] = {9'd30,-10'd170};
ram[21792] = {9'd33,-10'd167};
ram[21793] = {9'd36,-10'd164};
ram[21794] = {9'd40,-10'd161};
ram[21795] = {9'd43,-10'd158};
ram[21796] = {9'd46,-10'd154};
ram[21797] = {9'd49,-10'd151};
ram[21798] = {9'd52,-10'd148};
ram[21799] = {9'd55,-10'd145};
ram[21800] = {9'd58,-10'd142};
ram[21801] = {9'd62,-10'd139};
ram[21802] = {9'd65,-10'd136};
ram[21803] = {9'd68,-10'd132};
ram[21804] = {9'd71,-10'd129};
ram[21805] = {9'd74,-10'd126};
ram[21806] = {9'd77,-10'd123};
ram[21807] = {9'd80,-10'd120};
ram[21808] = {9'd84,-10'd117};
ram[21809] = {9'd87,-10'd114};
ram[21810] = {9'd90,-10'd110};
ram[21811] = {9'd93,-10'd107};
ram[21812] = {9'd96,-10'd104};
ram[21813] = {9'd99,-10'd101};
ram[21814] = {-9'd98,-10'd98};
ram[21815] = {-9'd95,-10'd95};
ram[21816] = {-9'd92,-10'd92};
ram[21817] = {-9'd88,-10'd88};
ram[21818] = {-9'd85,-10'd85};
ram[21819] = {-9'd82,-10'd82};
ram[21820] = {-9'd79,-10'd79};
ram[21821] = {-9'd76,-10'd76};
ram[21822] = {-9'd73,-10'd73};
ram[21823] = {-9'd70,-10'd70};
ram[21824] = {-9'd66,-10'd66};
ram[21825] = {-9'd63,-10'd63};
ram[21826] = {-9'd60,-10'd60};
ram[21827] = {-9'd57,-10'd57};
ram[21828] = {-9'd54,-10'd54};
ram[21829] = {-9'd51,-10'd51};
ram[21830] = {-9'd48,-10'd48};
ram[21831] = {-9'd44,-10'd44};
ram[21832] = {-9'd41,-10'd41};
ram[21833] = {-9'd38,-10'd38};
ram[21834] = {-9'd35,-10'd35};
ram[21835] = {-9'd32,-10'd32};
ram[21836] = {-9'd29,-10'd29};
ram[21837] = {-9'd26,-10'd26};
ram[21838] = {-9'd22,-10'd22};
ram[21839] = {-9'd19,-10'd19};
ram[21840] = {-9'd16,-10'd16};
ram[21841] = {-9'd13,-10'd13};
ram[21842] = {-9'd10,-10'd10};
ram[21843] = {-9'd7,-10'd7};
ram[21844] = {-9'd4,-10'd4};
ram[21845] = {9'd0,10'd0};
ram[21846] = {9'd3,10'd3};
ram[21847] = {9'd6,10'd6};
ram[21848] = {9'd9,10'd9};
ram[21849] = {9'd12,10'd12};
ram[21850] = {9'd15,10'd15};
ram[21851] = {9'd18,10'd18};
ram[21852] = {9'd21,10'd21};
ram[21853] = {9'd25,10'd25};
ram[21854] = {9'd28,10'd28};
ram[21855] = {9'd31,10'd31};
ram[21856] = {9'd34,10'd34};
ram[21857] = {9'd37,10'd37};
ram[21858] = {9'd40,10'd40};
ram[21859] = {9'd43,10'd43};
ram[21860] = {9'd47,10'd47};
ram[21861] = {9'd50,10'd50};
ram[21862] = {9'd53,10'd53};
ram[21863] = {9'd56,10'd56};
ram[21864] = {9'd59,10'd59};
ram[21865] = {9'd62,10'd62};
ram[21866] = {9'd65,10'd65};
ram[21867] = {9'd69,10'd69};
ram[21868] = {9'd72,10'd72};
ram[21869] = {9'd75,10'd75};
ram[21870] = {9'd78,10'd78};
ram[21871] = {9'd81,10'd81};
ram[21872] = {9'd84,10'd84};
ram[21873] = {9'd87,10'd87};
ram[21874] = {9'd91,10'd91};
ram[21875] = {9'd94,10'd94};
ram[21876] = {9'd97,10'd97};
ram[21877] = {-9'd100,10'd100};
ram[21878] = {-9'd97,10'd103};
ram[21879] = {-9'd94,10'd106};
ram[21880] = {-9'd91,10'd109};
ram[21881] = {-9'd88,10'd113};
ram[21882] = {-9'd85,10'd116};
ram[21883] = {-9'd81,10'd119};
ram[21884] = {-9'd78,10'd122};
ram[21885] = {-9'd75,10'd125};
ram[21886] = {-9'd72,10'd128};
ram[21887] = {-9'd69,10'd131};
ram[21888] = {-9'd69,10'd131};
ram[21889] = {-9'd66,10'd135};
ram[21890] = {-9'd63,10'd138};
ram[21891] = {-9'd59,10'd141};
ram[21892] = {-9'd56,10'd144};
ram[21893] = {-9'd53,10'd147};
ram[21894] = {-9'd50,10'd150};
ram[21895] = {-9'd47,10'd153};
ram[21896] = {-9'd44,10'd157};
ram[21897] = {-9'd41,10'd160};
ram[21898] = {-9'd37,10'd163};
ram[21899] = {-9'd34,10'd166};
ram[21900] = {-9'd31,10'd169};
ram[21901] = {-9'd28,10'd172};
ram[21902] = {-9'd25,10'd175};
ram[21903] = {-9'd22,10'd179};
ram[21904] = {-9'd19,10'd182};
ram[21905] = {-9'd15,10'd185};
ram[21906] = {-9'd12,10'd188};
ram[21907] = {-9'd9,10'd191};
ram[21908] = {-9'd6,10'd194};
ram[21909] = {-9'd3,10'd197};
ram[21910] = {9'd0,10'd201};
ram[21911] = {9'd3,10'd204};
ram[21912] = {9'd7,10'd207};
ram[21913] = {9'd10,10'd210};
ram[21914] = {9'd13,10'd213};
ram[21915] = {9'd16,10'd216};
ram[21916] = {9'd19,10'd219};
ram[21917] = {9'd22,10'd223};
ram[21918] = {9'd25,10'd226};
ram[21919] = {9'd29,10'd229};
ram[21920] = {9'd32,10'd232};
ram[21921] = {9'd35,10'd235};
ram[21922] = {9'd38,10'd238};
ram[21923] = {9'd41,10'd241};
ram[21924] = {9'd44,10'd245};
ram[21925] = {9'd47,10'd248};
ram[21926] = {9'd51,10'd251};
ram[21927] = {9'd54,10'd254};
ram[21928] = {9'd57,10'd257};
ram[21929] = {9'd60,10'd260};
ram[21930] = {9'd63,10'd263};
ram[21931] = {9'd66,10'd267};
ram[21932] = {9'd69,10'd270};
ram[21933] = {9'd73,10'd273};
ram[21934] = {9'd76,10'd276};
ram[21935] = {9'd79,10'd279};
ram[21936] = {9'd82,10'd282};
ram[21937] = {9'd85,10'd285};
ram[21938] = {9'd88,10'd289};
ram[21939] = {9'd91,10'd292};
ram[21940] = {9'd95,10'd295};
ram[21941] = {9'd98,10'd298};
ram[21942] = {-9'd99,10'd301};
ram[21943] = {-9'd96,10'd304};
ram[21944] = {-9'd93,10'd307};
ram[21945] = {-9'd90,10'd311};
ram[21946] = {-9'd87,10'd314};
ram[21947] = {-9'd84,10'd317};
ram[21948] = {-9'd81,10'd320};
ram[21949] = {-9'd77,10'd323};
ram[21950] = {-9'd74,10'd326};
ram[21951] = {-9'd71,10'd329};
ram[21952] = {-9'd68,10'd333};
ram[21953] = {-9'd65,10'd336};
ram[21954] = {-9'd62,10'd339};
ram[21955] = {-9'd59,10'd342};
ram[21956] = {-9'd55,10'd345};
ram[21957] = {-9'd52,10'd348};
ram[21958] = {-9'd49,10'd351};
ram[21959] = {-9'd46,10'd354};
ram[21960] = {-9'd43,10'd358};
ram[21961] = {-9'd40,10'd361};
ram[21962] = {-9'd37,10'd364};
ram[21963] = {-9'd33,10'd367};
ram[21964] = {-9'd30,10'd370};
ram[21965] = {-9'd27,10'd373};
ram[21966] = {-9'd24,10'd376};
ram[21967] = {-9'd21,10'd380};
ram[21968] = {-9'd18,10'd383};
ram[21969] = {-9'd15,10'd386};
ram[21970] = {-9'd11,10'd389};
ram[21971] = {-9'd8,10'd392};
ram[21972] = {-9'd5,10'd395};
ram[21973] = {-9'd2,10'd398};
ram[21974] = {9'd1,-10'd399};
ram[21975] = {9'd4,-10'd396};
ram[21976] = {9'd7,-10'd393};
ram[21977] = {9'd10,-10'd390};
ram[21978] = {9'd14,-10'd387};
ram[21979] = {9'd17,-10'd384};
ram[21980] = {9'd20,-10'd381};
ram[21981] = {9'd23,-10'd377};
ram[21982] = {9'd26,-10'd374};
ram[21983] = {9'd29,-10'd371};
ram[21984] = {9'd32,-10'd368};
ram[21985] = {9'd36,-10'd365};
ram[21986] = {9'd39,-10'd362};
ram[21987] = {9'd42,-10'd359};
ram[21988] = {9'd45,-10'd355};
ram[21989] = {9'd48,-10'd352};
ram[21990] = {9'd51,-10'd349};
ram[21991] = {9'd54,-10'd346};
ram[21992] = {9'd58,-10'd343};
ram[21993] = {9'd61,-10'd340};
ram[21994] = {9'd64,-10'd337};
ram[21995] = {9'd67,-10'd334};
ram[21996] = {9'd70,-10'd330};
ram[21997] = {9'd73,-10'd327};
ram[21998] = {9'd76,-10'd324};
ram[21999] = {9'd80,-10'd321};
ram[22000] = {9'd83,-10'd318};
ram[22001] = {9'd86,-10'd315};
ram[22002] = {9'd89,-10'd312};
ram[22003] = {9'd92,-10'd308};
ram[22004] = {9'd95,-10'd305};
ram[22005] = {9'd98,-10'd302};
ram[22006] = {-9'd99,-10'd299};
ram[22007] = {-9'd96,-10'd296};
ram[22008] = {-9'd92,-10'd293};
ram[22009] = {-9'd89,-10'd290};
ram[22010] = {-9'd86,-10'd286};
ram[22011] = {-9'd83,-10'd283};
ram[22012] = {-9'd80,-10'd280};
ram[22013] = {-9'd77,-10'd277};
ram[22014] = {-9'd74,-10'd274};
ram[22015] = {-9'd70,-10'd271};
ram[22016] = {-9'd70,-10'd271};
ram[22017] = {-9'd67,-10'd268};
ram[22018] = {-9'd64,-10'd264};
ram[22019] = {-9'd61,-10'd261};
ram[22020] = {-9'd58,-10'd258};
ram[22021] = {-9'd55,-10'd255};
ram[22022] = {-9'd52,-10'd252};
ram[22023] = {-9'd48,-10'd249};
ram[22024] = {-9'd45,-10'd246};
ram[22025] = {-9'd42,-10'd242};
ram[22026] = {-9'd39,-10'd239};
ram[22027] = {-9'd36,-10'd236};
ram[22028] = {-9'd33,-10'd233};
ram[22029] = {-9'd30,-10'd230};
ram[22030] = {-9'd26,-10'd227};
ram[22031] = {-9'd23,-10'd224};
ram[22032] = {-9'd20,-10'd220};
ram[22033] = {-9'd17,-10'd217};
ram[22034] = {-9'd14,-10'd214};
ram[22035] = {-9'd11,-10'd211};
ram[22036] = {-9'd8,-10'd208};
ram[22037] = {-9'd4,-10'd205};
ram[22038] = {-9'd1,-10'd202};
ram[22039] = {9'd2,-10'd198};
ram[22040] = {9'd5,-10'd195};
ram[22041] = {9'd8,-10'd192};
ram[22042] = {9'd11,-10'd189};
ram[22043] = {9'd14,-10'd186};
ram[22044] = {9'd18,-10'd183};
ram[22045] = {9'd21,-10'd180};
ram[22046] = {9'd24,-10'd176};
ram[22047] = {9'd27,-10'd173};
ram[22048] = {9'd30,-10'd170};
ram[22049] = {9'd33,-10'd167};
ram[22050] = {9'd36,-10'd164};
ram[22051] = {9'd40,-10'd161};
ram[22052] = {9'd43,-10'd158};
ram[22053] = {9'd46,-10'd154};
ram[22054] = {9'd49,-10'd151};
ram[22055] = {9'd52,-10'd148};
ram[22056] = {9'd55,-10'd145};
ram[22057] = {9'd58,-10'd142};
ram[22058] = {9'd62,-10'd139};
ram[22059] = {9'd65,-10'd136};
ram[22060] = {9'd68,-10'd132};
ram[22061] = {9'd71,-10'd129};
ram[22062] = {9'd74,-10'd126};
ram[22063] = {9'd77,-10'd123};
ram[22064] = {9'd80,-10'd120};
ram[22065] = {9'd84,-10'd117};
ram[22066] = {9'd87,-10'd114};
ram[22067] = {9'd90,-10'd110};
ram[22068] = {9'd93,-10'd107};
ram[22069] = {9'd96,-10'd104};
ram[22070] = {9'd99,-10'd101};
ram[22071] = {-9'd98,-10'd98};
ram[22072] = {-9'd95,-10'd95};
ram[22073] = {-9'd92,-10'd92};
ram[22074] = {-9'd88,-10'd88};
ram[22075] = {-9'd85,-10'd85};
ram[22076] = {-9'd82,-10'd82};
ram[22077] = {-9'd79,-10'd79};
ram[22078] = {-9'd76,-10'd76};
ram[22079] = {-9'd73,-10'd73};
ram[22080] = {-9'd70,-10'd70};
ram[22081] = {-9'd66,-10'd66};
ram[22082] = {-9'd63,-10'd63};
ram[22083] = {-9'd60,-10'd60};
ram[22084] = {-9'd57,-10'd57};
ram[22085] = {-9'd54,-10'd54};
ram[22086] = {-9'd51,-10'd51};
ram[22087] = {-9'd48,-10'd48};
ram[22088] = {-9'd44,-10'd44};
ram[22089] = {-9'd41,-10'd41};
ram[22090] = {-9'd38,-10'd38};
ram[22091] = {-9'd35,-10'd35};
ram[22092] = {-9'd32,-10'd32};
ram[22093] = {-9'd29,-10'd29};
ram[22094] = {-9'd26,-10'd26};
ram[22095] = {-9'd22,-10'd22};
ram[22096] = {-9'd19,-10'd19};
ram[22097] = {-9'd16,-10'd16};
ram[22098] = {-9'd13,-10'd13};
ram[22099] = {-9'd10,-10'd10};
ram[22100] = {-9'd7,-10'd7};
ram[22101] = {-9'd4,-10'd4};
ram[22102] = {9'd0,10'd0};
ram[22103] = {9'd3,10'd3};
ram[22104] = {9'd6,10'd6};
ram[22105] = {9'd9,10'd9};
ram[22106] = {9'd12,10'd12};
ram[22107] = {9'd15,10'd15};
ram[22108] = {9'd18,10'd18};
ram[22109] = {9'd21,10'd21};
ram[22110] = {9'd25,10'd25};
ram[22111] = {9'd28,10'd28};
ram[22112] = {9'd31,10'd31};
ram[22113] = {9'd34,10'd34};
ram[22114] = {9'd37,10'd37};
ram[22115] = {9'd40,10'd40};
ram[22116] = {9'd43,10'd43};
ram[22117] = {9'd47,10'd47};
ram[22118] = {9'd50,10'd50};
ram[22119] = {9'd53,10'd53};
ram[22120] = {9'd56,10'd56};
ram[22121] = {9'd59,10'd59};
ram[22122] = {9'd62,10'd62};
ram[22123] = {9'd65,10'd65};
ram[22124] = {9'd69,10'd69};
ram[22125] = {9'd72,10'd72};
ram[22126] = {9'd75,10'd75};
ram[22127] = {9'd78,10'd78};
ram[22128] = {9'd81,10'd81};
ram[22129] = {9'd84,10'd84};
ram[22130] = {9'd87,10'd87};
ram[22131] = {9'd91,10'd91};
ram[22132] = {9'd94,10'd94};
ram[22133] = {9'd97,10'd97};
ram[22134] = {-9'd100,10'd100};
ram[22135] = {-9'd97,10'd103};
ram[22136] = {-9'd94,10'd106};
ram[22137] = {-9'd91,10'd109};
ram[22138] = {-9'd88,10'd113};
ram[22139] = {-9'd85,10'd116};
ram[22140] = {-9'd81,10'd119};
ram[22141] = {-9'd78,10'd122};
ram[22142] = {-9'd75,10'd125};
ram[22143] = {-9'd72,10'd128};
ram[22144] = {-9'd72,10'd128};
ram[22145] = {-9'd69,10'd131};
ram[22146] = {-9'd66,10'd135};
ram[22147] = {-9'd63,10'd138};
ram[22148] = {-9'd59,10'd141};
ram[22149] = {-9'd56,10'd144};
ram[22150] = {-9'd53,10'd147};
ram[22151] = {-9'd50,10'd150};
ram[22152] = {-9'd47,10'd153};
ram[22153] = {-9'd44,10'd157};
ram[22154] = {-9'd41,10'd160};
ram[22155] = {-9'd37,10'd163};
ram[22156] = {-9'd34,10'd166};
ram[22157] = {-9'd31,10'd169};
ram[22158] = {-9'd28,10'd172};
ram[22159] = {-9'd25,10'd175};
ram[22160] = {-9'd22,10'd179};
ram[22161] = {-9'd19,10'd182};
ram[22162] = {-9'd15,10'd185};
ram[22163] = {-9'd12,10'd188};
ram[22164] = {-9'd9,10'd191};
ram[22165] = {-9'd6,10'd194};
ram[22166] = {-9'd3,10'd197};
ram[22167] = {9'd0,10'd201};
ram[22168] = {9'd3,10'd204};
ram[22169] = {9'd7,10'd207};
ram[22170] = {9'd10,10'd210};
ram[22171] = {9'd13,10'd213};
ram[22172] = {9'd16,10'd216};
ram[22173] = {9'd19,10'd219};
ram[22174] = {9'd22,10'd223};
ram[22175] = {9'd25,10'd226};
ram[22176] = {9'd29,10'd229};
ram[22177] = {9'd32,10'd232};
ram[22178] = {9'd35,10'd235};
ram[22179] = {9'd38,10'd238};
ram[22180] = {9'd41,10'd241};
ram[22181] = {9'd44,10'd245};
ram[22182] = {9'd47,10'd248};
ram[22183] = {9'd51,10'd251};
ram[22184] = {9'd54,10'd254};
ram[22185] = {9'd57,10'd257};
ram[22186] = {9'd60,10'd260};
ram[22187] = {9'd63,10'd263};
ram[22188] = {9'd66,10'd267};
ram[22189] = {9'd69,10'd270};
ram[22190] = {9'd73,10'd273};
ram[22191] = {9'd76,10'd276};
ram[22192] = {9'd79,10'd279};
ram[22193] = {9'd82,10'd282};
ram[22194] = {9'd85,10'd285};
ram[22195] = {9'd88,10'd289};
ram[22196] = {9'd91,10'd292};
ram[22197] = {9'd95,10'd295};
ram[22198] = {9'd98,10'd298};
ram[22199] = {-9'd99,10'd301};
ram[22200] = {-9'd96,10'd304};
ram[22201] = {-9'd93,10'd307};
ram[22202] = {-9'd90,10'd311};
ram[22203] = {-9'd87,10'd314};
ram[22204] = {-9'd84,10'd317};
ram[22205] = {-9'd81,10'd320};
ram[22206] = {-9'd77,10'd323};
ram[22207] = {-9'd74,10'd326};
ram[22208] = {-9'd71,10'd329};
ram[22209] = {-9'd68,10'd333};
ram[22210] = {-9'd65,10'd336};
ram[22211] = {-9'd62,10'd339};
ram[22212] = {-9'd59,10'd342};
ram[22213] = {-9'd55,10'd345};
ram[22214] = {-9'd52,10'd348};
ram[22215] = {-9'd49,10'd351};
ram[22216] = {-9'd46,10'd354};
ram[22217] = {-9'd43,10'd358};
ram[22218] = {-9'd40,10'd361};
ram[22219] = {-9'd37,10'd364};
ram[22220] = {-9'd33,10'd367};
ram[22221] = {-9'd30,10'd370};
ram[22222] = {-9'd27,10'd373};
ram[22223] = {-9'd24,10'd376};
ram[22224] = {-9'd21,10'd380};
ram[22225] = {-9'd18,10'd383};
ram[22226] = {-9'd15,10'd386};
ram[22227] = {-9'd11,10'd389};
ram[22228] = {-9'd8,10'd392};
ram[22229] = {-9'd5,10'd395};
ram[22230] = {-9'd2,10'd398};
ram[22231] = {9'd1,-10'd399};
ram[22232] = {9'd4,-10'd396};
ram[22233] = {9'd7,-10'd393};
ram[22234] = {9'd10,-10'd390};
ram[22235] = {9'd14,-10'd387};
ram[22236] = {9'd17,-10'd384};
ram[22237] = {9'd20,-10'd381};
ram[22238] = {9'd23,-10'd377};
ram[22239] = {9'd26,-10'd374};
ram[22240] = {9'd29,-10'd371};
ram[22241] = {9'd32,-10'd368};
ram[22242] = {9'd36,-10'd365};
ram[22243] = {9'd39,-10'd362};
ram[22244] = {9'd42,-10'd359};
ram[22245] = {9'd45,-10'd355};
ram[22246] = {9'd48,-10'd352};
ram[22247] = {9'd51,-10'd349};
ram[22248] = {9'd54,-10'd346};
ram[22249] = {9'd58,-10'd343};
ram[22250] = {9'd61,-10'd340};
ram[22251] = {9'd64,-10'd337};
ram[22252] = {9'd67,-10'd334};
ram[22253] = {9'd70,-10'd330};
ram[22254] = {9'd73,-10'd327};
ram[22255] = {9'd76,-10'd324};
ram[22256] = {9'd80,-10'd321};
ram[22257] = {9'd83,-10'd318};
ram[22258] = {9'd86,-10'd315};
ram[22259] = {9'd89,-10'd312};
ram[22260] = {9'd92,-10'd308};
ram[22261] = {9'd95,-10'd305};
ram[22262] = {9'd98,-10'd302};
ram[22263] = {-9'd99,-10'd299};
ram[22264] = {-9'd96,-10'd296};
ram[22265] = {-9'd92,-10'd293};
ram[22266] = {-9'd89,-10'd290};
ram[22267] = {-9'd86,-10'd286};
ram[22268] = {-9'd83,-10'd283};
ram[22269] = {-9'd80,-10'd280};
ram[22270] = {-9'd77,-10'd277};
ram[22271] = {-9'd74,-10'd274};
ram[22272] = {-9'd74,-10'd274};
ram[22273] = {-9'd70,-10'd271};
ram[22274] = {-9'd67,-10'd268};
ram[22275] = {-9'd64,-10'd264};
ram[22276] = {-9'd61,-10'd261};
ram[22277] = {-9'd58,-10'd258};
ram[22278] = {-9'd55,-10'd255};
ram[22279] = {-9'd52,-10'd252};
ram[22280] = {-9'd48,-10'd249};
ram[22281] = {-9'd45,-10'd246};
ram[22282] = {-9'd42,-10'd242};
ram[22283] = {-9'd39,-10'd239};
ram[22284] = {-9'd36,-10'd236};
ram[22285] = {-9'd33,-10'd233};
ram[22286] = {-9'd30,-10'd230};
ram[22287] = {-9'd26,-10'd227};
ram[22288] = {-9'd23,-10'd224};
ram[22289] = {-9'd20,-10'd220};
ram[22290] = {-9'd17,-10'd217};
ram[22291] = {-9'd14,-10'd214};
ram[22292] = {-9'd11,-10'd211};
ram[22293] = {-9'd8,-10'd208};
ram[22294] = {-9'd4,-10'd205};
ram[22295] = {-9'd1,-10'd202};
ram[22296] = {9'd2,-10'd198};
ram[22297] = {9'd5,-10'd195};
ram[22298] = {9'd8,-10'd192};
ram[22299] = {9'd11,-10'd189};
ram[22300] = {9'd14,-10'd186};
ram[22301] = {9'd18,-10'd183};
ram[22302] = {9'd21,-10'd180};
ram[22303] = {9'd24,-10'd176};
ram[22304] = {9'd27,-10'd173};
ram[22305] = {9'd30,-10'd170};
ram[22306] = {9'd33,-10'd167};
ram[22307] = {9'd36,-10'd164};
ram[22308] = {9'd40,-10'd161};
ram[22309] = {9'd43,-10'd158};
ram[22310] = {9'd46,-10'd154};
ram[22311] = {9'd49,-10'd151};
ram[22312] = {9'd52,-10'd148};
ram[22313] = {9'd55,-10'd145};
ram[22314] = {9'd58,-10'd142};
ram[22315] = {9'd62,-10'd139};
ram[22316] = {9'd65,-10'd136};
ram[22317] = {9'd68,-10'd132};
ram[22318] = {9'd71,-10'd129};
ram[22319] = {9'd74,-10'd126};
ram[22320] = {9'd77,-10'd123};
ram[22321] = {9'd80,-10'd120};
ram[22322] = {9'd84,-10'd117};
ram[22323] = {9'd87,-10'd114};
ram[22324] = {9'd90,-10'd110};
ram[22325] = {9'd93,-10'd107};
ram[22326] = {9'd96,-10'd104};
ram[22327] = {9'd99,-10'd101};
ram[22328] = {-9'd98,-10'd98};
ram[22329] = {-9'd95,-10'd95};
ram[22330] = {-9'd92,-10'd92};
ram[22331] = {-9'd88,-10'd88};
ram[22332] = {-9'd85,-10'd85};
ram[22333] = {-9'd82,-10'd82};
ram[22334] = {-9'd79,-10'd79};
ram[22335] = {-9'd76,-10'd76};
ram[22336] = {-9'd73,-10'd73};
ram[22337] = {-9'd70,-10'd70};
ram[22338] = {-9'd66,-10'd66};
ram[22339] = {-9'd63,-10'd63};
ram[22340] = {-9'd60,-10'd60};
ram[22341] = {-9'd57,-10'd57};
ram[22342] = {-9'd54,-10'd54};
ram[22343] = {-9'd51,-10'd51};
ram[22344] = {-9'd48,-10'd48};
ram[22345] = {-9'd44,-10'd44};
ram[22346] = {-9'd41,-10'd41};
ram[22347] = {-9'd38,-10'd38};
ram[22348] = {-9'd35,-10'd35};
ram[22349] = {-9'd32,-10'd32};
ram[22350] = {-9'd29,-10'd29};
ram[22351] = {-9'd26,-10'd26};
ram[22352] = {-9'd22,-10'd22};
ram[22353] = {-9'd19,-10'd19};
ram[22354] = {-9'd16,-10'd16};
ram[22355] = {-9'd13,-10'd13};
ram[22356] = {-9'd10,-10'd10};
ram[22357] = {-9'd7,-10'd7};
ram[22358] = {-9'd4,-10'd4};
ram[22359] = {9'd0,10'd0};
ram[22360] = {9'd3,10'd3};
ram[22361] = {9'd6,10'd6};
ram[22362] = {9'd9,10'd9};
ram[22363] = {9'd12,10'd12};
ram[22364] = {9'd15,10'd15};
ram[22365] = {9'd18,10'd18};
ram[22366] = {9'd21,10'd21};
ram[22367] = {9'd25,10'd25};
ram[22368] = {9'd28,10'd28};
ram[22369] = {9'd31,10'd31};
ram[22370] = {9'd34,10'd34};
ram[22371] = {9'd37,10'd37};
ram[22372] = {9'd40,10'd40};
ram[22373] = {9'd43,10'd43};
ram[22374] = {9'd47,10'd47};
ram[22375] = {9'd50,10'd50};
ram[22376] = {9'd53,10'd53};
ram[22377] = {9'd56,10'd56};
ram[22378] = {9'd59,10'd59};
ram[22379] = {9'd62,10'd62};
ram[22380] = {9'd65,10'd65};
ram[22381] = {9'd69,10'd69};
ram[22382] = {9'd72,10'd72};
ram[22383] = {9'd75,10'd75};
ram[22384] = {9'd78,10'd78};
ram[22385] = {9'd81,10'd81};
ram[22386] = {9'd84,10'd84};
ram[22387] = {9'd87,10'd87};
ram[22388] = {9'd91,10'd91};
ram[22389] = {9'd94,10'd94};
ram[22390] = {9'd97,10'd97};
ram[22391] = {-9'd100,10'd100};
ram[22392] = {-9'd97,10'd103};
ram[22393] = {-9'd94,10'd106};
ram[22394] = {-9'd91,10'd109};
ram[22395] = {-9'd88,10'd113};
ram[22396] = {-9'd85,10'd116};
ram[22397] = {-9'd81,10'd119};
ram[22398] = {-9'd78,10'd122};
ram[22399] = {-9'd75,10'd125};
ram[22400] = {-9'd75,10'd125};
ram[22401] = {-9'd72,10'd128};
ram[22402] = {-9'd69,10'd131};
ram[22403] = {-9'd66,10'd135};
ram[22404] = {-9'd63,10'd138};
ram[22405] = {-9'd59,10'd141};
ram[22406] = {-9'd56,10'd144};
ram[22407] = {-9'd53,10'd147};
ram[22408] = {-9'd50,10'd150};
ram[22409] = {-9'd47,10'd153};
ram[22410] = {-9'd44,10'd157};
ram[22411] = {-9'd41,10'd160};
ram[22412] = {-9'd37,10'd163};
ram[22413] = {-9'd34,10'd166};
ram[22414] = {-9'd31,10'd169};
ram[22415] = {-9'd28,10'd172};
ram[22416] = {-9'd25,10'd175};
ram[22417] = {-9'd22,10'd179};
ram[22418] = {-9'd19,10'd182};
ram[22419] = {-9'd15,10'd185};
ram[22420] = {-9'd12,10'd188};
ram[22421] = {-9'd9,10'd191};
ram[22422] = {-9'd6,10'd194};
ram[22423] = {-9'd3,10'd197};
ram[22424] = {9'd0,10'd201};
ram[22425] = {9'd3,10'd204};
ram[22426] = {9'd7,10'd207};
ram[22427] = {9'd10,10'd210};
ram[22428] = {9'd13,10'd213};
ram[22429] = {9'd16,10'd216};
ram[22430] = {9'd19,10'd219};
ram[22431] = {9'd22,10'd223};
ram[22432] = {9'd25,10'd226};
ram[22433] = {9'd29,10'd229};
ram[22434] = {9'd32,10'd232};
ram[22435] = {9'd35,10'd235};
ram[22436] = {9'd38,10'd238};
ram[22437] = {9'd41,10'd241};
ram[22438] = {9'd44,10'd245};
ram[22439] = {9'd47,10'd248};
ram[22440] = {9'd51,10'd251};
ram[22441] = {9'd54,10'd254};
ram[22442] = {9'd57,10'd257};
ram[22443] = {9'd60,10'd260};
ram[22444] = {9'd63,10'd263};
ram[22445] = {9'd66,10'd267};
ram[22446] = {9'd69,10'd270};
ram[22447] = {9'd73,10'd273};
ram[22448] = {9'd76,10'd276};
ram[22449] = {9'd79,10'd279};
ram[22450] = {9'd82,10'd282};
ram[22451] = {9'd85,10'd285};
ram[22452] = {9'd88,10'd289};
ram[22453] = {9'd91,10'd292};
ram[22454] = {9'd95,10'd295};
ram[22455] = {9'd98,10'd298};
ram[22456] = {-9'd99,10'd301};
ram[22457] = {-9'd96,10'd304};
ram[22458] = {-9'd93,10'd307};
ram[22459] = {-9'd90,10'd311};
ram[22460] = {-9'd87,10'd314};
ram[22461] = {-9'd84,10'd317};
ram[22462] = {-9'd81,10'd320};
ram[22463] = {-9'd77,10'd323};
ram[22464] = {-9'd74,10'd326};
ram[22465] = {-9'd71,10'd329};
ram[22466] = {-9'd68,10'd333};
ram[22467] = {-9'd65,10'd336};
ram[22468] = {-9'd62,10'd339};
ram[22469] = {-9'd59,10'd342};
ram[22470] = {-9'd55,10'd345};
ram[22471] = {-9'd52,10'd348};
ram[22472] = {-9'd49,10'd351};
ram[22473] = {-9'd46,10'd354};
ram[22474] = {-9'd43,10'd358};
ram[22475] = {-9'd40,10'd361};
ram[22476] = {-9'd37,10'd364};
ram[22477] = {-9'd33,10'd367};
ram[22478] = {-9'd30,10'd370};
ram[22479] = {-9'd27,10'd373};
ram[22480] = {-9'd24,10'd376};
ram[22481] = {-9'd21,10'd380};
ram[22482] = {-9'd18,10'd383};
ram[22483] = {-9'd15,10'd386};
ram[22484] = {-9'd11,10'd389};
ram[22485] = {-9'd8,10'd392};
ram[22486] = {-9'd5,10'd395};
ram[22487] = {-9'd2,10'd398};
ram[22488] = {9'd1,-10'd399};
ram[22489] = {9'd4,-10'd396};
ram[22490] = {9'd7,-10'd393};
ram[22491] = {9'd10,-10'd390};
ram[22492] = {9'd14,-10'd387};
ram[22493] = {9'd17,-10'd384};
ram[22494] = {9'd20,-10'd381};
ram[22495] = {9'd23,-10'd377};
ram[22496] = {9'd26,-10'd374};
ram[22497] = {9'd29,-10'd371};
ram[22498] = {9'd32,-10'd368};
ram[22499] = {9'd36,-10'd365};
ram[22500] = {9'd39,-10'd362};
ram[22501] = {9'd42,-10'd359};
ram[22502] = {9'd45,-10'd355};
ram[22503] = {9'd48,-10'd352};
ram[22504] = {9'd51,-10'd349};
ram[22505] = {9'd54,-10'd346};
ram[22506] = {9'd58,-10'd343};
ram[22507] = {9'd61,-10'd340};
ram[22508] = {9'd64,-10'd337};
ram[22509] = {9'd67,-10'd334};
ram[22510] = {9'd70,-10'd330};
ram[22511] = {9'd73,-10'd327};
ram[22512] = {9'd76,-10'd324};
ram[22513] = {9'd80,-10'd321};
ram[22514] = {9'd83,-10'd318};
ram[22515] = {9'd86,-10'd315};
ram[22516] = {9'd89,-10'd312};
ram[22517] = {9'd92,-10'd308};
ram[22518] = {9'd95,-10'd305};
ram[22519] = {9'd98,-10'd302};
ram[22520] = {-9'd99,-10'd299};
ram[22521] = {-9'd96,-10'd296};
ram[22522] = {-9'd92,-10'd293};
ram[22523] = {-9'd89,-10'd290};
ram[22524] = {-9'd86,-10'd286};
ram[22525] = {-9'd83,-10'd283};
ram[22526] = {-9'd80,-10'd280};
ram[22527] = {-9'd77,-10'd277};
ram[22528] = {-9'd77,-10'd277};
ram[22529] = {-9'd74,-10'd274};
ram[22530] = {-9'd70,-10'd271};
ram[22531] = {-9'd67,-10'd268};
ram[22532] = {-9'd64,-10'd264};
ram[22533] = {-9'd61,-10'd261};
ram[22534] = {-9'd58,-10'd258};
ram[22535] = {-9'd55,-10'd255};
ram[22536] = {-9'd52,-10'd252};
ram[22537] = {-9'd48,-10'd249};
ram[22538] = {-9'd45,-10'd246};
ram[22539] = {-9'd42,-10'd242};
ram[22540] = {-9'd39,-10'd239};
ram[22541] = {-9'd36,-10'd236};
ram[22542] = {-9'd33,-10'd233};
ram[22543] = {-9'd30,-10'd230};
ram[22544] = {-9'd26,-10'd227};
ram[22545] = {-9'd23,-10'd224};
ram[22546] = {-9'd20,-10'd220};
ram[22547] = {-9'd17,-10'd217};
ram[22548] = {-9'd14,-10'd214};
ram[22549] = {-9'd11,-10'd211};
ram[22550] = {-9'd8,-10'd208};
ram[22551] = {-9'd4,-10'd205};
ram[22552] = {-9'd1,-10'd202};
ram[22553] = {9'd2,-10'd198};
ram[22554] = {9'd5,-10'd195};
ram[22555] = {9'd8,-10'd192};
ram[22556] = {9'd11,-10'd189};
ram[22557] = {9'd14,-10'd186};
ram[22558] = {9'd18,-10'd183};
ram[22559] = {9'd21,-10'd180};
ram[22560] = {9'd24,-10'd176};
ram[22561] = {9'd27,-10'd173};
ram[22562] = {9'd30,-10'd170};
ram[22563] = {9'd33,-10'd167};
ram[22564] = {9'd36,-10'd164};
ram[22565] = {9'd40,-10'd161};
ram[22566] = {9'd43,-10'd158};
ram[22567] = {9'd46,-10'd154};
ram[22568] = {9'd49,-10'd151};
ram[22569] = {9'd52,-10'd148};
ram[22570] = {9'd55,-10'd145};
ram[22571] = {9'd58,-10'd142};
ram[22572] = {9'd62,-10'd139};
ram[22573] = {9'd65,-10'd136};
ram[22574] = {9'd68,-10'd132};
ram[22575] = {9'd71,-10'd129};
ram[22576] = {9'd74,-10'd126};
ram[22577] = {9'd77,-10'd123};
ram[22578] = {9'd80,-10'd120};
ram[22579] = {9'd84,-10'd117};
ram[22580] = {9'd87,-10'd114};
ram[22581] = {9'd90,-10'd110};
ram[22582] = {9'd93,-10'd107};
ram[22583] = {9'd96,-10'd104};
ram[22584] = {9'd99,-10'd101};
ram[22585] = {-9'd98,-10'd98};
ram[22586] = {-9'd95,-10'd95};
ram[22587] = {-9'd92,-10'd92};
ram[22588] = {-9'd88,-10'd88};
ram[22589] = {-9'd85,-10'd85};
ram[22590] = {-9'd82,-10'd82};
ram[22591] = {-9'd79,-10'd79};
ram[22592] = {-9'd76,-10'd76};
ram[22593] = {-9'd73,-10'd73};
ram[22594] = {-9'd70,-10'd70};
ram[22595] = {-9'd66,-10'd66};
ram[22596] = {-9'd63,-10'd63};
ram[22597] = {-9'd60,-10'd60};
ram[22598] = {-9'd57,-10'd57};
ram[22599] = {-9'd54,-10'd54};
ram[22600] = {-9'd51,-10'd51};
ram[22601] = {-9'd48,-10'd48};
ram[22602] = {-9'd44,-10'd44};
ram[22603] = {-9'd41,-10'd41};
ram[22604] = {-9'd38,-10'd38};
ram[22605] = {-9'd35,-10'd35};
ram[22606] = {-9'd32,-10'd32};
ram[22607] = {-9'd29,-10'd29};
ram[22608] = {-9'd26,-10'd26};
ram[22609] = {-9'd22,-10'd22};
ram[22610] = {-9'd19,-10'd19};
ram[22611] = {-9'd16,-10'd16};
ram[22612] = {-9'd13,-10'd13};
ram[22613] = {-9'd10,-10'd10};
ram[22614] = {-9'd7,-10'd7};
ram[22615] = {-9'd4,-10'd4};
ram[22616] = {9'd0,10'd0};
ram[22617] = {9'd3,10'd3};
ram[22618] = {9'd6,10'd6};
ram[22619] = {9'd9,10'd9};
ram[22620] = {9'd12,10'd12};
ram[22621] = {9'd15,10'd15};
ram[22622] = {9'd18,10'd18};
ram[22623] = {9'd21,10'd21};
ram[22624] = {9'd25,10'd25};
ram[22625] = {9'd28,10'd28};
ram[22626] = {9'd31,10'd31};
ram[22627] = {9'd34,10'd34};
ram[22628] = {9'd37,10'd37};
ram[22629] = {9'd40,10'd40};
ram[22630] = {9'd43,10'd43};
ram[22631] = {9'd47,10'd47};
ram[22632] = {9'd50,10'd50};
ram[22633] = {9'd53,10'd53};
ram[22634] = {9'd56,10'd56};
ram[22635] = {9'd59,10'd59};
ram[22636] = {9'd62,10'd62};
ram[22637] = {9'd65,10'd65};
ram[22638] = {9'd69,10'd69};
ram[22639] = {9'd72,10'd72};
ram[22640] = {9'd75,10'd75};
ram[22641] = {9'd78,10'd78};
ram[22642] = {9'd81,10'd81};
ram[22643] = {9'd84,10'd84};
ram[22644] = {9'd87,10'd87};
ram[22645] = {9'd91,10'd91};
ram[22646] = {9'd94,10'd94};
ram[22647] = {9'd97,10'd97};
ram[22648] = {-9'd100,10'd100};
ram[22649] = {-9'd97,10'd103};
ram[22650] = {-9'd94,10'd106};
ram[22651] = {-9'd91,10'd109};
ram[22652] = {-9'd88,10'd113};
ram[22653] = {-9'd85,10'd116};
ram[22654] = {-9'd81,10'd119};
ram[22655] = {-9'd78,10'd122};
ram[22656] = {-9'd78,10'd122};
ram[22657] = {-9'd75,10'd125};
ram[22658] = {-9'd72,10'd128};
ram[22659] = {-9'd69,10'd131};
ram[22660] = {-9'd66,10'd135};
ram[22661] = {-9'd63,10'd138};
ram[22662] = {-9'd59,10'd141};
ram[22663] = {-9'd56,10'd144};
ram[22664] = {-9'd53,10'd147};
ram[22665] = {-9'd50,10'd150};
ram[22666] = {-9'd47,10'd153};
ram[22667] = {-9'd44,10'd157};
ram[22668] = {-9'd41,10'd160};
ram[22669] = {-9'd37,10'd163};
ram[22670] = {-9'd34,10'd166};
ram[22671] = {-9'd31,10'd169};
ram[22672] = {-9'd28,10'd172};
ram[22673] = {-9'd25,10'd175};
ram[22674] = {-9'd22,10'd179};
ram[22675] = {-9'd19,10'd182};
ram[22676] = {-9'd15,10'd185};
ram[22677] = {-9'd12,10'd188};
ram[22678] = {-9'd9,10'd191};
ram[22679] = {-9'd6,10'd194};
ram[22680] = {-9'd3,10'd197};
ram[22681] = {9'd0,10'd201};
ram[22682] = {9'd3,10'd204};
ram[22683] = {9'd7,10'd207};
ram[22684] = {9'd10,10'd210};
ram[22685] = {9'd13,10'd213};
ram[22686] = {9'd16,10'd216};
ram[22687] = {9'd19,10'd219};
ram[22688] = {9'd22,10'd223};
ram[22689] = {9'd25,10'd226};
ram[22690] = {9'd29,10'd229};
ram[22691] = {9'd32,10'd232};
ram[22692] = {9'd35,10'd235};
ram[22693] = {9'd38,10'd238};
ram[22694] = {9'd41,10'd241};
ram[22695] = {9'd44,10'd245};
ram[22696] = {9'd47,10'd248};
ram[22697] = {9'd51,10'd251};
ram[22698] = {9'd54,10'd254};
ram[22699] = {9'd57,10'd257};
ram[22700] = {9'd60,10'd260};
ram[22701] = {9'd63,10'd263};
ram[22702] = {9'd66,10'd267};
ram[22703] = {9'd69,10'd270};
ram[22704] = {9'd73,10'd273};
ram[22705] = {9'd76,10'd276};
ram[22706] = {9'd79,10'd279};
ram[22707] = {9'd82,10'd282};
ram[22708] = {9'd85,10'd285};
ram[22709] = {9'd88,10'd289};
ram[22710] = {9'd91,10'd292};
ram[22711] = {9'd95,10'd295};
ram[22712] = {9'd98,10'd298};
ram[22713] = {-9'd99,10'd301};
ram[22714] = {-9'd96,10'd304};
ram[22715] = {-9'd93,10'd307};
ram[22716] = {-9'd90,10'd311};
ram[22717] = {-9'd87,10'd314};
ram[22718] = {-9'd84,10'd317};
ram[22719] = {-9'd81,10'd320};
ram[22720] = {-9'd77,10'd323};
ram[22721] = {-9'd74,10'd326};
ram[22722] = {-9'd71,10'd329};
ram[22723] = {-9'd68,10'd333};
ram[22724] = {-9'd65,10'd336};
ram[22725] = {-9'd62,10'd339};
ram[22726] = {-9'd59,10'd342};
ram[22727] = {-9'd55,10'd345};
ram[22728] = {-9'd52,10'd348};
ram[22729] = {-9'd49,10'd351};
ram[22730] = {-9'd46,10'd354};
ram[22731] = {-9'd43,10'd358};
ram[22732] = {-9'd40,10'd361};
ram[22733] = {-9'd37,10'd364};
ram[22734] = {-9'd33,10'd367};
ram[22735] = {-9'd30,10'd370};
ram[22736] = {-9'd27,10'd373};
ram[22737] = {-9'd24,10'd376};
ram[22738] = {-9'd21,10'd380};
ram[22739] = {-9'd18,10'd383};
ram[22740] = {-9'd15,10'd386};
ram[22741] = {-9'd11,10'd389};
ram[22742] = {-9'd8,10'd392};
ram[22743] = {-9'd5,10'd395};
ram[22744] = {-9'd2,10'd398};
ram[22745] = {9'd1,-10'd399};
ram[22746] = {9'd4,-10'd396};
ram[22747] = {9'd7,-10'd393};
ram[22748] = {9'd10,-10'd390};
ram[22749] = {9'd14,-10'd387};
ram[22750] = {9'd17,-10'd384};
ram[22751] = {9'd20,-10'd381};
ram[22752] = {9'd23,-10'd377};
ram[22753] = {9'd26,-10'd374};
ram[22754] = {9'd29,-10'd371};
ram[22755] = {9'd32,-10'd368};
ram[22756] = {9'd36,-10'd365};
ram[22757] = {9'd39,-10'd362};
ram[22758] = {9'd42,-10'd359};
ram[22759] = {9'd45,-10'd355};
ram[22760] = {9'd48,-10'd352};
ram[22761] = {9'd51,-10'd349};
ram[22762] = {9'd54,-10'd346};
ram[22763] = {9'd58,-10'd343};
ram[22764] = {9'd61,-10'd340};
ram[22765] = {9'd64,-10'd337};
ram[22766] = {9'd67,-10'd334};
ram[22767] = {9'd70,-10'd330};
ram[22768] = {9'd73,-10'd327};
ram[22769] = {9'd76,-10'd324};
ram[22770] = {9'd80,-10'd321};
ram[22771] = {9'd83,-10'd318};
ram[22772] = {9'd86,-10'd315};
ram[22773] = {9'd89,-10'd312};
ram[22774] = {9'd92,-10'd308};
ram[22775] = {9'd95,-10'd305};
ram[22776] = {9'd98,-10'd302};
ram[22777] = {-9'd99,-10'd299};
ram[22778] = {-9'd96,-10'd296};
ram[22779] = {-9'd92,-10'd293};
ram[22780] = {-9'd89,-10'd290};
ram[22781] = {-9'd86,-10'd286};
ram[22782] = {-9'd83,-10'd283};
ram[22783] = {-9'd80,-10'd280};
ram[22784] = {-9'd80,-10'd280};
ram[22785] = {-9'd77,-10'd277};
ram[22786] = {-9'd74,-10'd274};
ram[22787] = {-9'd70,-10'd271};
ram[22788] = {-9'd67,-10'd268};
ram[22789] = {-9'd64,-10'd264};
ram[22790] = {-9'd61,-10'd261};
ram[22791] = {-9'd58,-10'd258};
ram[22792] = {-9'd55,-10'd255};
ram[22793] = {-9'd52,-10'd252};
ram[22794] = {-9'd48,-10'd249};
ram[22795] = {-9'd45,-10'd246};
ram[22796] = {-9'd42,-10'd242};
ram[22797] = {-9'd39,-10'd239};
ram[22798] = {-9'd36,-10'd236};
ram[22799] = {-9'd33,-10'd233};
ram[22800] = {-9'd30,-10'd230};
ram[22801] = {-9'd26,-10'd227};
ram[22802] = {-9'd23,-10'd224};
ram[22803] = {-9'd20,-10'd220};
ram[22804] = {-9'd17,-10'd217};
ram[22805] = {-9'd14,-10'd214};
ram[22806] = {-9'd11,-10'd211};
ram[22807] = {-9'd8,-10'd208};
ram[22808] = {-9'd4,-10'd205};
ram[22809] = {-9'd1,-10'd202};
ram[22810] = {9'd2,-10'd198};
ram[22811] = {9'd5,-10'd195};
ram[22812] = {9'd8,-10'd192};
ram[22813] = {9'd11,-10'd189};
ram[22814] = {9'd14,-10'd186};
ram[22815] = {9'd18,-10'd183};
ram[22816] = {9'd21,-10'd180};
ram[22817] = {9'd24,-10'd176};
ram[22818] = {9'd27,-10'd173};
ram[22819] = {9'd30,-10'd170};
ram[22820] = {9'd33,-10'd167};
ram[22821] = {9'd36,-10'd164};
ram[22822] = {9'd40,-10'd161};
ram[22823] = {9'd43,-10'd158};
ram[22824] = {9'd46,-10'd154};
ram[22825] = {9'd49,-10'd151};
ram[22826] = {9'd52,-10'd148};
ram[22827] = {9'd55,-10'd145};
ram[22828] = {9'd58,-10'd142};
ram[22829] = {9'd62,-10'd139};
ram[22830] = {9'd65,-10'd136};
ram[22831] = {9'd68,-10'd132};
ram[22832] = {9'd71,-10'd129};
ram[22833] = {9'd74,-10'd126};
ram[22834] = {9'd77,-10'd123};
ram[22835] = {9'd80,-10'd120};
ram[22836] = {9'd84,-10'd117};
ram[22837] = {9'd87,-10'd114};
ram[22838] = {9'd90,-10'd110};
ram[22839] = {9'd93,-10'd107};
ram[22840] = {9'd96,-10'd104};
ram[22841] = {9'd99,-10'd101};
ram[22842] = {-9'd98,-10'd98};
ram[22843] = {-9'd95,-10'd95};
ram[22844] = {-9'd92,-10'd92};
ram[22845] = {-9'd88,-10'd88};
ram[22846] = {-9'd85,-10'd85};
ram[22847] = {-9'd82,-10'd82};
ram[22848] = {-9'd79,-10'd79};
ram[22849] = {-9'd76,-10'd76};
ram[22850] = {-9'd73,-10'd73};
ram[22851] = {-9'd70,-10'd70};
ram[22852] = {-9'd66,-10'd66};
ram[22853] = {-9'd63,-10'd63};
ram[22854] = {-9'd60,-10'd60};
ram[22855] = {-9'd57,-10'd57};
ram[22856] = {-9'd54,-10'd54};
ram[22857] = {-9'd51,-10'd51};
ram[22858] = {-9'd48,-10'd48};
ram[22859] = {-9'd44,-10'd44};
ram[22860] = {-9'd41,-10'd41};
ram[22861] = {-9'd38,-10'd38};
ram[22862] = {-9'd35,-10'd35};
ram[22863] = {-9'd32,-10'd32};
ram[22864] = {-9'd29,-10'd29};
ram[22865] = {-9'd26,-10'd26};
ram[22866] = {-9'd22,-10'd22};
ram[22867] = {-9'd19,-10'd19};
ram[22868] = {-9'd16,-10'd16};
ram[22869] = {-9'd13,-10'd13};
ram[22870] = {-9'd10,-10'd10};
ram[22871] = {-9'd7,-10'd7};
ram[22872] = {-9'd4,-10'd4};
ram[22873] = {9'd0,10'd0};
ram[22874] = {9'd3,10'd3};
ram[22875] = {9'd6,10'd6};
ram[22876] = {9'd9,10'd9};
ram[22877] = {9'd12,10'd12};
ram[22878] = {9'd15,10'd15};
ram[22879] = {9'd18,10'd18};
ram[22880] = {9'd21,10'd21};
ram[22881] = {9'd25,10'd25};
ram[22882] = {9'd28,10'd28};
ram[22883] = {9'd31,10'd31};
ram[22884] = {9'd34,10'd34};
ram[22885] = {9'd37,10'd37};
ram[22886] = {9'd40,10'd40};
ram[22887] = {9'd43,10'd43};
ram[22888] = {9'd47,10'd47};
ram[22889] = {9'd50,10'd50};
ram[22890] = {9'd53,10'd53};
ram[22891] = {9'd56,10'd56};
ram[22892] = {9'd59,10'd59};
ram[22893] = {9'd62,10'd62};
ram[22894] = {9'd65,10'd65};
ram[22895] = {9'd69,10'd69};
ram[22896] = {9'd72,10'd72};
ram[22897] = {9'd75,10'd75};
ram[22898] = {9'd78,10'd78};
ram[22899] = {9'd81,10'd81};
ram[22900] = {9'd84,10'd84};
ram[22901] = {9'd87,10'd87};
ram[22902] = {9'd91,10'd91};
ram[22903] = {9'd94,10'd94};
ram[22904] = {9'd97,10'd97};
ram[22905] = {-9'd100,10'd100};
ram[22906] = {-9'd97,10'd103};
ram[22907] = {-9'd94,10'd106};
ram[22908] = {-9'd91,10'd109};
ram[22909] = {-9'd88,10'd113};
ram[22910] = {-9'd85,10'd116};
ram[22911] = {-9'd81,10'd119};
ram[22912] = {-9'd81,10'd119};
ram[22913] = {-9'd78,10'd122};
ram[22914] = {-9'd75,10'd125};
ram[22915] = {-9'd72,10'd128};
ram[22916] = {-9'd69,10'd131};
ram[22917] = {-9'd66,10'd135};
ram[22918] = {-9'd63,10'd138};
ram[22919] = {-9'd59,10'd141};
ram[22920] = {-9'd56,10'd144};
ram[22921] = {-9'd53,10'd147};
ram[22922] = {-9'd50,10'd150};
ram[22923] = {-9'd47,10'd153};
ram[22924] = {-9'd44,10'd157};
ram[22925] = {-9'd41,10'd160};
ram[22926] = {-9'd37,10'd163};
ram[22927] = {-9'd34,10'd166};
ram[22928] = {-9'd31,10'd169};
ram[22929] = {-9'd28,10'd172};
ram[22930] = {-9'd25,10'd175};
ram[22931] = {-9'd22,10'd179};
ram[22932] = {-9'd19,10'd182};
ram[22933] = {-9'd15,10'd185};
ram[22934] = {-9'd12,10'd188};
ram[22935] = {-9'd9,10'd191};
ram[22936] = {-9'd6,10'd194};
ram[22937] = {-9'd3,10'd197};
ram[22938] = {9'd0,10'd201};
ram[22939] = {9'd3,10'd204};
ram[22940] = {9'd7,10'd207};
ram[22941] = {9'd10,10'd210};
ram[22942] = {9'd13,10'd213};
ram[22943] = {9'd16,10'd216};
ram[22944] = {9'd19,10'd219};
ram[22945] = {9'd22,10'd223};
ram[22946] = {9'd25,10'd226};
ram[22947] = {9'd29,10'd229};
ram[22948] = {9'd32,10'd232};
ram[22949] = {9'd35,10'd235};
ram[22950] = {9'd38,10'd238};
ram[22951] = {9'd41,10'd241};
ram[22952] = {9'd44,10'd245};
ram[22953] = {9'd47,10'd248};
ram[22954] = {9'd51,10'd251};
ram[22955] = {9'd54,10'd254};
ram[22956] = {9'd57,10'd257};
ram[22957] = {9'd60,10'd260};
ram[22958] = {9'd63,10'd263};
ram[22959] = {9'd66,10'd267};
ram[22960] = {9'd69,10'd270};
ram[22961] = {9'd73,10'd273};
ram[22962] = {9'd76,10'd276};
ram[22963] = {9'd79,10'd279};
ram[22964] = {9'd82,10'd282};
ram[22965] = {9'd85,10'd285};
ram[22966] = {9'd88,10'd289};
ram[22967] = {9'd91,10'd292};
ram[22968] = {9'd95,10'd295};
ram[22969] = {9'd98,10'd298};
ram[22970] = {-9'd99,10'd301};
ram[22971] = {-9'd96,10'd304};
ram[22972] = {-9'd93,10'd307};
ram[22973] = {-9'd90,10'd311};
ram[22974] = {-9'd87,10'd314};
ram[22975] = {-9'd84,10'd317};
ram[22976] = {-9'd81,10'd320};
ram[22977] = {-9'd77,10'd323};
ram[22978] = {-9'd74,10'd326};
ram[22979] = {-9'd71,10'd329};
ram[22980] = {-9'd68,10'd333};
ram[22981] = {-9'd65,10'd336};
ram[22982] = {-9'd62,10'd339};
ram[22983] = {-9'd59,10'd342};
ram[22984] = {-9'd55,10'd345};
ram[22985] = {-9'd52,10'd348};
ram[22986] = {-9'd49,10'd351};
ram[22987] = {-9'd46,10'd354};
ram[22988] = {-9'd43,10'd358};
ram[22989] = {-9'd40,10'd361};
ram[22990] = {-9'd37,10'd364};
ram[22991] = {-9'd33,10'd367};
ram[22992] = {-9'd30,10'd370};
ram[22993] = {-9'd27,10'd373};
ram[22994] = {-9'd24,10'd376};
ram[22995] = {-9'd21,10'd380};
ram[22996] = {-9'd18,10'd383};
ram[22997] = {-9'd15,10'd386};
ram[22998] = {-9'd11,10'd389};
ram[22999] = {-9'd8,10'd392};
ram[23000] = {-9'd5,10'd395};
ram[23001] = {-9'd2,10'd398};
ram[23002] = {9'd1,-10'd399};
ram[23003] = {9'd4,-10'd396};
ram[23004] = {9'd7,-10'd393};
ram[23005] = {9'd10,-10'd390};
ram[23006] = {9'd14,-10'd387};
ram[23007] = {9'd17,-10'd384};
ram[23008] = {9'd20,-10'd381};
ram[23009] = {9'd23,-10'd377};
ram[23010] = {9'd26,-10'd374};
ram[23011] = {9'd29,-10'd371};
ram[23012] = {9'd32,-10'd368};
ram[23013] = {9'd36,-10'd365};
ram[23014] = {9'd39,-10'd362};
ram[23015] = {9'd42,-10'd359};
ram[23016] = {9'd45,-10'd355};
ram[23017] = {9'd48,-10'd352};
ram[23018] = {9'd51,-10'd349};
ram[23019] = {9'd54,-10'd346};
ram[23020] = {9'd58,-10'd343};
ram[23021] = {9'd61,-10'd340};
ram[23022] = {9'd64,-10'd337};
ram[23023] = {9'd67,-10'd334};
ram[23024] = {9'd70,-10'd330};
ram[23025] = {9'd73,-10'd327};
ram[23026] = {9'd76,-10'd324};
ram[23027] = {9'd80,-10'd321};
ram[23028] = {9'd83,-10'd318};
ram[23029] = {9'd86,-10'd315};
ram[23030] = {9'd89,-10'd312};
ram[23031] = {9'd92,-10'd308};
ram[23032] = {9'd95,-10'd305};
ram[23033] = {9'd98,-10'd302};
ram[23034] = {-9'd99,-10'd299};
ram[23035] = {-9'd96,-10'd296};
ram[23036] = {-9'd92,-10'd293};
ram[23037] = {-9'd89,-10'd290};
ram[23038] = {-9'd86,-10'd286};
ram[23039] = {-9'd83,-10'd283};
ram[23040] = {-9'd83,-10'd283};
ram[23041] = {-9'd80,-10'd280};
ram[23042] = {-9'd77,-10'd277};
ram[23043] = {-9'd74,-10'd274};
ram[23044] = {-9'd70,-10'd271};
ram[23045] = {-9'd67,-10'd268};
ram[23046] = {-9'd64,-10'd264};
ram[23047] = {-9'd61,-10'd261};
ram[23048] = {-9'd58,-10'd258};
ram[23049] = {-9'd55,-10'd255};
ram[23050] = {-9'd52,-10'd252};
ram[23051] = {-9'd48,-10'd249};
ram[23052] = {-9'd45,-10'd246};
ram[23053] = {-9'd42,-10'd242};
ram[23054] = {-9'd39,-10'd239};
ram[23055] = {-9'd36,-10'd236};
ram[23056] = {-9'd33,-10'd233};
ram[23057] = {-9'd30,-10'd230};
ram[23058] = {-9'd26,-10'd227};
ram[23059] = {-9'd23,-10'd224};
ram[23060] = {-9'd20,-10'd220};
ram[23061] = {-9'd17,-10'd217};
ram[23062] = {-9'd14,-10'd214};
ram[23063] = {-9'd11,-10'd211};
ram[23064] = {-9'd8,-10'd208};
ram[23065] = {-9'd4,-10'd205};
ram[23066] = {-9'd1,-10'd202};
ram[23067] = {9'd2,-10'd198};
ram[23068] = {9'd5,-10'd195};
ram[23069] = {9'd8,-10'd192};
ram[23070] = {9'd11,-10'd189};
ram[23071] = {9'd14,-10'd186};
ram[23072] = {9'd18,-10'd183};
ram[23073] = {9'd21,-10'd180};
ram[23074] = {9'd24,-10'd176};
ram[23075] = {9'd27,-10'd173};
ram[23076] = {9'd30,-10'd170};
ram[23077] = {9'd33,-10'd167};
ram[23078] = {9'd36,-10'd164};
ram[23079] = {9'd40,-10'd161};
ram[23080] = {9'd43,-10'd158};
ram[23081] = {9'd46,-10'd154};
ram[23082] = {9'd49,-10'd151};
ram[23083] = {9'd52,-10'd148};
ram[23084] = {9'd55,-10'd145};
ram[23085] = {9'd58,-10'd142};
ram[23086] = {9'd62,-10'd139};
ram[23087] = {9'd65,-10'd136};
ram[23088] = {9'd68,-10'd132};
ram[23089] = {9'd71,-10'd129};
ram[23090] = {9'd74,-10'd126};
ram[23091] = {9'd77,-10'd123};
ram[23092] = {9'd80,-10'd120};
ram[23093] = {9'd84,-10'd117};
ram[23094] = {9'd87,-10'd114};
ram[23095] = {9'd90,-10'd110};
ram[23096] = {9'd93,-10'd107};
ram[23097] = {9'd96,-10'd104};
ram[23098] = {9'd99,-10'd101};
ram[23099] = {-9'd98,-10'd98};
ram[23100] = {-9'd95,-10'd95};
ram[23101] = {-9'd92,-10'd92};
ram[23102] = {-9'd88,-10'd88};
ram[23103] = {-9'd85,-10'd85};
ram[23104] = {-9'd82,-10'd82};
ram[23105] = {-9'd79,-10'd79};
ram[23106] = {-9'd76,-10'd76};
ram[23107] = {-9'd73,-10'd73};
ram[23108] = {-9'd70,-10'd70};
ram[23109] = {-9'd66,-10'd66};
ram[23110] = {-9'd63,-10'd63};
ram[23111] = {-9'd60,-10'd60};
ram[23112] = {-9'd57,-10'd57};
ram[23113] = {-9'd54,-10'd54};
ram[23114] = {-9'd51,-10'd51};
ram[23115] = {-9'd48,-10'd48};
ram[23116] = {-9'd44,-10'd44};
ram[23117] = {-9'd41,-10'd41};
ram[23118] = {-9'd38,-10'd38};
ram[23119] = {-9'd35,-10'd35};
ram[23120] = {-9'd32,-10'd32};
ram[23121] = {-9'd29,-10'd29};
ram[23122] = {-9'd26,-10'd26};
ram[23123] = {-9'd22,-10'd22};
ram[23124] = {-9'd19,-10'd19};
ram[23125] = {-9'd16,-10'd16};
ram[23126] = {-9'd13,-10'd13};
ram[23127] = {-9'd10,-10'd10};
ram[23128] = {-9'd7,-10'd7};
ram[23129] = {-9'd4,-10'd4};
ram[23130] = {9'd0,10'd0};
ram[23131] = {9'd3,10'd3};
ram[23132] = {9'd6,10'd6};
ram[23133] = {9'd9,10'd9};
ram[23134] = {9'd12,10'd12};
ram[23135] = {9'd15,10'd15};
ram[23136] = {9'd18,10'd18};
ram[23137] = {9'd21,10'd21};
ram[23138] = {9'd25,10'd25};
ram[23139] = {9'd28,10'd28};
ram[23140] = {9'd31,10'd31};
ram[23141] = {9'd34,10'd34};
ram[23142] = {9'd37,10'd37};
ram[23143] = {9'd40,10'd40};
ram[23144] = {9'd43,10'd43};
ram[23145] = {9'd47,10'd47};
ram[23146] = {9'd50,10'd50};
ram[23147] = {9'd53,10'd53};
ram[23148] = {9'd56,10'd56};
ram[23149] = {9'd59,10'd59};
ram[23150] = {9'd62,10'd62};
ram[23151] = {9'd65,10'd65};
ram[23152] = {9'd69,10'd69};
ram[23153] = {9'd72,10'd72};
ram[23154] = {9'd75,10'd75};
ram[23155] = {9'd78,10'd78};
ram[23156] = {9'd81,10'd81};
ram[23157] = {9'd84,10'd84};
ram[23158] = {9'd87,10'd87};
ram[23159] = {9'd91,10'd91};
ram[23160] = {9'd94,10'd94};
ram[23161] = {9'd97,10'd97};
ram[23162] = {-9'd100,10'd100};
ram[23163] = {-9'd97,10'd103};
ram[23164] = {-9'd94,10'd106};
ram[23165] = {-9'd91,10'd109};
ram[23166] = {-9'd88,10'd113};
ram[23167] = {-9'd85,10'd116};
ram[23168] = {-9'd85,10'd116};
ram[23169] = {-9'd81,10'd119};
ram[23170] = {-9'd78,10'd122};
ram[23171] = {-9'd75,10'd125};
ram[23172] = {-9'd72,10'd128};
ram[23173] = {-9'd69,10'd131};
ram[23174] = {-9'd66,10'd135};
ram[23175] = {-9'd63,10'd138};
ram[23176] = {-9'd59,10'd141};
ram[23177] = {-9'd56,10'd144};
ram[23178] = {-9'd53,10'd147};
ram[23179] = {-9'd50,10'd150};
ram[23180] = {-9'd47,10'd153};
ram[23181] = {-9'd44,10'd157};
ram[23182] = {-9'd41,10'd160};
ram[23183] = {-9'd37,10'd163};
ram[23184] = {-9'd34,10'd166};
ram[23185] = {-9'd31,10'd169};
ram[23186] = {-9'd28,10'd172};
ram[23187] = {-9'd25,10'd175};
ram[23188] = {-9'd22,10'd179};
ram[23189] = {-9'd19,10'd182};
ram[23190] = {-9'd15,10'd185};
ram[23191] = {-9'd12,10'd188};
ram[23192] = {-9'd9,10'd191};
ram[23193] = {-9'd6,10'd194};
ram[23194] = {-9'd3,10'd197};
ram[23195] = {9'd0,10'd201};
ram[23196] = {9'd3,10'd204};
ram[23197] = {9'd7,10'd207};
ram[23198] = {9'd10,10'd210};
ram[23199] = {9'd13,10'd213};
ram[23200] = {9'd16,10'd216};
ram[23201] = {9'd19,10'd219};
ram[23202] = {9'd22,10'd223};
ram[23203] = {9'd25,10'd226};
ram[23204] = {9'd29,10'd229};
ram[23205] = {9'd32,10'd232};
ram[23206] = {9'd35,10'd235};
ram[23207] = {9'd38,10'd238};
ram[23208] = {9'd41,10'd241};
ram[23209] = {9'd44,10'd245};
ram[23210] = {9'd47,10'd248};
ram[23211] = {9'd51,10'd251};
ram[23212] = {9'd54,10'd254};
ram[23213] = {9'd57,10'd257};
ram[23214] = {9'd60,10'd260};
ram[23215] = {9'd63,10'd263};
ram[23216] = {9'd66,10'd267};
ram[23217] = {9'd69,10'd270};
ram[23218] = {9'd73,10'd273};
ram[23219] = {9'd76,10'd276};
ram[23220] = {9'd79,10'd279};
ram[23221] = {9'd82,10'd282};
ram[23222] = {9'd85,10'd285};
ram[23223] = {9'd88,10'd289};
ram[23224] = {9'd91,10'd292};
ram[23225] = {9'd95,10'd295};
ram[23226] = {9'd98,10'd298};
ram[23227] = {-9'd99,10'd301};
ram[23228] = {-9'd96,10'd304};
ram[23229] = {-9'd93,10'd307};
ram[23230] = {-9'd90,10'd311};
ram[23231] = {-9'd87,10'd314};
ram[23232] = {-9'd84,10'd317};
ram[23233] = {-9'd81,10'd320};
ram[23234] = {-9'd77,10'd323};
ram[23235] = {-9'd74,10'd326};
ram[23236] = {-9'd71,10'd329};
ram[23237] = {-9'd68,10'd333};
ram[23238] = {-9'd65,10'd336};
ram[23239] = {-9'd62,10'd339};
ram[23240] = {-9'd59,10'd342};
ram[23241] = {-9'd55,10'd345};
ram[23242] = {-9'd52,10'd348};
ram[23243] = {-9'd49,10'd351};
ram[23244] = {-9'd46,10'd354};
ram[23245] = {-9'd43,10'd358};
ram[23246] = {-9'd40,10'd361};
ram[23247] = {-9'd37,10'd364};
ram[23248] = {-9'd33,10'd367};
ram[23249] = {-9'd30,10'd370};
ram[23250] = {-9'd27,10'd373};
ram[23251] = {-9'd24,10'd376};
ram[23252] = {-9'd21,10'd380};
ram[23253] = {-9'd18,10'd383};
ram[23254] = {-9'd15,10'd386};
ram[23255] = {-9'd11,10'd389};
ram[23256] = {-9'd8,10'd392};
ram[23257] = {-9'd5,10'd395};
ram[23258] = {-9'd2,10'd398};
ram[23259] = {9'd1,-10'd399};
ram[23260] = {9'd4,-10'd396};
ram[23261] = {9'd7,-10'd393};
ram[23262] = {9'd10,-10'd390};
ram[23263] = {9'd14,-10'd387};
ram[23264] = {9'd17,-10'd384};
ram[23265] = {9'd20,-10'd381};
ram[23266] = {9'd23,-10'd377};
ram[23267] = {9'd26,-10'd374};
ram[23268] = {9'd29,-10'd371};
ram[23269] = {9'd32,-10'd368};
ram[23270] = {9'd36,-10'd365};
ram[23271] = {9'd39,-10'd362};
ram[23272] = {9'd42,-10'd359};
ram[23273] = {9'd45,-10'd355};
ram[23274] = {9'd48,-10'd352};
ram[23275] = {9'd51,-10'd349};
ram[23276] = {9'd54,-10'd346};
ram[23277] = {9'd58,-10'd343};
ram[23278] = {9'd61,-10'd340};
ram[23279] = {9'd64,-10'd337};
ram[23280] = {9'd67,-10'd334};
ram[23281] = {9'd70,-10'd330};
ram[23282] = {9'd73,-10'd327};
ram[23283] = {9'd76,-10'd324};
ram[23284] = {9'd80,-10'd321};
ram[23285] = {9'd83,-10'd318};
ram[23286] = {9'd86,-10'd315};
ram[23287] = {9'd89,-10'd312};
ram[23288] = {9'd92,-10'd308};
ram[23289] = {9'd95,-10'd305};
ram[23290] = {9'd98,-10'd302};
ram[23291] = {-9'd99,-10'd299};
ram[23292] = {-9'd96,-10'd296};
ram[23293] = {-9'd92,-10'd293};
ram[23294] = {-9'd89,-10'd290};
ram[23295] = {-9'd86,-10'd286};
ram[23296] = {-9'd86,-10'd286};
ram[23297] = {-9'd83,-10'd283};
ram[23298] = {-9'd80,-10'd280};
ram[23299] = {-9'd77,-10'd277};
ram[23300] = {-9'd74,-10'd274};
ram[23301] = {-9'd70,-10'd271};
ram[23302] = {-9'd67,-10'd268};
ram[23303] = {-9'd64,-10'd264};
ram[23304] = {-9'd61,-10'd261};
ram[23305] = {-9'd58,-10'd258};
ram[23306] = {-9'd55,-10'd255};
ram[23307] = {-9'd52,-10'd252};
ram[23308] = {-9'd48,-10'd249};
ram[23309] = {-9'd45,-10'd246};
ram[23310] = {-9'd42,-10'd242};
ram[23311] = {-9'd39,-10'd239};
ram[23312] = {-9'd36,-10'd236};
ram[23313] = {-9'd33,-10'd233};
ram[23314] = {-9'd30,-10'd230};
ram[23315] = {-9'd26,-10'd227};
ram[23316] = {-9'd23,-10'd224};
ram[23317] = {-9'd20,-10'd220};
ram[23318] = {-9'd17,-10'd217};
ram[23319] = {-9'd14,-10'd214};
ram[23320] = {-9'd11,-10'd211};
ram[23321] = {-9'd8,-10'd208};
ram[23322] = {-9'd4,-10'd205};
ram[23323] = {-9'd1,-10'd202};
ram[23324] = {9'd2,-10'd198};
ram[23325] = {9'd5,-10'd195};
ram[23326] = {9'd8,-10'd192};
ram[23327] = {9'd11,-10'd189};
ram[23328] = {9'd14,-10'd186};
ram[23329] = {9'd18,-10'd183};
ram[23330] = {9'd21,-10'd180};
ram[23331] = {9'd24,-10'd176};
ram[23332] = {9'd27,-10'd173};
ram[23333] = {9'd30,-10'd170};
ram[23334] = {9'd33,-10'd167};
ram[23335] = {9'd36,-10'd164};
ram[23336] = {9'd40,-10'd161};
ram[23337] = {9'd43,-10'd158};
ram[23338] = {9'd46,-10'd154};
ram[23339] = {9'd49,-10'd151};
ram[23340] = {9'd52,-10'd148};
ram[23341] = {9'd55,-10'd145};
ram[23342] = {9'd58,-10'd142};
ram[23343] = {9'd62,-10'd139};
ram[23344] = {9'd65,-10'd136};
ram[23345] = {9'd68,-10'd132};
ram[23346] = {9'd71,-10'd129};
ram[23347] = {9'd74,-10'd126};
ram[23348] = {9'd77,-10'd123};
ram[23349] = {9'd80,-10'd120};
ram[23350] = {9'd84,-10'd117};
ram[23351] = {9'd87,-10'd114};
ram[23352] = {9'd90,-10'd110};
ram[23353] = {9'd93,-10'd107};
ram[23354] = {9'd96,-10'd104};
ram[23355] = {9'd99,-10'd101};
ram[23356] = {-9'd98,-10'd98};
ram[23357] = {-9'd95,-10'd95};
ram[23358] = {-9'd92,-10'd92};
ram[23359] = {-9'd88,-10'd88};
ram[23360] = {-9'd85,-10'd85};
ram[23361] = {-9'd82,-10'd82};
ram[23362] = {-9'd79,-10'd79};
ram[23363] = {-9'd76,-10'd76};
ram[23364] = {-9'd73,-10'd73};
ram[23365] = {-9'd70,-10'd70};
ram[23366] = {-9'd66,-10'd66};
ram[23367] = {-9'd63,-10'd63};
ram[23368] = {-9'd60,-10'd60};
ram[23369] = {-9'd57,-10'd57};
ram[23370] = {-9'd54,-10'd54};
ram[23371] = {-9'd51,-10'd51};
ram[23372] = {-9'd48,-10'd48};
ram[23373] = {-9'd44,-10'd44};
ram[23374] = {-9'd41,-10'd41};
ram[23375] = {-9'd38,-10'd38};
ram[23376] = {-9'd35,-10'd35};
ram[23377] = {-9'd32,-10'd32};
ram[23378] = {-9'd29,-10'd29};
ram[23379] = {-9'd26,-10'd26};
ram[23380] = {-9'd22,-10'd22};
ram[23381] = {-9'd19,-10'd19};
ram[23382] = {-9'd16,-10'd16};
ram[23383] = {-9'd13,-10'd13};
ram[23384] = {-9'd10,-10'd10};
ram[23385] = {-9'd7,-10'd7};
ram[23386] = {-9'd4,-10'd4};
ram[23387] = {9'd0,10'd0};
ram[23388] = {9'd3,10'd3};
ram[23389] = {9'd6,10'd6};
ram[23390] = {9'd9,10'd9};
ram[23391] = {9'd12,10'd12};
ram[23392] = {9'd15,10'd15};
ram[23393] = {9'd18,10'd18};
ram[23394] = {9'd21,10'd21};
ram[23395] = {9'd25,10'd25};
ram[23396] = {9'd28,10'd28};
ram[23397] = {9'd31,10'd31};
ram[23398] = {9'd34,10'd34};
ram[23399] = {9'd37,10'd37};
ram[23400] = {9'd40,10'd40};
ram[23401] = {9'd43,10'd43};
ram[23402] = {9'd47,10'd47};
ram[23403] = {9'd50,10'd50};
ram[23404] = {9'd53,10'd53};
ram[23405] = {9'd56,10'd56};
ram[23406] = {9'd59,10'd59};
ram[23407] = {9'd62,10'd62};
ram[23408] = {9'd65,10'd65};
ram[23409] = {9'd69,10'd69};
ram[23410] = {9'd72,10'd72};
ram[23411] = {9'd75,10'd75};
ram[23412] = {9'd78,10'd78};
ram[23413] = {9'd81,10'd81};
ram[23414] = {9'd84,10'd84};
ram[23415] = {9'd87,10'd87};
ram[23416] = {9'd91,10'd91};
ram[23417] = {9'd94,10'd94};
ram[23418] = {9'd97,10'd97};
ram[23419] = {-9'd100,10'd100};
ram[23420] = {-9'd97,10'd103};
ram[23421] = {-9'd94,10'd106};
ram[23422] = {-9'd91,10'd109};
ram[23423] = {-9'd88,10'd113};
ram[23424] = {-9'd88,10'd113};
ram[23425] = {-9'd85,10'd116};
ram[23426] = {-9'd81,10'd119};
ram[23427] = {-9'd78,10'd122};
ram[23428] = {-9'd75,10'd125};
ram[23429] = {-9'd72,10'd128};
ram[23430] = {-9'd69,10'd131};
ram[23431] = {-9'd66,10'd135};
ram[23432] = {-9'd63,10'd138};
ram[23433] = {-9'd59,10'd141};
ram[23434] = {-9'd56,10'd144};
ram[23435] = {-9'd53,10'd147};
ram[23436] = {-9'd50,10'd150};
ram[23437] = {-9'd47,10'd153};
ram[23438] = {-9'd44,10'd157};
ram[23439] = {-9'd41,10'd160};
ram[23440] = {-9'd37,10'd163};
ram[23441] = {-9'd34,10'd166};
ram[23442] = {-9'd31,10'd169};
ram[23443] = {-9'd28,10'd172};
ram[23444] = {-9'd25,10'd175};
ram[23445] = {-9'd22,10'd179};
ram[23446] = {-9'd19,10'd182};
ram[23447] = {-9'd15,10'd185};
ram[23448] = {-9'd12,10'd188};
ram[23449] = {-9'd9,10'd191};
ram[23450] = {-9'd6,10'd194};
ram[23451] = {-9'd3,10'd197};
ram[23452] = {9'd0,10'd201};
ram[23453] = {9'd3,10'd204};
ram[23454] = {9'd7,10'd207};
ram[23455] = {9'd10,10'd210};
ram[23456] = {9'd13,10'd213};
ram[23457] = {9'd16,10'd216};
ram[23458] = {9'd19,10'd219};
ram[23459] = {9'd22,10'd223};
ram[23460] = {9'd25,10'd226};
ram[23461] = {9'd29,10'd229};
ram[23462] = {9'd32,10'd232};
ram[23463] = {9'd35,10'd235};
ram[23464] = {9'd38,10'd238};
ram[23465] = {9'd41,10'd241};
ram[23466] = {9'd44,10'd245};
ram[23467] = {9'd47,10'd248};
ram[23468] = {9'd51,10'd251};
ram[23469] = {9'd54,10'd254};
ram[23470] = {9'd57,10'd257};
ram[23471] = {9'd60,10'd260};
ram[23472] = {9'd63,10'd263};
ram[23473] = {9'd66,10'd267};
ram[23474] = {9'd69,10'd270};
ram[23475] = {9'd73,10'd273};
ram[23476] = {9'd76,10'd276};
ram[23477] = {9'd79,10'd279};
ram[23478] = {9'd82,10'd282};
ram[23479] = {9'd85,10'd285};
ram[23480] = {9'd88,10'd289};
ram[23481] = {9'd91,10'd292};
ram[23482] = {9'd95,10'd295};
ram[23483] = {9'd98,10'd298};
ram[23484] = {-9'd99,10'd301};
ram[23485] = {-9'd96,10'd304};
ram[23486] = {-9'd93,10'd307};
ram[23487] = {-9'd90,10'd311};
ram[23488] = {-9'd87,10'd314};
ram[23489] = {-9'd84,10'd317};
ram[23490] = {-9'd81,10'd320};
ram[23491] = {-9'd77,10'd323};
ram[23492] = {-9'd74,10'd326};
ram[23493] = {-9'd71,10'd329};
ram[23494] = {-9'd68,10'd333};
ram[23495] = {-9'd65,10'd336};
ram[23496] = {-9'd62,10'd339};
ram[23497] = {-9'd59,10'd342};
ram[23498] = {-9'd55,10'd345};
ram[23499] = {-9'd52,10'd348};
ram[23500] = {-9'd49,10'd351};
ram[23501] = {-9'd46,10'd354};
ram[23502] = {-9'd43,10'd358};
ram[23503] = {-9'd40,10'd361};
ram[23504] = {-9'd37,10'd364};
ram[23505] = {-9'd33,10'd367};
ram[23506] = {-9'd30,10'd370};
ram[23507] = {-9'd27,10'd373};
ram[23508] = {-9'd24,10'd376};
ram[23509] = {-9'd21,10'd380};
ram[23510] = {-9'd18,10'd383};
ram[23511] = {-9'd15,10'd386};
ram[23512] = {-9'd11,10'd389};
ram[23513] = {-9'd8,10'd392};
ram[23514] = {-9'd5,10'd395};
ram[23515] = {-9'd2,10'd398};
ram[23516] = {9'd1,-10'd399};
ram[23517] = {9'd4,-10'd396};
ram[23518] = {9'd7,-10'd393};
ram[23519] = {9'd10,-10'd390};
ram[23520] = {9'd14,-10'd387};
ram[23521] = {9'd17,-10'd384};
ram[23522] = {9'd20,-10'd381};
ram[23523] = {9'd23,-10'd377};
ram[23524] = {9'd26,-10'd374};
ram[23525] = {9'd29,-10'd371};
ram[23526] = {9'd32,-10'd368};
ram[23527] = {9'd36,-10'd365};
ram[23528] = {9'd39,-10'd362};
ram[23529] = {9'd42,-10'd359};
ram[23530] = {9'd45,-10'd355};
ram[23531] = {9'd48,-10'd352};
ram[23532] = {9'd51,-10'd349};
ram[23533] = {9'd54,-10'd346};
ram[23534] = {9'd58,-10'd343};
ram[23535] = {9'd61,-10'd340};
ram[23536] = {9'd64,-10'd337};
ram[23537] = {9'd67,-10'd334};
ram[23538] = {9'd70,-10'd330};
ram[23539] = {9'd73,-10'd327};
ram[23540] = {9'd76,-10'd324};
ram[23541] = {9'd80,-10'd321};
ram[23542] = {9'd83,-10'd318};
ram[23543] = {9'd86,-10'd315};
ram[23544] = {9'd89,-10'd312};
ram[23545] = {9'd92,-10'd308};
ram[23546] = {9'd95,-10'd305};
ram[23547] = {9'd98,-10'd302};
ram[23548] = {-9'd99,-10'd299};
ram[23549] = {-9'd96,-10'd296};
ram[23550] = {-9'd92,-10'd293};
ram[23551] = {-9'd89,-10'd290};
ram[23552] = {-9'd89,-10'd290};
ram[23553] = {-9'd86,-10'd286};
ram[23554] = {-9'd83,-10'd283};
ram[23555] = {-9'd80,-10'd280};
ram[23556] = {-9'd77,-10'd277};
ram[23557] = {-9'd74,-10'd274};
ram[23558] = {-9'd70,-10'd271};
ram[23559] = {-9'd67,-10'd268};
ram[23560] = {-9'd64,-10'd264};
ram[23561] = {-9'd61,-10'd261};
ram[23562] = {-9'd58,-10'd258};
ram[23563] = {-9'd55,-10'd255};
ram[23564] = {-9'd52,-10'd252};
ram[23565] = {-9'd48,-10'd249};
ram[23566] = {-9'd45,-10'd246};
ram[23567] = {-9'd42,-10'd242};
ram[23568] = {-9'd39,-10'd239};
ram[23569] = {-9'd36,-10'd236};
ram[23570] = {-9'd33,-10'd233};
ram[23571] = {-9'd30,-10'd230};
ram[23572] = {-9'd26,-10'd227};
ram[23573] = {-9'd23,-10'd224};
ram[23574] = {-9'd20,-10'd220};
ram[23575] = {-9'd17,-10'd217};
ram[23576] = {-9'd14,-10'd214};
ram[23577] = {-9'd11,-10'd211};
ram[23578] = {-9'd8,-10'd208};
ram[23579] = {-9'd4,-10'd205};
ram[23580] = {-9'd1,-10'd202};
ram[23581] = {9'd2,-10'd198};
ram[23582] = {9'd5,-10'd195};
ram[23583] = {9'd8,-10'd192};
ram[23584] = {9'd11,-10'd189};
ram[23585] = {9'd14,-10'd186};
ram[23586] = {9'd18,-10'd183};
ram[23587] = {9'd21,-10'd180};
ram[23588] = {9'd24,-10'd176};
ram[23589] = {9'd27,-10'd173};
ram[23590] = {9'd30,-10'd170};
ram[23591] = {9'd33,-10'd167};
ram[23592] = {9'd36,-10'd164};
ram[23593] = {9'd40,-10'd161};
ram[23594] = {9'd43,-10'd158};
ram[23595] = {9'd46,-10'd154};
ram[23596] = {9'd49,-10'd151};
ram[23597] = {9'd52,-10'd148};
ram[23598] = {9'd55,-10'd145};
ram[23599] = {9'd58,-10'd142};
ram[23600] = {9'd62,-10'd139};
ram[23601] = {9'd65,-10'd136};
ram[23602] = {9'd68,-10'd132};
ram[23603] = {9'd71,-10'd129};
ram[23604] = {9'd74,-10'd126};
ram[23605] = {9'd77,-10'd123};
ram[23606] = {9'd80,-10'd120};
ram[23607] = {9'd84,-10'd117};
ram[23608] = {9'd87,-10'd114};
ram[23609] = {9'd90,-10'd110};
ram[23610] = {9'd93,-10'd107};
ram[23611] = {9'd96,-10'd104};
ram[23612] = {9'd99,-10'd101};
ram[23613] = {-9'd98,-10'd98};
ram[23614] = {-9'd95,-10'd95};
ram[23615] = {-9'd92,-10'd92};
ram[23616] = {-9'd88,-10'd88};
ram[23617] = {-9'd85,-10'd85};
ram[23618] = {-9'd82,-10'd82};
ram[23619] = {-9'd79,-10'd79};
ram[23620] = {-9'd76,-10'd76};
ram[23621] = {-9'd73,-10'd73};
ram[23622] = {-9'd70,-10'd70};
ram[23623] = {-9'd66,-10'd66};
ram[23624] = {-9'd63,-10'd63};
ram[23625] = {-9'd60,-10'd60};
ram[23626] = {-9'd57,-10'd57};
ram[23627] = {-9'd54,-10'd54};
ram[23628] = {-9'd51,-10'd51};
ram[23629] = {-9'd48,-10'd48};
ram[23630] = {-9'd44,-10'd44};
ram[23631] = {-9'd41,-10'd41};
ram[23632] = {-9'd38,-10'd38};
ram[23633] = {-9'd35,-10'd35};
ram[23634] = {-9'd32,-10'd32};
ram[23635] = {-9'd29,-10'd29};
ram[23636] = {-9'd26,-10'd26};
ram[23637] = {-9'd22,-10'd22};
ram[23638] = {-9'd19,-10'd19};
ram[23639] = {-9'd16,-10'd16};
ram[23640] = {-9'd13,-10'd13};
ram[23641] = {-9'd10,-10'd10};
ram[23642] = {-9'd7,-10'd7};
ram[23643] = {-9'd4,-10'd4};
ram[23644] = {9'd0,10'd0};
ram[23645] = {9'd3,10'd3};
ram[23646] = {9'd6,10'd6};
ram[23647] = {9'd9,10'd9};
ram[23648] = {9'd12,10'd12};
ram[23649] = {9'd15,10'd15};
ram[23650] = {9'd18,10'd18};
ram[23651] = {9'd21,10'd21};
ram[23652] = {9'd25,10'd25};
ram[23653] = {9'd28,10'd28};
ram[23654] = {9'd31,10'd31};
ram[23655] = {9'd34,10'd34};
ram[23656] = {9'd37,10'd37};
ram[23657] = {9'd40,10'd40};
ram[23658] = {9'd43,10'd43};
ram[23659] = {9'd47,10'd47};
ram[23660] = {9'd50,10'd50};
ram[23661] = {9'd53,10'd53};
ram[23662] = {9'd56,10'd56};
ram[23663] = {9'd59,10'd59};
ram[23664] = {9'd62,10'd62};
ram[23665] = {9'd65,10'd65};
ram[23666] = {9'd69,10'd69};
ram[23667] = {9'd72,10'd72};
ram[23668] = {9'd75,10'd75};
ram[23669] = {9'd78,10'd78};
ram[23670] = {9'd81,10'd81};
ram[23671] = {9'd84,10'd84};
ram[23672] = {9'd87,10'd87};
ram[23673] = {9'd91,10'd91};
ram[23674] = {9'd94,10'd94};
ram[23675] = {9'd97,10'd97};
ram[23676] = {-9'd100,10'd100};
ram[23677] = {-9'd97,10'd103};
ram[23678] = {-9'd94,10'd106};
ram[23679] = {-9'd91,10'd109};
ram[23680] = {-9'd91,10'd109};
ram[23681] = {-9'd88,10'd113};
ram[23682] = {-9'd85,10'd116};
ram[23683] = {-9'd81,10'd119};
ram[23684] = {-9'd78,10'd122};
ram[23685] = {-9'd75,10'd125};
ram[23686] = {-9'd72,10'd128};
ram[23687] = {-9'd69,10'd131};
ram[23688] = {-9'd66,10'd135};
ram[23689] = {-9'd63,10'd138};
ram[23690] = {-9'd59,10'd141};
ram[23691] = {-9'd56,10'd144};
ram[23692] = {-9'd53,10'd147};
ram[23693] = {-9'd50,10'd150};
ram[23694] = {-9'd47,10'd153};
ram[23695] = {-9'd44,10'd157};
ram[23696] = {-9'd41,10'd160};
ram[23697] = {-9'd37,10'd163};
ram[23698] = {-9'd34,10'd166};
ram[23699] = {-9'd31,10'd169};
ram[23700] = {-9'd28,10'd172};
ram[23701] = {-9'd25,10'd175};
ram[23702] = {-9'd22,10'd179};
ram[23703] = {-9'd19,10'd182};
ram[23704] = {-9'd15,10'd185};
ram[23705] = {-9'd12,10'd188};
ram[23706] = {-9'd9,10'd191};
ram[23707] = {-9'd6,10'd194};
ram[23708] = {-9'd3,10'd197};
ram[23709] = {9'd0,10'd201};
ram[23710] = {9'd3,10'd204};
ram[23711] = {9'd7,10'd207};
ram[23712] = {9'd10,10'd210};
ram[23713] = {9'd13,10'd213};
ram[23714] = {9'd16,10'd216};
ram[23715] = {9'd19,10'd219};
ram[23716] = {9'd22,10'd223};
ram[23717] = {9'd25,10'd226};
ram[23718] = {9'd29,10'd229};
ram[23719] = {9'd32,10'd232};
ram[23720] = {9'd35,10'd235};
ram[23721] = {9'd38,10'd238};
ram[23722] = {9'd41,10'd241};
ram[23723] = {9'd44,10'd245};
ram[23724] = {9'd47,10'd248};
ram[23725] = {9'd51,10'd251};
ram[23726] = {9'd54,10'd254};
ram[23727] = {9'd57,10'd257};
ram[23728] = {9'd60,10'd260};
ram[23729] = {9'd63,10'd263};
ram[23730] = {9'd66,10'd267};
ram[23731] = {9'd69,10'd270};
ram[23732] = {9'd73,10'd273};
ram[23733] = {9'd76,10'd276};
ram[23734] = {9'd79,10'd279};
ram[23735] = {9'd82,10'd282};
ram[23736] = {9'd85,10'd285};
ram[23737] = {9'd88,10'd289};
ram[23738] = {9'd91,10'd292};
ram[23739] = {9'd95,10'd295};
ram[23740] = {9'd98,10'd298};
ram[23741] = {-9'd99,10'd301};
ram[23742] = {-9'd96,10'd304};
ram[23743] = {-9'd93,10'd307};
ram[23744] = {-9'd90,10'd311};
ram[23745] = {-9'd87,10'd314};
ram[23746] = {-9'd84,10'd317};
ram[23747] = {-9'd81,10'd320};
ram[23748] = {-9'd77,10'd323};
ram[23749] = {-9'd74,10'd326};
ram[23750] = {-9'd71,10'd329};
ram[23751] = {-9'd68,10'd333};
ram[23752] = {-9'd65,10'd336};
ram[23753] = {-9'd62,10'd339};
ram[23754] = {-9'd59,10'd342};
ram[23755] = {-9'd55,10'd345};
ram[23756] = {-9'd52,10'd348};
ram[23757] = {-9'd49,10'd351};
ram[23758] = {-9'd46,10'd354};
ram[23759] = {-9'd43,10'd358};
ram[23760] = {-9'd40,10'd361};
ram[23761] = {-9'd37,10'd364};
ram[23762] = {-9'd33,10'd367};
ram[23763] = {-9'd30,10'd370};
ram[23764] = {-9'd27,10'd373};
ram[23765] = {-9'd24,10'd376};
ram[23766] = {-9'd21,10'd380};
ram[23767] = {-9'd18,10'd383};
ram[23768] = {-9'd15,10'd386};
ram[23769] = {-9'd11,10'd389};
ram[23770] = {-9'd8,10'd392};
ram[23771] = {-9'd5,10'd395};
ram[23772] = {-9'd2,10'd398};
ram[23773] = {9'd1,-10'd399};
ram[23774] = {9'd4,-10'd396};
ram[23775] = {9'd7,-10'd393};
ram[23776] = {9'd10,-10'd390};
ram[23777] = {9'd14,-10'd387};
ram[23778] = {9'd17,-10'd384};
ram[23779] = {9'd20,-10'd381};
ram[23780] = {9'd23,-10'd377};
ram[23781] = {9'd26,-10'd374};
ram[23782] = {9'd29,-10'd371};
ram[23783] = {9'd32,-10'd368};
ram[23784] = {9'd36,-10'd365};
ram[23785] = {9'd39,-10'd362};
ram[23786] = {9'd42,-10'd359};
ram[23787] = {9'd45,-10'd355};
ram[23788] = {9'd48,-10'd352};
ram[23789] = {9'd51,-10'd349};
ram[23790] = {9'd54,-10'd346};
ram[23791] = {9'd58,-10'd343};
ram[23792] = {9'd61,-10'd340};
ram[23793] = {9'd64,-10'd337};
ram[23794] = {9'd67,-10'd334};
ram[23795] = {9'd70,-10'd330};
ram[23796] = {9'd73,-10'd327};
ram[23797] = {9'd76,-10'd324};
ram[23798] = {9'd80,-10'd321};
ram[23799] = {9'd83,-10'd318};
ram[23800] = {9'd86,-10'd315};
ram[23801] = {9'd89,-10'd312};
ram[23802] = {9'd92,-10'd308};
ram[23803] = {9'd95,-10'd305};
ram[23804] = {9'd98,-10'd302};
ram[23805] = {-9'd99,-10'd299};
ram[23806] = {-9'd96,-10'd296};
ram[23807] = {-9'd92,-10'd293};
ram[23808] = {-9'd92,-10'd293};
ram[23809] = {-9'd89,-10'd290};
ram[23810] = {-9'd86,-10'd286};
ram[23811] = {-9'd83,-10'd283};
ram[23812] = {-9'd80,-10'd280};
ram[23813] = {-9'd77,-10'd277};
ram[23814] = {-9'd74,-10'd274};
ram[23815] = {-9'd70,-10'd271};
ram[23816] = {-9'd67,-10'd268};
ram[23817] = {-9'd64,-10'd264};
ram[23818] = {-9'd61,-10'd261};
ram[23819] = {-9'd58,-10'd258};
ram[23820] = {-9'd55,-10'd255};
ram[23821] = {-9'd52,-10'd252};
ram[23822] = {-9'd48,-10'd249};
ram[23823] = {-9'd45,-10'd246};
ram[23824] = {-9'd42,-10'd242};
ram[23825] = {-9'd39,-10'd239};
ram[23826] = {-9'd36,-10'd236};
ram[23827] = {-9'd33,-10'd233};
ram[23828] = {-9'd30,-10'd230};
ram[23829] = {-9'd26,-10'd227};
ram[23830] = {-9'd23,-10'd224};
ram[23831] = {-9'd20,-10'd220};
ram[23832] = {-9'd17,-10'd217};
ram[23833] = {-9'd14,-10'd214};
ram[23834] = {-9'd11,-10'd211};
ram[23835] = {-9'd8,-10'd208};
ram[23836] = {-9'd4,-10'd205};
ram[23837] = {-9'd1,-10'd202};
ram[23838] = {9'd2,-10'd198};
ram[23839] = {9'd5,-10'd195};
ram[23840] = {9'd8,-10'd192};
ram[23841] = {9'd11,-10'd189};
ram[23842] = {9'd14,-10'd186};
ram[23843] = {9'd18,-10'd183};
ram[23844] = {9'd21,-10'd180};
ram[23845] = {9'd24,-10'd176};
ram[23846] = {9'd27,-10'd173};
ram[23847] = {9'd30,-10'd170};
ram[23848] = {9'd33,-10'd167};
ram[23849] = {9'd36,-10'd164};
ram[23850] = {9'd40,-10'd161};
ram[23851] = {9'd43,-10'd158};
ram[23852] = {9'd46,-10'd154};
ram[23853] = {9'd49,-10'd151};
ram[23854] = {9'd52,-10'd148};
ram[23855] = {9'd55,-10'd145};
ram[23856] = {9'd58,-10'd142};
ram[23857] = {9'd62,-10'd139};
ram[23858] = {9'd65,-10'd136};
ram[23859] = {9'd68,-10'd132};
ram[23860] = {9'd71,-10'd129};
ram[23861] = {9'd74,-10'd126};
ram[23862] = {9'd77,-10'd123};
ram[23863] = {9'd80,-10'd120};
ram[23864] = {9'd84,-10'd117};
ram[23865] = {9'd87,-10'd114};
ram[23866] = {9'd90,-10'd110};
ram[23867] = {9'd93,-10'd107};
ram[23868] = {9'd96,-10'd104};
ram[23869] = {9'd99,-10'd101};
ram[23870] = {-9'd98,-10'd98};
ram[23871] = {-9'd95,-10'd95};
ram[23872] = {-9'd92,-10'd92};
ram[23873] = {-9'd88,-10'd88};
ram[23874] = {-9'd85,-10'd85};
ram[23875] = {-9'd82,-10'd82};
ram[23876] = {-9'd79,-10'd79};
ram[23877] = {-9'd76,-10'd76};
ram[23878] = {-9'd73,-10'd73};
ram[23879] = {-9'd70,-10'd70};
ram[23880] = {-9'd66,-10'd66};
ram[23881] = {-9'd63,-10'd63};
ram[23882] = {-9'd60,-10'd60};
ram[23883] = {-9'd57,-10'd57};
ram[23884] = {-9'd54,-10'd54};
ram[23885] = {-9'd51,-10'd51};
ram[23886] = {-9'd48,-10'd48};
ram[23887] = {-9'd44,-10'd44};
ram[23888] = {-9'd41,-10'd41};
ram[23889] = {-9'd38,-10'd38};
ram[23890] = {-9'd35,-10'd35};
ram[23891] = {-9'd32,-10'd32};
ram[23892] = {-9'd29,-10'd29};
ram[23893] = {-9'd26,-10'd26};
ram[23894] = {-9'd22,-10'd22};
ram[23895] = {-9'd19,-10'd19};
ram[23896] = {-9'd16,-10'd16};
ram[23897] = {-9'd13,-10'd13};
ram[23898] = {-9'd10,-10'd10};
ram[23899] = {-9'd7,-10'd7};
ram[23900] = {-9'd4,-10'd4};
ram[23901] = {9'd0,10'd0};
ram[23902] = {9'd3,10'd3};
ram[23903] = {9'd6,10'd6};
ram[23904] = {9'd9,10'd9};
ram[23905] = {9'd12,10'd12};
ram[23906] = {9'd15,10'd15};
ram[23907] = {9'd18,10'd18};
ram[23908] = {9'd21,10'd21};
ram[23909] = {9'd25,10'd25};
ram[23910] = {9'd28,10'd28};
ram[23911] = {9'd31,10'd31};
ram[23912] = {9'd34,10'd34};
ram[23913] = {9'd37,10'd37};
ram[23914] = {9'd40,10'd40};
ram[23915] = {9'd43,10'd43};
ram[23916] = {9'd47,10'd47};
ram[23917] = {9'd50,10'd50};
ram[23918] = {9'd53,10'd53};
ram[23919] = {9'd56,10'd56};
ram[23920] = {9'd59,10'd59};
ram[23921] = {9'd62,10'd62};
ram[23922] = {9'd65,10'd65};
ram[23923] = {9'd69,10'd69};
ram[23924] = {9'd72,10'd72};
ram[23925] = {9'd75,10'd75};
ram[23926] = {9'd78,10'd78};
ram[23927] = {9'd81,10'd81};
ram[23928] = {9'd84,10'd84};
ram[23929] = {9'd87,10'd87};
ram[23930] = {9'd91,10'd91};
ram[23931] = {9'd94,10'd94};
ram[23932] = {9'd97,10'd97};
ram[23933] = {-9'd100,10'd100};
ram[23934] = {-9'd97,10'd103};
ram[23935] = {-9'd94,10'd106};
ram[23936] = {-9'd94,10'd106};
ram[23937] = {-9'd91,10'd109};
ram[23938] = {-9'd88,10'd113};
ram[23939] = {-9'd85,10'd116};
ram[23940] = {-9'd81,10'd119};
ram[23941] = {-9'd78,10'd122};
ram[23942] = {-9'd75,10'd125};
ram[23943] = {-9'd72,10'd128};
ram[23944] = {-9'd69,10'd131};
ram[23945] = {-9'd66,10'd135};
ram[23946] = {-9'd63,10'd138};
ram[23947] = {-9'd59,10'd141};
ram[23948] = {-9'd56,10'd144};
ram[23949] = {-9'd53,10'd147};
ram[23950] = {-9'd50,10'd150};
ram[23951] = {-9'd47,10'd153};
ram[23952] = {-9'd44,10'd157};
ram[23953] = {-9'd41,10'd160};
ram[23954] = {-9'd37,10'd163};
ram[23955] = {-9'd34,10'd166};
ram[23956] = {-9'd31,10'd169};
ram[23957] = {-9'd28,10'd172};
ram[23958] = {-9'd25,10'd175};
ram[23959] = {-9'd22,10'd179};
ram[23960] = {-9'd19,10'd182};
ram[23961] = {-9'd15,10'd185};
ram[23962] = {-9'd12,10'd188};
ram[23963] = {-9'd9,10'd191};
ram[23964] = {-9'd6,10'd194};
ram[23965] = {-9'd3,10'd197};
ram[23966] = {9'd0,10'd201};
ram[23967] = {9'd3,10'd204};
ram[23968] = {9'd7,10'd207};
ram[23969] = {9'd10,10'd210};
ram[23970] = {9'd13,10'd213};
ram[23971] = {9'd16,10'd216};
ram[23972] = {9'd19,10'd219};
ram[23973] = {9'd22,10'd223};
ram[23974] = {9'd25,10'd226};
ram[23975] = {9'd29,10'd229};
ram[23976] = {9'd32,10'd232};
ram[23977] = {9'd35,10'd235};
ram[23978] = {9'd38,10'd238};
ram[23979] = {9'd41,10'd241};
ram[23980] = {9'd44,10'd245};
ram[23981] = {9'd47,10'd248};
ram[23982] = {9'd51,10'd251};
ram[23983] = {9'd54,10'd254};
ram[23984] = {9'd57,10'd257};
ram[23985] = {9'd60,10'd260};
ram[23986] = {9'd63,10'd263};
ram[23987] = {9'd66,10'd267};
ram[23988] = {9'd69,10'd270};
ram[23989] = {9'd73,10'd273};
ram[23990] = {9'd76,10'd276};
ram[23991] = {9'd79,10'd279};
ram[23992] = {9'd82,10'd282};
ram[23993] = {9'd85,10'd285};
ram[23994] = {9'd88,10'd289};
ram[23995] = {9'd91,10'd292};
ram[23996] = {9'd95,10'd295};
ram[23997] = {9'd98,10'd298};
ram[23998] = {-9'd99,10'd301};
ram[23999] = {-9'd96,10'd304};
ram[24000] = {-9'd93,10'd307};
ram[24001] = {-9'd90,10'd311};
ram[24002] = {-9'd87,10'd314};
ram[24003] = {-9'd84,10'd317};
ram[24004] = {-9'd81,10'd320};
ram[24005] = {-9'd77,10'd323};
ram[24006] = {-9'd74,10'd326};
ram[24007] = {-9'd71,10'd329};
ram[24008] = {-9'd68,10'd333};
ram[24009] = {-9'd65,10'd336};
ram[24010] = {-9'd62,10'd339};
ram[24011] = {-9'd59,10'd342};
ram[24012] = {-9'd55,10'd345};
ram[24013] = {-9'd52,10'd348};
ram[24014] = {-9'd49,10'd351};
ram[24015] = {-9'd46,10'd354};
ram[24016] = {-9'd43,10'd358};
ram[24017] = {-9'd40,10'd361};
ram[24018] = {-9'd37,10'd364};
ram[24019] = {-9'd33,10'd367};
ram[24020] = {-9'd30,10'd370};
ram[24021] = {-9'd27,10'd373};
ram[24022] = {-9'd24,10'd376};
ram[24023] = {-9'd21,10'd380};
ram[24024] = {-9'd18,10'd383};
ram[24025] = {-9'd15,10'd386};
ram[24026] = {-9'd11,10'd389};
ram[24027] = {-9'd8,10'd392};
ram[24028] = {-9'd5,10'd395};
ram[24029] = {-9'd2,10'd398};
ram[24030] = {9'd1,-10'd399};
ram[24031] = {9'd4,-10'd396};
ram[24032] = {9'd7,-10'd393};
ram[24033] = {9'd10,-10'd390};
ram[24034] = {9'd14,-10'd387};
ram[24035] = {9'd17,-10'd384};
ram[24036] = {9'd20,-10'd381};
ram[24037] = {9'd23,-10'd377};
ram[24038] = {9'd26,-10'd374};
ram[24039] = {9'd29,-10'd371};
ram[24040] = {9'd32,-10'd368};
ram[24041] = {9'd36,-10'd365};
ram[24042] = {9'd39,-10'd362};
ram[24043] = {9'd42,-10'd359};
ram[24044] = {9'd45,-10'd355};
ram[24045] = {9'd48,-10'd352};
ram[24046] = {9'd51,-10'd349};
ram[24047] = {9'd54,-10'd346};
ram[24048] = {9'd58,-10'd343};
ram[24049] = {9'd61,-10'd340};
ram[24050] = {9'd64,-10'd337};
ram[24051] = {9'd67,-10'd334};
ram[24052] = {9'd70,-10'd330};
ram[24053] = {9'd73,-10'd327};
ram[24054] = {9'd76,-10'd324};
ram[24055] = {9'd80,-10'd321};
ram[24056] = {9'd83,-10'd318};
ram[24057] = {9'd86,-10'd315};
ram[24058] = {9'd89,-10'd312};
ram[24059] = {9'd92,-10'd308};
ram[24060] = {9'd95,-10'd305};
ram[24061] = {9'd98,-10'd302};
ram[24062] = {-9'd99,-10'd299};
ram[24063] = {-9'd96,-10'd296};
ram[24064] = {-9'd96,-10'd296};
ram[24065] = {-9'd92,-10'd293};
ram[24066] = {-9'd89,-10'd290};
ram[24067] = {-9'd86,-10'd286};
ram[24068] = {-9'd83,-10'd283};
ram[24069] = {-9'd80,-10'd280};
ram[24070] = {-9'd77,-10'd277};
ram[24071] = {-9'd74,-10'd274};
ram[24072] = {-9'd70,-10'd271};
ram[24073] = {-9'd67,-10'd268};
ram[24074] = {-9'd64,-10'd264};
ram[24075] = {-9'd61,-10'd261};
ram[24076] = {-9'd58,-10'd258};
ram[24077] = {-9'd55,-10'd255};
ram[24078] = {-9'd52,-10'd252};
ram[24079] = {-9'd48,-10'd249};
ram[24080] = {-9'd45,-10'd246};
ram[24081] = {-9'd42,-10'd242};
ram[24082] = {-9'd39,-10'd239};
ram[24083] = {-9'd36,-10'd236};
ram[24084] = {-9'd33,-10'd233};
ram[24085] = {-9'd30,-10'd230};
ram[24086] = {-9'd26,-10'd227};
ram[24087] = {-9'd23,-10'd224};
ram[24088] = {-9'd20,-10'd220};
ram[24089] = {-9'd17,-10'd217};
ram[24090] = {-9'd14,-10'd214};
ram[24091] = {-9'd11,-10'd211};
ram[24092] = {-9'd8,-10'd208};
ram[24093] = {-9'd4,-10'd205};
ram[24094] = {-9'd1,-10'd202};
ram[24095] = {9'd2,-10'd198};
ram[24096] = {9'd5,-10'd195};
ram[24097] = {9'd8,-10'd192};
ram[24098] = {9'd11,-10'd189};
ram[24099] = {9'd14,-10'd186};
ram[24100] = {9'd18,-10'd183};
ram[24101] = {9'd21,-10'd180};
ram[24102] = {9'd24,-10'd176};
ram[24103] = {9'd27,-10'd173};
ram[24104] = {9'd30,-10'd170};
ram[24105] = {9'd33,-10'd167};
ram[24106] = {9'd36,-10'd164};
ram[24107] = {9'd40,-10'd161};
ram[24108] = {9'd43,-10'd158};
ram[24109] = {9'd46,-10'd154};
ram[24110] = {9'd49,-10'd151};
ram[24111] = {9'd52,-10'd148};
ram[24112] = {9'd55,-10'd145};
ram[24113] = {9'd58,-10'd142};
ram[24114] = {9'd62,-10'd139};
ram[24115] = {9'd65,-10'd136};
ram[24116] = {9'd68,-10'd132};
ram[24117] = {9'd71,-10'd129};
ram[24118] = {9'd74,-10'd126};
ram[24119] = {9'd77,-10'd123};
ram[24120] = {9'd80,-10'd120};
ram[24121] = {9'd84,-10'd117};
ram[24122] = {9'd87,-10'd114};
ram[24123] = {9'd90,-10'd110};
ram[24124] = {9'd93,-10'd107};
ram[24125] = {9'd96,-10'd104};
ram[24126] = {9'd99,-10'd101};
ram[24127] = {-9'd98,-10'd98};
ram[24128] = {-9'd95,-10'd95};
ram[24129] = {-9'd92,-10'd92};
ram[24130] = {-9'd88,-10'd88};
ram[24131] = {-9'd85,-10'd85};
ram[24132] = {-9'd82,-10'd82};
ram[24133] = {-9'd79,-10'd79};
ram[24134] = {-9'd76,-10'd76};
ram[24135] = {-9'd73,-10'd73};
ram[24136] = {-9'd70,-10'd70};
ram[24137] = {-9'd66,-10'd66};
ram[24138] = {-9'd63,-10'd63};
ram[24139] = {-9'd60,-10'd60};
ram[24140] = {-9'd57,-10'd57};
ram[24141] = {-9'd54,-10'd54};
ram[24142] = {-9'd51,-10'd51};
ram[24143] = {-9'd48,-10'd48};
ram[24144] = {-9'd44,-10'd44};
ram[24145] = {-9'd41,-10'd41};
ram[24146] = {-9'd38,-10'd38};
ram[24147] = {-9'd35,-10'd35};
ram[24148] = {-9'd32,-10'd32};
ram[24149] = {-9'd29,-10'd29};
ram[24150] = {-9'd26,-10'd26};
ram[24151] = {-9'd22,-10'd22};
ram[24152] = {-9'd19,-10'd19};
ram[24153] = {-9'd16,-10'd16};
ram[24154] = {-9'd13,-10'd13};
ram[24155] = {-9'd10,-10'd10};
ram[24156] = {-9'd7,-10'd7};
ram[24157] = {-9'd4,-10'd4};
ram[24158] = {9'd0,10'd0};
ram[24159] = {9'd3,10'd3};
ram[24160] = {9'd6,10'd6};
ram[24161] = {9'd9,10'd9};
ram[24162] = {9'd12,10'd12};
ram[24163] = {9'd15,10'd15};
ram[24164] = {9'd18,10'd18};
ram[24165] = {9'd21,10'd21};
ram[24166] = {9'd25,10'd25};
ram[24167] = {9'd28,10'd28};
ram[24168] = {9'd31,10'd31};
ram[24169] = {9'd34,10'd34};
ram[24170] = {9'd37,10'd37};
ram[24171] = {9'd40,10'd40};
ram[24172] = {9'd43,10'd43};
ram[24173] = {9'd47,10'd47};
ram[24174] = {9'd50,10'd50};
ram[24175] = {9'd53,10'd53};
ram[24176] = {9'd56,10'd56};
ram[24177] = {9'd59,10'd59};
ram[24178] = {9'd62,10'd62};
ram[24179] = {9'd65,10'd65};
ram[24180] = {9'd69,10'd69};
ram[24181] = {9'd72,10'd72};
ram[24182] = {9'd75,10'd75};
ram[24183] = {9'd78,10'd78};
ram[24184] = {9'd81,10'd81};
ram[24185] = {9'd84,10'd84};
ram[24186] = {9'd87,10'd87};
ram[24187] = {9'd91,10'd91};
ram[24188] = {9'd94,10'd94};
ram[24189] = {9'd97,10'd97};
ram[24190] = {-9'd100,10'd100};
ram[24191] = {-9'd97,10'd103};
ram[24192] = {-9'd97,10'd103};
ram[24193] = {-9'd94,10'd106};
ram[24194] = {-9'd91,10'd109};
ram[24195] = {-9'd88,10'd113};
ram[24196] = {-9'd85,10'd116};
ram[24197] = {-9'd81,10'd119};
ram[24198] = {-9'd78,10'd122};
ram[24199] = {-9'd75,10'd125};
ram[24200] = {-9'd72,10'd128};
ram[24201] = {-9'd69,10'd131};
ram[24202] = {-9'd66,10'd135};
ram[24203] = {-9'd63,10'd138};
ram[24204] = {-9'd59,10'd141};
ram[24205] = {-9'd56,10'd144};
ram[24206] = {-9'd53,10'd147};
ram[24207] = {-9'd50,10'd150};
ram[24208] = {-9'd47,10'd153};
ram[24209] = {-9'd44,10'd157};
ram[24210] = {-9'd41,10'd160};
ram[24211] = {-9'd37,10'd163};
ram[24212] = {-9'd34,10'd166};
ram[24213] = {-9'd31,10'd169};
ram[24214] = {-9'd28,10'd172};
ram[24215] = {-9'd25,10'd175};
ram[24216] = {-9'd22,10'd179};
ram[24217] = {-9'd19,10'd182};
ram[24218] = {-9'd15,10'd185};
ram[24219] = {-9'd12,10'd188};
ram[24220] = {-9'd9,10'd191};
ram[24221] = {-9'd6,10'd194};
ram[24222] = {-9'd3,10'd197};
ram[24223] = {9'd0,10'd201};
ram[24224] = {9'd3,10'd204};
ram[24225] = {9'd7,10'd207};
ram[24226] = {9'd10,10'd210};
ram[24227] = {9'd13,10'd213};
ram[24228] = {9'd16,10'd216};
ram[24229] = {9'd19,10'd219};
ram[24230] = {9'd22,10'd223};
ram[24231] = {9'd25,10'd226};
ram[24232] = {9'd29,10'd229};
ram[24233] = {9'd32,10'd232};
ram[24234] = {9'd35,10'd235};
ram[24235] = {9'd38,10'd238};
ram[24236] = {9'd41,10'd241};
ram[24237] = {9'd44,10'd245};
ram[24238] = {9'd47,10'd248};
ram[24239] = {9'd51,10'd251};
ram[24240] = {9'd54,10'd254};
ram[24241] = {9'd57,10'd257};
ram[24242] = {9'd60,10'd260};
ram[24243] = {9'd63,10'd263};
ram[24244] = {9'd66,10'd267};
ram[24245] = {9'd69,10'd270};
ram[24246] = {9'd73,10'd273};
ram[24247] = {9'd76,10'd276};
ram[24248] = {9'd79,10'd279};
ram[24249] = {9'd82,10'd282};
ram[24250] = {9'd85,10'd285};
ram[24251] = {9'd88,10'd289};
ram[24252] = {9'd91,10'd292};
ram[24253] = {9'd95,10'd295};
ram[24254] = {9'd98,10'd298};
ram[24255] = {-9'd99,10'd301};
ram[24256] = {-9'd96,10'd304};
ram[24257] = {-9'd93,10'd307};
ram[24258] = {-9'd90,10'd311};
ram[24259] = {-9'd87,10'd314};
ram[24260] = {-9'd84,10'd317};
ram[24261] = {-9'd81,10'd320};
ram[24262] = {-9'd77,10'd323};
ram[24263] = {-9'd74,10'd326};
ram[24264] = {-9'd71,10'd329};
ram[24265] = {-9'd68,10'd333};
ram[24266] = {-9'd65,10'd336};
ram[24267] = {-9'd62,10'd339};
ram[24268] = {-9'd59,10'd342};
ram[24269] = {-9'd55,10'd345};
ram[24270] = {-9'd52,10'd348};
ram[24271] = {-9'd49,10'd351};
ram[24272] = {-9'd46,10'd354};
ram[24273] = {-9'd43,10'd358};
ram[24274] = {-9'd40,10'd361};
ram[24275] = {-9'd37,10'd364};
ram[24276] = {-9'd33,10'd367};
ram[24277] = {-9'd30,10'd370};
ram[24278] = {-9'd27,10'd373};
ram[24279] = {-9'd24,10'd376};
ram[24280] = {-9'd21,10'd380};
ram[24281] = {-9'd18,10'd383};
ram[24282] = {-9'd15,10'd386};
ram[24283] = {-9'd11,10'd389};
ram[24284] = {-9'd8,10'd392};
ram[24285] = {-9'd5,10'd395};
ram[24286] = {-9'd2,10'd398};
ram[24287] = {9'd1,-10'd399};
ram[24288] = {9'd4,-10'd396};
ram[24289] = {9'd7,-10'd393};
ram[24290] = {9'd10,-10'd390};
ram[24291] = {9'd14,-10'd387};
ram[24292] = {9'd17,-10'd384};
ram[24293] = {9'd20,-10'd381};
ram[24294] = {9'd23,-10'd377};
ram[24295] = {9'd26,-10'd374};
ram[24296] = {9'd29,-10'd371};
ram[24297] = {9'd32,-10'd368};
ram[24298] = {9'd36,-10'd365};
ram[24299] = {9'd39,-10'd362};
ram[24300] = {9'd42,-10'd359};
ram[24301] = {9'd45,-10'd355};
ram[24302] = {9'd48,-10'd352};
ram[24303] = {9'd51,-10'd349};
ram[24304] = {9'd54,-10'd346};
ram[24305] = {9'd58,-10'd343};
ram[24306] = {9'd61,-10'd340};
ram[24307] = {9'd64,-10'd337};
ram[24308] = {9'd67,-10'd334};
ram[24309] = {9'd70,-10'd330};
ram[24310] = {9'd73,-10'd327};
ram[24311] = {9'd76,-10'd324};
ram[24312] = {9'd80,-10'd321};
ram[24313] = {9'd83,-10'd318};
ram[24314] = {9'd86,-10'd315};
ram[24315] = {9'd89,-10'd312};
ram[24316] = {9'd92,-10'd308};
ram[24317] = {9'd95,-10'd305};
ram[24318] = {9'd98,-10'd302};
ram[24319] = {-9'd99,-10'd299};
ram[24320] = {-9'd99,-10'd299};
ram[24321] = {-9'd96,-10'd296};
ram[24322] = {-9'd92,-10'd293};
ram[24323] = {-9'd89,-10'd290};
ram[24324] = {-9'd86,-10'd286};
ram[24325] = {-9'd83,-10'd283};
ram[24326] = {-9'd80,-10'd280};
ram[24327] = {-9'd77,-10'd277};
ram[24328] = {-9'd74,-10'd274};
ram[24329] = {-9'd70,-10'd271};
ram[24330] = {-9'd67,-10'd268};
ram[24331] = {-9'd64,-10'd264};
ram[24332] = {-9'd61,-10'd261};
ram[24333] = {-9'd58,-10'd258};
ram[24334] = {-9'd55,-10'd255};
ram[24335] = {-9'd52,-10'd252};
ram[24336] = {-9'd48,-10'd249};
ram[24337] = {-9'd45,-10'd246};
ram[24338] = {-9'd42,-10'd242};
ram[24339] = {-9'd39,-10'd239};
ram[24340] = {-9'd36,-10'd236};
ram[24341] = {-9'd33,-10'd233};
ram[24342] = {-9'd30,-10'd230};
ram[24343] = {-9'd26,-10'd227};
ram[24344] = {-9'd23,-10'd224};
ram[24345] = {-9'd20,-10'd220};
ram[24346] = {-9'd17,-10'd217};
ram[24347] = {-9'd14,-10'd214};
ram[24348] = {-9'd11,-10'd211};
ram[24349] = {-9'd8,-10'd208};
ram[24350] = {-9'd4,-10'd205};
ram[24351] = {-9'd1,-10'd202};
ram[24352] = {9'd2,-10'd198};
ram[24353] = {9'd5,-10'd195};
ram[24354] = {9'd8,-10'd192};
ram[24355] = {9'd11,-10'd189};
ram[24356] = {9'd14,-10'd186};
ram[24357] = {9'd18,-10'd183};
ram[24358] = {9'd21,-10'd180};
ram[24359] = {9'd24,-10'd176};
ram[24360] = {9'd27,-10'd173};
ram[24361] = {9'd30,-10'd170};
ram[24362] = {9'd33,-10'd167};
ram[24363] = {9'd36,-10'd164};
ram[24364] = {9'd40,-10'd161};
ram[24365] = {9'd43,-10'd158};
ram[24366] = {9'd46,-10'd154};
ram[24367] = {9'd49,-10'd151};
ram[24368] = {9'd52,-10'd148};
ram[24369] = {9'd55,-10'd145};
ram[24370] = {9'd58,-10'd142};
ram[24371] = {9'd62,-10'd139};
ram[24372] = {9'd65,-10'd136};
ram[24373] = {9'd68,-10'd132};
ram[24374] = {9'd71,-10'd129};
ram[24375] = {9'd74,-10'd126};
ram[24376] = {9'd77,-10'd123};
ram[24377] = {9'd80,-10'd120};
ram[24378] = {9'd84,-10'd117};
ram[24379] = {9'd87,-10'd114};
ram[24380] = {9'd90,-10'd110};
ram[24381] = {9'd93,-10'd107};
ram[24382] = {9'd96,-10'd104};
ram[24383] = {9'd99,-10'd101};
ram[24384] = {-9'd98,-10'd98};
ram[24385] = {-9'd95,-10'd95};
ram[24386] = {-9'd92,-10'd92};
ram[24387] = {-9'd88,-10'd88};
ram[24388] = {-9'd85,-10'd85};
ram[24389] = {-9'd82,-10'd82};
ram[24390] = {-9'd79,-10'd79};
ram[24391] = {-9'd76,-10'd76};
ram[24392] = {-9'd73,-10'd73};
ram[24393] = {-9'd70,-10'd70};
ram[24394] = {-9'd66,-10'd66};
ram[24395] = {-9'd63,-10'd63};
ram[24396] = {-9'd60,-10'd60};
ram[24397] = {-9'd57,-10'd57};
ram[24398] = {-9'd54,-10'd54};
ram[24399] = {-9'd51,-10'd51};
ram[24400] = {-9'd48,-10'd48};
ram[24401] = {-9'd44,-10'd44};
ram[24402] = {-9'd41,-10'd41};
ram[24403] = {-9'd38,-10'd38};
ram[24404] = {-9'd35,-10'd35};
ram[24405] = {-9'd32,-10'd32};
ram[24406] = {-9'd29,-10'd29};
ram[24407] = {-9'd26,-10'd26};
ram[24408] = {-9'd22,-10'd22};
ram[24409] = {-9'd19,-10'd19};
ram[24410] = {-9'd16,-10'd16};
ram[24411] = {-9'd13,-10'd13};
ram[24412] = {-9'd10,-10'd10};
ram[24413] = {-9'd7,-10'd7};
ram[24414] = {-9'd4,-10'd4};
ram[24415] = {9'd0,10'd0};
ram[24416] = {9'd3,10'd3};
ram[24417] = {9'd6,10'd6};
ram[24418] = {9'd9,10'd9};
ram[24419] = {9'd12,10'd12};
ram[24420] = {9'd15,10'd15};
ram[24421] = {9'd18,10'd18};
ram[24422] = {9'd21,10'd21};
ram[24423] = {9'd25,10'd25};
ram[24424] = {9'd28,10'd28};
ram[24425] = {9'd31,10'd31};
ram[24426] = {9'd34,10'd34};
ram[24427] = {9'd37,10'd37};
ram[24428] = {9'd40,10'd40};
ram[24429] = {9'd43,10'd43};
ram[24430] = {9'd47,10'd47};
ram[24431] = {9'd50,10'd50};
ram[24432] = {9'd53,10'd53};
ram[24433] = {9'd56,10'd56};
ram[24434] = {9'd59,10'd59};
ram[24435] = {9'd62,10'd62};
ram[24436] = {9'd65,10'd65};
ram[24437] = {9'd69,10'd69};
ram[24438] = {9'd72,10'd72};
ram[24439] = {9'd75,10'd75};
ram[24440] = {9'd78,10'd78};
ram[24441] = {9'd81,10'd81};
ram[24442] = {9'd84,10'd84};
ram[24443] = {9'd87,10'd87};
ram[24444] = {9'd91,10'd91};
ram[24445] = {9'd94,10'd94};
ram[24446] = {9'd97,10'd97};
ram[24447] = {-9'd100,10'd100};
ram[24448] = {-9'd100,10'd100};
ram[24449] = {-9'd97,10'd103};
ram[24450] = {-9'd94,10'd106};
ram[24451] = {-9'd91,10'd109};
ram[24452] = {-9'd88,10'd113};
ram[24453] = {-9'd85,10'd116};
ram[24454] = {-9'd81,10'd119};
ram[24455] = {-9'd78,10'd122};
ram[24456] = {-9'd75,10'd125};
ram[24457] = {-9'd72,10'd128};
ram[24458] = {-9'd69,10'd131};
ram[24459] = {-9'd66,10'd135};
ram[24460] = {-9'd63,10'd138};
ram[24461] = {-9'd59,10'd141};
ram[24462] = {-9'd56,10'd144};
ram[24463] = {-9'd53,10'd147};
ram[24464] = {-9'd50,10'd150};
ram[24465] = {-9'd47,10'd153};
ram[24466] = {-9'd44,10'd157};
ram[24467] = {-9'd41,10'd160};
ram[24468] = {-9'd37,10'd163};
ram[24469] = {-9'd34,10'd166};
ram[24470] = {-9'd31,10'd169};
ram[24471] = {-9'd28,10'd172};
ram[24472] = {-9'd25,10'd175};
ram[24473] = {-9'd22,10'd179};
ram[24474] = {-9'd19,10'd182};
ram[24475] = {-9'd15,10'd185};
ram[24476] = {-9'd12,10'd188};
ram[24477] = {-9'd9,10'd191};
ram[24478] = {-9'd6,10'd194};
ram[24479] = {-9'd3,10'd197};
ram[24480] = {9'd0,10'd201};
ram[24481] = {9'd3,10'd204};
ram[24482] = {9'd7,10'd207};
ram[24483] = {9'd10,10'd210};
ram[24484] = {9'd13,10'd213};
ram[24485] = {9'd16,10'd216};
ram[24486] = {9'd19,10'd219};
ram[24487] = {9'd22,10'd223};
ram[24488] = {9'd25,10'd226};
ram[24489] = {9'd29,10'd229};
ram[24490] = {9'd32,10'd232};
ram[24491] = {9'd35,10'd235};
ram[24492] = {9'd38,10'd238};
ram[24493] = {9'd41,10'd241};
ram[24494] = {9'd44,10'd245};
ram[24495] = {9'd47,10'd248};
ram[24496] = {9'd51,10'd251};
ram[24497] = {9'd54,10'd254};
ram[24498] = {9'd57,10'd257};
ram[24499] = {9'd60,10'd260};
ram[24500] = {9'd63,10'd263};
ram[24501] = {9'd66,10'd267};
ram[24502] = {9'd69,10'd270};
ram[24503] = {9'd73,10'd273};
ram[24504] = {9'd76,10'd276};
ram[24505] = {9'd79,10'd279};
ram[24506] = {9'd82,10'd282};
ram[24507] = {9'd85,10'd285};
ram[24508] = {9'd88,10'd289};
ram[24509] = {9'd91,10'd292};
ram[24510] = {9'd95,10'd295};
ram[24511] = {9'd98,10'd298};
ram[24512] = {-9'd99,10'd301};
ram[24513] = {-9'd96,10'd304};
ram[24514] = {-9'd93,10'd307};
ram[24515] = {-9'd90,10'd311};
ram[24516] = {-9'd87,10'd314};
ram[24517] = {-9'd84,10'd317};
ram[24518] = {-9'd81,10'd320};
ram[24519] = {-9'd77,10'd323};
ram[24520] = {-9'd74,10'd326};
ram[24521] = {-9'd71,10'd329};
ram[24522] = {-9'd68,10'd333};
ram[24523] = {-9'd65,10'd336};
ram[24524] = {-9'd62,10'd339};
ram[24525] = {-9'd59,10'd342};
ram[24526] = {-9'd55,10'd345};
ram[24527] = {-9'd52,10'd348};
ram[24528] = {-9'd49,10'd351};
ram[24529] = {-9'd46,10'd354};
ram[24530] = {-9'd43,10'd358};
ram[24531] = {-9'd40,10'd361};
ram[24532] = {-9'd37,10'd364};
ram[24533] = {-9'd33,10'd367};
ram[24534] = {-9'd30,10'd370};
ram[24535] = {-9'd27,10'd373};
ram[24536] = {-9'd24,10'd376};
ram[24537] = {-9'd21,10'd380};
ram[24538] = {-9'd18,10'd383};
ram[24539] = {-9'd15,10'd386};
ram[24540] = {-9'd11,10'd389};
ram[24541] = {-9'd8,10'd392};
ram[24542] = {-9'd5,10'd395};
ram[24543] = {-9'd2,10'd398};
ram[24544] = {9'd1,-10'd399};
ram[24545] = {9'd4,-10'd396};
ram[24546] = {9'd7,-10'd393};
ram[24547] = {9'd10,-10'd390};
ram[24548] = {9'd14,-10'd387};
ram[24549] = {9'd17,-10'd384};
ram[24550] = {9'd20,-10'd381};
ram[24551] = {9'd23,-10'd377};
ram[24552] = {9'd26,-10'd374};
ram[24553] = {9'd29,-10'd371};
ram[24554] = {9'd32,-10'd368};
ram[24555] = {9'd36,-10'd365};
ram[24556] = {9'd39,-10'd362};
ram[24557] = {9'd42,-10'd359};
ram[24558] = {9'd45,-10'd355};
ram[24559] = {9'd48,-10'd352};
ram[24560] = {9'd51,-10'd349};
ram[24561] = {9'd54,-10'd346};
ram[24562] = {9'd58,-10'd343};
ram[24563] = {9'd61,-10'd340};
ram[24564] = {9'd64,-10'd337};
ram[24565] = {9'd67,-10'd334};
ram[24566] = {9'd70,-10'd330};
ram[24567] = {9'd73,-10'd327};
ram[24568] = {9'd76,-10'd324};
ram[24569] = {9'd80,-10'd321};
ram[24570] = {9'd83,-10'd318};
ram[24571] = {9'd86,-10'd315};
ram[24572] = {9'd89,-10'd312};
ram[24573] = {9'd92,-10'd308};
ram[24574] = {9'd95,-10'd305};
ram[24575] = {9'd98,-10'd302};
ram[24576] = {9'd98,-10'd302};
ram[24577] = {-9'd99,-10'd299};
ram[24578] = {-9'd96,-10'd296};
ram[24579] = {-9'd92,-10'd293};
ram[24580] = {-9'd89,-10'd290};
ram[24581] = {-9'd86,-10'd286};
ram[24582] = {-9'd83,-10'd283};
ram[24583] = {-9'd80,-10'd280};
ram[24584] = {-9'd77,-10'd277};
ram[24585] = {-9'd74,-10'd274};
ram[24586] = {-9'd70,-10'd271};
ram[24587] = {-9'd67,-10'd268};
ram[24588] = {-9'd64,-10'd264};
ram[24589] = {-9'd61,-10'd261};
ram[24590] = {-9'd58,-10'd258};
ram[24591] = {-9'd55,-10'd255};
ram[24592] = {-9'd52,-10'd252};
ram[24593] = {-9'd48,-10'd249};
ram[24594] = {-9'd45,-10'd246};
ram[24595] = {-9'd42,-10'd242};
ram[24596] = {-9'd39,-10'd239};
ram[24597] = {-9'd36,-10'd236};
ram[24598] = {-9'd33,-10'd233};
ram[24599] = {-9'd30,-10'd230};
ram[24600] = {-9'd26,-10'd227};
ram[24601] = {-9'd23,-10'd224};
ram[24602] = {-9'd20,-10'd220};
ram[24603] = {-9'd17,-10'd217};
ram[24604] = {-9'd14,-10'd214};
ram[24605] = {-9'd11,-10'd211};
ram[24606] = {-9'd8,-10'd208};
ram[24607] = {-9'd4,-10'd205};
ram[24608] = {-9'd1,-10'd202};
ram[24609] = {9'd2,-10'd198};
ram[24610] = {9'd5,-10'd195};
ram[24611] = {9'd8,-10'd192};
ram[24612] = {9'd11,-10'd189};
ram[24613] = {9'd14,-10'd186};
ram[24614] = {9'd18,-10'd183};
ram[24615] = {9'd21,-10'd180};
ram[24616] = {9'd24,-10'd176};
ram[24617] = {9'd27,-10'd173};
ram[24618] = {9'd30,-10'd170};
ram[24619] = {9'd33,-10'd167};
ram[24620] = {9'd36,-10'd164};
ram[24621] = {9'd40,-10'd161};
ram[24622] = {9'd43,-10'd158};
ram[24623] = {9'd46,-10'd154};
ram[24624] = {9'd49,-10'd151};
ram[24625] = {9'd52,-10'd148};
ram[24626] = {9'd55,-10'd145};
ram[24627] = {9'd58,-10'd142};
ram[24628] = {9'd62,-10'd139};
ram[24629] = {9'd65,-10'd136};
ram[24630] = {9'd68,-10'd132};
ram[24631] = {9'd71,-10'd129};
ram[24632] = {9'd74,-10'd126};
ram[24633] = {9'd77,-10'd123};
ram[24634] = {9'd80,-10'd120};
ram[24635] = {9'd84,-10'd117};
ram[24636] = {9'd87,-10'd114};
ram[24637] = {9'd90,-10'd110};
ram[24638] = {9'd93,-10'd107};
ram[24639] = {9'd96,-10'd104};
ram[24640] = {9'd99,-10'd101};
ram[24641] = {-9'd98,-10'd98};
ram[24642] = {-9'd95,-10'd95};
ram[24643] = {-9'd92,-10'd92};
ram[24644] = {-9'd88,-10'd88};
ram[24645] = {-9'd85,-10'd85};
ram[24646] = {-9'd82,-10'd82};
ram[24647] = {-9'd79,-10'd79};
ram[24648] = {-9'd76,-10'd76};
ram[24649] = {-9'd73,-10'd73};
ram[24650] = {-9'd70,-10'd70};
ram[24651] = {-9'd66,-10'd66};
ram[24652] = {-9'd63,-10'd63};
ram[24653] = {-9'd60,-10'd60};
ram[24654] = {-9'd57,-10'd57};
ram[24655] = {-9'd54,-10'd54};
ram[24656] = {-9'd51,-10'd51};
ram[24657] = {-9'd48,-10'd48};
ram[24658] = {-9'd44,-10'd44};
ram[24659] = {-9'd41,-10'd41};
ram[24660] = {-9'd38,-10'd38};
ram[24661] = {-9'd35,-10'd35};
ram[24662] = {-9'd32,-10'd32};
ram[24663] = {-9'd29,-10'd29};
ram[24664] = {-9'd26,-10'd26};
ram[24665] = {-9'd22,-10'd22};
ram[24666] = {-9'd19,-10'd19};
ram[24667] = {-9'd16,-10'd16};
ram[24668] = {-9'd13,-10'd13};
ram[24669] = {-9'd10,-10'd10};
ram[24670] = {-9'd7,-10'd7};
ram[24671] = {-9'd4,-10'd4};
ram[24672] = {9'd0,10'd0};
ram[24673] = {9'd3,10'd3};
ram[24674] = {9'd6,10'd6};
ram[24675] = {9'd9,10'd9};
ram[24676] = {9'd12,10'd12};
ram[24677] = {9'd15,10'd15};
ram[24678] = {9'd18,10'd18};
ram[24679] = {9'd21,10'd21};
ram[24680] = {9'd25,10'd25};
ram[24681] = {9'd28,10'd28};
ram[24682] = {9'd31,10'd31};
ram[24683] = {9'd34,10'd34};
ram[24684] = {9'd37,10'd37};
ram[24685] = {9'd40,10'd40};
ram[24686] = {9'd43,10'd43};
ram[24687] = {9'd47,10'd47};
ram[24688] = {9'd50,10'd50};
ram[24689] = {9'd53,10'd53};
ram[24690] = {9'd56,10'd56};
ram[24691] = {9'd59,10'd59};
ram[24692] = {9'd62,10'd62};
ram[24693] = {9'd65,10'd65};
ram[24694] = {9'd69,10'd69};
ram[24695] = {9'd72,10'd72};
ram[24696] = {9'd75,10'd75};
ram[24697] = {9'd78,10'd78};
ram[24698] = {9'd81,10'd81};
ram[24699] = {9'd84,10'd84};
ram[24700] = {9'd87,10'd87};
ram[24701] = {9'd91,10'd91};
ram[24702] = {9'd94,10'd94};
ram[24703] = {9'd97,10'd97};
ram[24704] = {9'd97,10'd97};
ram[24705] = {-9'd100,10'd100};
ram[24706] = {-9'd97,10'd103};
ram[24707] = {-9'd94,10'd106};
ram[24708] = {-9'd91,10'd109};
ram[24709] = {-9'd88,10'd113};
ram[24710] = {-9'd85,10'd116};
ram[24711] = {-9'd81,10'd119};
ram[24712] = {-9'd78,10'd122};
ram[24713] = {-9'd75,10'd125};
ram[24714] = {-9'd72,10'd128};
ram[24715] = {-9'd69,10'd131};
ram[24716] = {-9'd66,10'd135};
ram[24717] = {-9'd63,10'd138};
ram[24718] = {-9'd59,10'd141};
ram[24719] = {-9'd56,10'd144};
ram[24720] = {-9'd53,10'd147};
ram[24721] = {-9'd50,10'd150};
ram[24722] = {-9'd47,10'd153};
ram[24723] = {-9'd44,10'd157};
ram[24724] = {-9'd41,10'd160};
ram[24725] = {-9'd37,10'd163};
ram[24726] = {-9'd34,10'd166};
ram[24727] = {-9'd31,10'd169};
ram[24728] = {-9'd28,10'd172};
ram[24729] = {-9'd25,10'd175};
ram[24730] = {-9'd22,10'd179};
ram[24731] = {-9'd19,10'd182};
ram[24732] = {-9'd15,10'd185};
ram[24733] = {-9'd12,10'd188};
ram[24734] = {-9'd9,10'd191};
ram[24735] = {-9'd6,10'd194};
ram[24736] = {-9'd3,10'd197};
ram[24737] = {9'd0,10'd201};
ram[24738] = {9'd3,10'd204};
ram[24739] = {9'd7,10'd207};
ram[24740] = {9'd10,10'd210};
ram[24741] = {9'd13,10'd213};
ram[24742] = {9'd16,10'd216};
ram[24743] = {9'd19,10'd219};
ram[24744] = {9'd22,10'd223};
ram[24745] = {9'd25,10'd226};
ram[24746] = {9'd29,10'd229};
ram[24747] = {9'd32,10'd232};
ram[24748] = {9'd35,10'd235};
ram[24749] = {9'd38,10'd238};
ram[24750] = {9'd41,10'd241};
ram[24751] = {9'd44,10'd245};
ram[24752] = {9'd47,10'd248};
ram[24753] = {9'd51,10'd251};
ram[24754] = {9'd54,10'd254};
ram[24755] = {9'd57,10'd257};
ram[24756] = {9'd60,10'd260};
ram[24757] = {9'd63,10'd263};
ram[24758] = {9'd66,10'd267};
ram[24759] = {9'd69,10'd270};
ram[24760] = {9'd73,10'd273};
ram[24761] = {9'd76,10'd276};
ram[24762] = {9'd79,10'd279};
ram[24763] = {9'd82,10'd282};
ram[24764] = {9'd85,10'd285};
ram[24765] = {9'd88,10'd289};
ram[24766] = {9'd91,10'd292};
ram[24767] = {9'd95,10'd295};
ram[24768] = {9'd98,10'd298};
ram[24769] = {-9'd99,10'd301};
ram[24770] = {-9'd96,10'd304};
ram[24771] = {-9'd93,10'd307};
ram[24772] = {-9'd90,10'd311};
ram[24773] = {-9'd87,10'd314};
ram[24774] = {-9'd84,10'd317};
ram[24775] = {-9'd81,10'd320};
ram[24776] = {-9'd77,10'd323};
ram[24777] = {-9'd74,10'd326};
ram[24778] = {-9'd71,10'd329};
ram[24779] = {-9'd68,10'd333};
ram[24780] = {-9'd65,10'd336};
ram[24781] = {-9'd62,10'd339};
ram[24782] = {-9'd59,10'd342};
ram[24783] = {-9'd55,10'd345};
ram[24784] = {-9'd52,10'd348};
ram[24785] = {-9'd49,10'd351};
ram[24786] = {-9'd46,10'd354};
ram[24787] = {-9'd43,10'd358};
ram[24788] = {-9'd40,10'd361};
ram[24789] = {-9'd37,10'd364};
ram[24790] = {-9'd33,10'd367};
ram[24791] = {-9'd30,10'd370};
ram[24792] = {-9'd27,10'd373};
ram[24793] = {-9'd24,10'd376};
ram[24794] = {-9'd21,10'd380};
ram[24795] = {-9'd18,10'd383};
ram[24796] = {-9'd15,10'd386};
ram[24797] = {-9'd11,10'd389};
ram[24798] = {-9'd8,10'd392};
ram[24799] = {-9'd5,10'd395};
ram[24800] = {-9'd2,10'd398};
ram[24801] = {9'd1,-10'd399};
ram[24802] = {9'd4,-10'd396};
ram[24803] = {9'd7,-10'd393};
ram[24804] = {9'd10,-10'd390};
ram[24805] = {9'd14,-10'd387};
ram[24806] = {9'd17,-10'd384};
ram[24807] = {9'd20,-10'd381};
ram[24808] = {9'd23,-10'd377};
ram[24809] = {9'd26,-10'd374};
ram[24810] = {9'd29,-10'd371};
ram[24811] = {9'd32,-10'd368};
ram[24812] = {9'd36,-10'd365};
ram[24813] = {9'd39,-10'd362};
ram[24814] = {9'd42,-10'd359};
ram[24815] = {9'd45,-10'd355};
ram[24816] = {9'd48,-10'd352};
ram[24817] = {9'd51,-10'd349};
ram[24818] = {9'd54,-10'd346};
ram[24819] = {9'd58,-10'd343};
ram[24820] = {9'd61,-10'd340};
ram[24821] = {9'd64,-10'd337};
ram[24822] = {9'd67,-10'd334};
ram[24823] = {9'd70,-10'd330};
ram[24824] = {9'd73,-10'd327};
ram[24825] = {9'd76,-10'd324};
ram[24826] = {9'd80,-10'd321};
ram[24827] = {9'd83,-10'd318};
ram[24828] = {9'd86,-10'd315};
ram[24829] = {9'd89,-10'd312};
ram[24830] = {9'd92,-10'd308};
ram[24831] = {9'd95,-10'd305};
ram[24832] = {9'd95,-10'd305};
ram[24833] = {9'd98,-10'd302};
ram[24834] = {-9'd99,-10'd299};
ram[24835] = {-9'd96,-10'd296};
ram[24836] = {-9'd92,-10'd293};
ram[24837] = {-9'd89,-10'd290};
ram[24838] = {-9'd86,-10'd286};
ram[24839] = {-9'd83,-10'd283};
ram[24840] = {-9'd80,-10'd280};
ram[24841] = {-9'd77,-10'd277};
ram[24842] = {-9'd74,-10'd274};
ram[24843] = {-9'd70,-10'd271};
ram[24844] = {-9'd67,-10'd268};
ram[24845] = {-9'd64,-10'd264};
ram[24846] = {-9'd61,-10'd261};
ram[24847] = {-9'd58,-10'd258};
ram[24848] = {-9'd55,-10'd255};
ram[24849] = {-9'd52,-10'd252};
ram[24850] = {-9'd48,-10'd249};
ram[24851] = {-9'd45,-10'd246};
ram[24852] = {-9'd42,-10'd242};
ram[24853] = {-9'd39,-10'd239};
ram[24854] = {-9'd36,-10'd236};
ram[24855] = {-9'd33,-10'd233};
ram[24856] = {-9'd30,-10'd230};
ram[24857] = {-9'd26,-10'd227};
ram[24858] = {-9'd23,-10'd224};
ram[24859] = {-9'd20,-10'd220};
ram[24860] = {-9'd17,-10'd217};
ram[24861] = {-9'd14,-10'd214};
ram[24862] = {-9'd11,-10'd211};
ram[24863] = {-9'd8,-10'd208};
ram[24864] = {-9'd4,-10'd205};
ram[24865] = {-9'd1,-10'd202};
ram[24866] = {9'd2,-10'd198};
ram[24867] = {9'd5,-10'd195};
ram[24868] = {9'd8,-10'd192};
ram[24869] = {9'd11,-10'd189};
ram[24870] = {9'd14,-10'd186};
ram[24871] = {9'd18,-10'd183};
ram[24872] = {9'd21,-10'd180};
ram[24873] = {9'd24,-10'd176};
ram[24874] = {9'd27,-10'd173};
ram[24875] = {9'd30,-10'd170};
ram[24876] = {9'd33,-10'd167};
ram[24877] = {9'd36,-10'd164};
ram[24878] = {9'd40,-10'd161};
ram[24879] = {9'd43,-10'd158};
ram[24880] = {9'd46,-10'd154};
ram[24881] = {9'd49,-10'd151};
ram[24882] = {9'd52,-10'd148};
ram[24883] = {9'd55,-10'd145};
ram[24884] = {9'd58,-10'd142};
ram[24885] = {9'd62,-10'd139};
ram[24886] = {9'd65,-10'd136};
ram[24887] = {9'd68,-10'd132};
ram[24888] = {9'd71,-10'd129};
ram[24889] = {9'd74,-10'd126};
ram[24890] = {9'd77,-10'd123};
ram[24891] = {9'd80,-10'd120};
ram[24892] = {9'd84,-10'd117};
ram[24893] = {9'd87,-10'd114};
ram[24894] = {9'd90,-10'd110};
ram[24895] = {9'd93,-10'd107};
ram[24896] = {9'd96,-10'd104};
ram[24897] = {9'd99,-10'd101};
ram[24898] = {-9'd98,-10'd98};
ram[24899] = {-9'd95,-10'd95};
ram[24900] = {-9'd92,-10'd92};
ram[24901] = {-9'd88,-10'd88};
ram[24902] = {-9'd85,-10'd85};
ram[24903] = {-9'd82,-10'd82};
ram[24904] = {-9'd79,-10'd79};
ram[24905] = {-9'd76,-10'd76};
ram[24906] = {-9'd73,-10'd73};
ram[24907] = {-9'd70,-10'd70};
ram[24908] = {-9'd66,-10'd66};
ram[24909] = {-9'd63,-10'd63};
ram[24910] = {-9'd60,-10'd60};
ram[24911] = {-9'd57,-10'd57};
ram[24912] = {-9'd54,-10'd54};
ram[24913] = {-9'd51,-10'd51};
ram[24914] = {-9'd48,-10'd48};
ram[24915] = {-9'd44,-10'd44};
ram[24916] = {-9'd41,-10'd41};
ram[24917] = {-9'd38,-10'd38};
ram[24918] = {-9'd35,-10'd35};
ram[24919] = {-9'd32,-10'd32};
ram[24920] = {-9'd29,-10'd29};
ram[24921] = {-9'd26,-10'd26};
ram[24922] = {-9'd22,-10'd22};
ram[24923] = {-9'd19,-10'd19};
ram[24924] = {-9'd16,-10'd16};
ram[24925] = {-9'd13,-10'd13};
ram[24926] = {-9'd10,-10'd10};
ram[24927] = {-9'd7,-10'd7};
ram[24928] = {-9'd4,-10'd4};
ram[24929] = {9'd0,10'd0};
ram[24930] = {9'd3,10'd3};
ram[24931] = {9'd6,10'd6};
ram[24932] = {9'd9,10'd9};
ram[24933] = {9'd12,10'd12};
ram[24934] = {9'd15,10'd15};
ram[24935] = {9'd18,10'd18};
ram[24936] = {9'd21,10'd21};
ram[24937] = {9'd25,10'd25};
ram[24938] = {9'd28,10'd28};
ram[24939] = {9'd31,10'd31};
ram[24940] = {9'd34,10'd34};
ram[24941] = {9'd37,10'd37};
ram[24942] = {9'd40,10'd40};
ram[24943] = {9'd43,10'd43};
ram[24944] = {9'd47,10'd47};
ram[24945] = {9'd50,10'd50};
ram[24946] = {9'd53,10'd53};
ram[24947] = {9'd56,10'd56};
ram[24948] = {9'd59,10'd59};
ram[24949] = {9'd62,10'd62};
ram[24950] = {9'd65,10'd65};
ram[24951] = {9'd69,10'd69};
ram[24952] = {9'd72,10'd72};
ram[24953] = {9'd75,10'd75};
ram[24954] = {9'd78,10'd78};
ram[24955] = {9'd81,10'd81};
ram[24956] = {9'd84,10'd84};
ram[24957] = {9'd87,10'd87};
ram[24958] = {9'd91,10'd91};
ram[24959] = {9'd94,10'd94};
ram[24960] = {9'd94,10'd94};
ram[24961] = {9'd97,10'd97};
ram[24962] = {-9'd100,10'd100};
ram[24963] = {-9'd97,10'd103};
ram[24964] = {-9'd94,10'd106};
ram[24965] = {-9'd91,10'd109};
ram[24966] = {-9'd88,10'd113};
ram[24967] = {-9'd85,10'd116};
ram[24968] = {-9'd81,10'd119};
ram[24969] = {-9'd78,10'd122};
ram[24970] = {-9'd75,10'd125};
ram[24971] = {-9'd72,10'd128};
ram[24972] = {-9'd69,10'd131};
ram[24973] = {-9'd66,10'd135};
ram[24974] = {-9'd63,10'd138};
ram[24975] = {-9'd59,10'd141};
ram[24976] = {-9'd56,10'd144};
ram[24977] = {-9'd53,10'd147};
ram[24978] = {-9'd50,10'd150};
ram[24979] = {-9'd47,10'd153};
ram[24980] = {-9'd44,10'd157};
ram[24981] = {-9'd41,10'd160};
ram[24982] = {-9'd37,10'd163};
ram[24983] = {-9'd34,10'd166};
ram[24984] = {-9'd31,10'd169};
ram[24985] = {-9'd28,10'd172};
ram[24986] = {-9'd25,10'd175};
ram[24987] = {-9'd22,10'd179};
ram[24988] = {-9'd19,10'd182};
ram[24989] = {-9'd15,10'd185};
ram[24990] = {-9'd12,10'd188};
ram[24991] = {-9'd9,10'd191};
ram[24992] = {-9'd6,10'd194};
ram[24993] = {-9'd3,10'd197};
ram[24994] = {9'd0,10'd201};
ram[24995] = {9'd3,10'd204};
ram[24996] = {9'd7,10'd207};
ram[24997] = {9'd10,10'd210};
ram[24998] = {9'd13,10'd213};
ram[24999] = {9'd16,10'd216};
ram[25000] = {9'd19,10'd219};
ram[25001] = {9'd22,10'd223};
ram[25002] = {9'd25,10'd226};
ram[25003] = {9'd29,10'd229};
ram[25004] = {9'd32,10'd232};
ram[25005] = {9'd35,10'd235};
ram[25006] = {9'd38,10'd238};
ram[25007] = {9'd41,10'd241};
ram[25008] = {9'd44,10'd245};
ram[25009] = {9'd47,10'd248};
ram[25010] = {9'd51,10'd251};
ram[25011] = {9'd54,10'd254};
ram[25012] = {9'd57,10'd257};
ram[25013] = {9'd60,10'd260};
ram[25014] = {9'd63,10'd263};
ram[25015] = {9'd66,10'd267};
ram[25016] = {9'd69,10'd270};
ram[25017] = {9'd73,10'd273};
ram[25018] = {9'd76,10'd276};
ram[25019] = {9'd79,10'd279};
ram[25020] = {9'd82,10'd282};
ram[25021] = {9'd85,10'd285};
ram[25022] = {9'd88,10'd289};
ram[25023] = {9'd91,10'd292};
ram[25024] = {9'd95,10'd295};
ram[25025] = {9'd98,10'd298};
ram[25026] = {-9'd99,10'd301};
ram[25027] = {-9'd96,10'd304};
ram[25028] = {-9'd93,10'd307};
ram[25029] = {-9'd90,10'd311};
ram[25030] = {-9'd87,10'd314};
ram[25031] = {-9'd84,10'd317};
ram[25032] = {-9'd81,10'd320};
ram[25033] = {-9'd77,10'd323};
ram[25034] = {-9'd74,10'd326};
ram[25035] = {-9'd71,10'd329};
ram[25036] = {-9'd68,10'd333};
ram[25037] = {-9'd65,10'd336};
ram[25038] = {-9'd62,10'd339};
ram[25039] = {-9'd59,10'd342};
ram[25040] = {-9'd55,10'd345};
ram[25041] = {-9'd52,10'd348};
ram[25042] = {-9'd49,10'd351};
ram[25043] = {-9'd46,10'd354};
ram[25044] = {-9'd43,10'd358};
ram[25045] = {-9'd40,10'd361};
ram[25046] = {-9'd37,10'd364};
ram[25047] = {-9'd33,10'd367};
ram[25048] = {-9'd30,10'd370};
ram[25049] = {-9'd27,10'd373};
ram[25050] = {-9'd24,10'd376};
ram[25051] = {-9'd21,10'd380};
ram[25052] = {-9'd18,10'd383};
ram[25053] = {-9'd15,10'd386};
ram[25054] = {-9'd11,10'd389};
ram[25055] = {-9'd8,10'd392};
ram[25056] = {-9'd5,10'd395};
ram[25057] = {-9'd2,10'd398};
ram[25058] = {9'd1,-10'd399};
ram[25059] = {9'd4,-10'd396};
ram[25060] = {9'd7,-10'd393};
ram[25061] = {9'd10,-10'd390};
ram[25062] = {9'd14,-10'd387};
ram[25063] = {9'd17,-10'd384};
ram[25064] = {9'd20,-10'd381};
ram[25065] = {9'd23,-10'd377};
ram[25066] = {9'd26,-10'd374};
ram[25067] = {9'd29,-10'd371};
ram[25068] = {9'd32,-10'd368};
ram[25069] = {9'd36,-10'd365};
ram[25070] = {9'd39,-10'd362};
ram[25071] = {9'd42,-10'd359};
ram[25072] = {9'd45,-10'd355};
ram[25073] = {9'd48,-10'd352};
ram[25074] = {9'd51,-10'd349};
ram[25075] = {9'd54,-10'd346};
ram[25076] = {9'd58,-10'd343};
ram[25077] = {9'd61,-10'd340};
ram[25078] = {9'd64,-10'd337};
ram[25079] = {9'd67,-10'd334};
ram[25080] = {9'd70,-10'd330};
ram[25081] = {9'd73,-10'd327};
ram[25082] = {9'd76,-10'd324};
ram[25083] = {9'd80,-10'd321};
ram[25084] = {9'd83,-10'd318};
ram[25085] = {9'd86,-10'd315};
ram[25086] = {9'd89,-10'd312};
ram[25087] = {9'd92,-10'd308};
ram[25088] = {9'd92,-10'd308};
ram[25089] = {9'd95,-10'd305};
ram[25090] = {9'd98,-10'd302};
ram[25091] = {-9'd99,-10'd299};
ram[25092] = {-9'd96,-10'd296};
ram[25093] = {-9'd92,-10'd293};
ram[25094] = {-9'd89,-10'd290};
ram[25095] = {-9'd86,-10'd286};
ram[25096] = {-9'd83,-10'd283};
ram[25097] = {-9'd80,-10'd280};
ram[25098] = {-9'd77,-10'd277};
ram[25099] = {-9'd74,-10'd274};
ram[25100] = {-9'd70,-10'd271};
ram[25101] = {-9'd67,-10'd268};
ram[25102] = {-9'd64,-10'd264};
ram[25103] = {-9'd61,-10'd261};
ram[25104] = {-9'd58,-10'd258};
ram[25105] = {-9'd55,-10'd255};
ram[25106] = {-9'd52,-10'd252};
ram[25107] = {-9'd48,-10'd249};
ram[25108] = {-9'd45,-10'd246};
ram[25109] = {-9'd42,-10'd242};
ram[25110] = {-9'd39,-10'd239};
ram[25111] = {-9'd36,-10'd236};
ram[25112] = {-9'd33,-10'd233};
ram[25113] = {-9'd30,-10'd230};
ram[25114] = {-9'd26,-10'd227};
ram[25115] = {-9'd23,-10'd224};
ram[25116] = {-9'd20,-10'd220};
ram[25117] = {-9'd17,-10'd217};
ram[25118] = {-9'd14,-10'd214};
ram[25119] = {-9'd11,-10'd211};
ram[25120] = {-9'd8,-10'd208};
ram[25121] = {-9'd4,-10'd205};
ram[25122] = {-9'd1,-10'd202};
ram[25123] = {9'd2,-10'd198};
ram[25124] = {9'd5,-10'd195};
ram[25125] = {9'd8,-10'd192};
ram[25126] = {9'd11,-10'd189};
ram[25127] = {9'd14,-10'd186};
ram[25128] = {9'd18,-10'd183};
ram[25129] = {9'd21,-10'd180};
ram[25130] = {9'd24,-10'd176};
ram[25131] = {9'd27,-10'd173};
ram[25132] = {9'd30,-10'd170};
ram[25133] = {9'd33,-10'd167};
ram[25134] = {9'd36,-10'd164};
ram[25135] = {9'd40,-10'd161};
ram[25136] = {9'd43,-10'd158};
ram[25137] = {9'd46,-10'd154};
ram[25138] = {9'd49,-10'd151};
ram[25139] = {9'd52,-10'd148};
ram[25140] = {9'd55,-10'd145};
ram[25141] = {9'd58,-10'd142};
ram[25142] = {9'd62,-10'd139};
ram[25143] = {9'd65,-10'd136};
ram[25144] = {9'd68,-10'd132};
ram[25145] = {9'd71,-10'd129};
ram[25146] = {9'd74,-10'd126};
ram[25147] = {9'd77,-10'd123};
ram[25148] = {9'd80,-10'd120};
ram[25149] = {9'd84,-10'd117};
ram[25150] = {9'd87,-10'd114};
ram[25151] = {9'd90,-10'd110};
ram[25152] = {9'd93,-10'd107};
ram[25153] = {9'd96,-10'd104};
ram[25154] = {9'd99,-10'd101};
ram[25155] = {-9'd98,-10'd98};
ram[25156] = {-9'd95,-10'd95};
ram[25157] = {-9'd92,-10'd92};
ram[25158] = {-9'd88,-10'd88};
ram[25159] = {-9'd85,-10'd85};
ram[25160] = {-9'd82,-10'd82};
ram[25161] = {-9'd79,-10'd79};
ram[25162] = {-9'd76,-10'd76};
ram[25163] = {-9'd73,-10'd73};
ram[25164] = {-9'd70,-10'd70};
ram[25165] = {-9'd66,-10'd66};
ram[25166] = {-9'd63,-10'd63};
ram[25167] = {-9'd60,-10'd60};
ram[25168] = {-9'd57,-10'd57};
ram[25169] = {-9'd54,-10'd54};
ram[25170] = {-9'd51,-10'd51};
ram[25171] = {-9'd48,-10'd48};
ram[25172] = {-9'd44,-10'd44};
ram[25173] = {-9'd41,-10'd41};
ram[25174] = {-9'd38,-10'd38};
ram[25175] = {-9'd35,-10'd35};
ram[25176] = {-9'd32,-10'd32};
ram[25177] = {-9'd29,-10'd29};
ram[25178] = {-9'd26,-10'd26};
ram[25179] = {-9'd22,-10'd22};
ram[25180] = {-9'd19,-10'd19};
ram[25181] = {-9'd16,-10'd16};
ram[25182] = {-9'd13,-10'd13};
ram[25183] = {-9'd10,-10'd10};
ram[25184] = {-9'd7,-10'd7};
ram[25185] = {-9'd4,-10'd4};
ram[25186] = {9'd0,10'd0};
ram[25187] = {9'd3,10'd3};
ram[25188] = {9'd6,10'd6};
ram[25189] = {9'd9,10'd9};
ram[25190] = {9'd12,10'd12};
ram[25191] = {9'd15,10'd15};
ram[25192] = {9'd18,10'd18};
ram[25193] = {9'd21,10'd21};
ram[25194] = {9'd25,10'd25};
ram[25195] = {9'd28,10'd28};
ram[25196] = {9'd31,10'd31};
ram[25197] = {9'd34,10'd34};
ram[25198] = {9'd37,10'd37};
ram[25199] = {9'd40,10'd40};
ram[25200] = {9'd43,10'd43};
ram[25201] = {9'd47,10'd47};
ram[25202] = {9'd50,10'd50};
ram[25203] = {9'd53,10'd53};
ram[25204] = {9'd56,10'd56};
ram[25205] = {9'd59,10'd59};
ram[25206] = {9'd62,10'd62};
ram[25207] = {9'd65,10'd65};
ram[25208] = {9'd69,10'd69};
ram[25209] = {9'd72,10'd72};
ram[25210] = {9'd75,10'd75};
ram[25211] = {9'd78,10'd78};
ram[25212] = {9'd81,10'd81};
ram[25213] = {9'd84,10'd84};
ram[25214] = {9'd87,10'd87};
ram[25215] = {9'd91,10'd91};
ram[25216] = {9'd91,10'd91};
ram[25217] = {9'd94,10'd94};
ram[25218] = {9'd97,10'd97};
ram[25219] = {-9'd100,10'd100};
ram[25220] = {-9'd97,10'd103};
ram[25221] = {-9'd94,10'd106};
ram[25222] = {-9'd91,10'd109};
ram[25223] = {-9'd88,10'd113};
ram[25224] = {-9'd85,10'd116};
ram[25225] = {-9'd81,10'd119};
ram[25226] = {-9'd78,10'd122};
ram[25227] = {-9'd75,10'd125};
ram[25228] = {-9'd72,10'd128};
ram[25229] = {-9'd69,10'd131};
ram[25230] = {-9'd66,10'd135};
ram[25231] = {-9'd63,10'd138};
ram[25232] = {-9'd59,10'd141};
ram[25233] = {-9'd56,10'd144};
ram[25234] = {-9'd53,10'd147};
ram[25235] = {-9'd50,10'd150};
ram[25236] = {-9'd47,10'd153};
ram[25237] = {-9'd44,10'd157};
ram[25238] = {-9'd41,10'd160};
ram[25239] = {-9'd37,10'd163};
ram[25240] = {-9'd34,10'd166};
ram[25241] = {-9'd31,10'd169};
ram[25242] = {-9'd28,10'd172};
ram[25243] = {-9'd25,10'd175};
ram[25244] = {-9'd22,10'd179};
ram[25245] = {-9'd19,10'd182};
ram[25246] = {-9'd15,10'd185};
ram[25247] = {-9'd12,10'd188};
ram[25248] = {-9'd9,10'd191};
ram[25249] = {-9'd6,10'd194};
ram[25250] = {-9'd3,10'd197};
ram[25251] = {9'd0,10'd201};
ram[25252] = {9'd3,10'd204};
ram[25253] = {9'd7,10'd207};
ram[25254] = {9'd10,10'd210};
ram[25255] = {9'd13,10'd213};
ram[25256] = {9'd16,10'd216};
ram[25257] = {9'd19,10'd219};
ram[25258] = {9'd22,10'd223};
ram[25259] = {9'd25,10'd226};
ram[25260] = {9'd29,10'd229};
ram[25261] = {9'd32,10'd232};
ram[25262] = {9'd35,10'd235};
ram[25263] = {9'd38,10'd238};
ram[25264] = {9'd41,10'd241};
ram[25265] = {9'd44,10'd245};
ram[25266] = {9'd47,10'd248};
ram[25267] = {9'd51,10'd251};
ram[25268] = {9'd54,10'd254};
ram[25269] = {9'd57,10'd257};
ram[25270] = {9'd60,10'd260};
ram[25271] = {9'd63,10'd263};
ram[25272] = {9'd66,10'd267};
ram[25273] = {9'd69,10'd270};
ram[25274] = {9'd73,10'd273};
ram[25275] = {9'd76,10'd276};
ram[25276] = {9'd79,10'd279};
ram[25277] = {9'd82,10'd282};
ram[25278] = {9'd85,10'd285};
ram[25279] = {9'd88,10'd289};
ram[25280] = {9'd91,10'd292};
ram[25281] = {9'd95,10'd295};
ram[25282] = {9'd98,10'd298};
ram[25283] = {-9'd99,10'd301};
ram[25284] = {-9'd96,10'd304};
ram[25285] = {-9'd93,10'd307};
ram[25286] = {-9'd90,10'd311};
ram[25287] = {-9'd87,10'd314};
ram[25288] = {-9'd84,10'd317};
ram[25289] = {-9'd81,10'd320};
ram[25290] = {-9'd77,10'd323};
ram[25291] = {-9'd74,10'd326};
ram[25292] = {-9'd71,10'd329};
ram[25293] = {-9'd68,10'd333};
ram[25294] = {-9'd65,10'd336};
ram[25295] = {-9'd62,10'd339};
ram[25296] = {-9'd59,10'd342};
ram[25297] = {-9'd55,10'd345};
ram[25298] = {-9'd52,10'd348};
ram[25299] = {-9'd49,10'd351};
ram[25300] = {-9'd46,10'd354};
ram[25301] = {-9'd43,10'd358};
ram[25302] = {-9'd40,10'd361};
ram[25303] = {-9'd37,10'd364};
ram[25304] = {-9'd33,10'd367};
ram[25305] = {-9'd30,10'd370};
ram[25306] = {-9'd27,10'd373};
ram[25307] = {-9'd24,10'd376};
ram[25308] = {-9'd21,10'd380};
ram[25309] = {-9'd18,10'd383};
ram[25310] = {-9'd15,10'd386};
ram[25311] = {-9'd11,10'd389};
ram[25312] = {-9'd8,10'd392};
ram[25313] = {-9'd5,10'd395};
ram[25314] = {-9'd2,10'd398};
ram[25315] = {9'd1,-10'd399};
ram[25316] = {9'd4,-10'd396};
ram[25317] = {9'd7,-10'd393};
ram[25318] = {9'd10,-10'd390};
ram[25319] = {9'd14,-10'd387};
ram[25320] = {9'd17,-10'd384};
ram[25321] = {9'd20,-10'd381};
ram[25322] = {9'd23,-10'd377};
ram[25323] = {9'd26,-10'd374};
ram[25324] = {9'd29,-10'd371};
ram[25325] = {9'd32,-10'd368};
ram[25326] = {9'd36,-10'd365};
ram[25327] = {9'd39,-10'd362};
ram[25328] = {9'd42,-10'd359};
ram[25329] = {9'd45,-10'd355};
ram[25330] = {9'd48,-10'd352};
ram[25331] = {9'd51,-10'd349};
ram[25332] = {9'd54,-10'd346};
ram[25333] = {9'd58,-10'd343};
ram[25334] = {9'd61,-10'd340};
ram[25335] = {9'd64,-10'd337};
ram[25336] = {9'd67,-10'd334};
ram[25337] = {9'd70,-10'd330};
ram[25338] = {9'd73,-10'd327};
ram[25339] = {9'd76,-10'd324};
ram[25340] = {9'd80,-10'd321};
ram[25341] = {9'd83,-10'd318};
ram[25342] = {9'd86,-10'd315};
ram[25343] = {9'd89,-10'd312};
ram[25344] = {9'd89,-10'd312};
ram[25345] = {9'd92,-10'd308};
ram[25346] = {9'd95,-10'd305};
ram[25347] = {9'd98,-10'd302};
ram[25348] = {-9'd99,-10'd299};
ram[25349] = {-9'd96,-10'd296};
ram[25350] = {-9'd92,-10'd293};
ram[25351] = {-9'd89,-10'd290};
ram[25352] = {-9'd86,-10'd286};
ram[25353] = {-9'd83,-10'd283};
ram[25354] = {-9'd80,-10'd280};
ram[25355] = {-9'd77,-10'd277};
ram[25356] = {-9'd74,-10'd274};
ram[25357] = {-9'd70,-10'd271};
ram[25358] = {-9'd67,-10'd268};
ram[25359] = {-9'd64,-10'd264};
ram[25360] = {-9'd61,-10'd261};
ram[25361] = {-9'd58,-10'd258};
ram[25362] = {-9'd55,-10'd255};
ram[25363] = {-9'd52,-10'd252};
ram[25364] = {-9'd48,-10'd249};
ram[25365] = {-9'd45,-10'd246};
ram[25366] = {-9'd42,-10'd242};
ram[25367] = {-9'd39,-10'd239};
ram[25368] = {-9'd36,-10'd236};
ram[25369] = {-9'd33,-10'd233};
ram[25370] = {-9'd30,-10'd230};
ram[25371] = {-9'd26,-10'd227};
ram[25372] = {-9'd23,-10'd224};
ram[25373] = {-9'd20,-10'd220};
ram[25374] = {-9'd17,-10'd217};
ram[25375] = {-9'd14,-10'd214};
ram[25376] = {-9'd11,-10'd211};
ram[25377] = {-9'd8,-10'd208};
ram[25378] = {-9'd4,-10'd205};
ram[25379] = {-9'd1,-10'd202};
ram[25380] = {9'd2,-10'd198};
ram[25381] = {9'd5,-10'd195};
ram[25382] = {9'd8,-10'd192};
ram[25383] = {9'd11,-10'd189};
ram[25384] = {9'd14,-10'd186};
ram[25385] = {9'd18,-10'd183};
ram[25386] = {9'd21,-10'd180};
ram[25387] = {9'd24,-10'd176};
ram[25388] = {9'd27,-10'd173};
ram[25389] = {9'd30,-10'd170};
ram[25390] = {9'd33,-10'd167};
ram[25391] = {9'd36,-10'd164};
ram[25392] = {9'd40,-10'd161};
ram[25393] = {9'd43,-10'd158};
ram[25394] = {9'd46,-10'd154};
ram[25395] = {9'd49,-10'd151};
ram[25396] = {9'd52,-10'd148};
ram[25397] = {9'd55,-10'd145};
ram[25398] = {9'd58,-10'd142};
ram[25399] = {9'd62,-10'd139};
ram[25400] = {9'd65,-10'd136};
ram[25401] = {9'd68,-10'd132};
ram[25402] = {9'd71,-10'd129};
ram[25403] = {9'd74,-10'd126};
ram[25404] = {9'd77,-10'd123};
ram[25405] = {9'd80,-10'd120};
ram[25406] = {9'd84,-10'd117};
ram[25407] = {9'd87,-10'd114};
ram[25408] = {9'd90,-10'd110};
ram[25409] = {9'd93,-10'd107};
ram[25410] = {9'd96,-10'd104};
ram[25411] = {9'd99,-10'd101};
ram[25412] = {-9'd98,-10'd98};
ram[25413] = {-9'd95,-10'd95};
ram[25414] = {-9'd92,-10'd92};
ram[25415] = {-9'd88,-10'd88};
ram[25416] = {-9'd85,-10'd85};
ram[25417] = {-9'd82,-10'd82};
ram[25418] = {-9'd79,-10'd79};
ram[25419] = {-9'd76,-10'd76};
ram[25420] = {-9'd73,-10'd73};
ram[25421] = {-9'd70,-10'd70};
ram[25422] = {-9'd66,-10'd66};
ram[25423] = {-9'd63,-10'd63};
ram[25424] = {-9'd60,-10'd60};
ram[25425] = {-9'd57,-10'd57};
ram[25426] = {-9'd54,-10'd54};
ram[25427] = {-9'd51,-10'd51};
ram[25428] = {-9'd48,-10'd48};
ram[25429] = {-9'd44,-10'd44};
ram[25430] = {-9'd41,-10'd41};
ram[25431] = {-9'd38,-10'd38};
ram[25432] = {-9'd35,-10'd35};
ram[25433] = {-9'd32,-10'd32};
ram[25434] = {-9'd29,-10'd29};
ram[25435] = {-9'd26,-10'd26};
ram[25436] = {-9'd22,-10'd22};
ram[25437] = {-9'd19,-10'd19};
ram[25438] = {-9'd16,-10'd16};
ram[25439] = {-9'd13,-10'd13};
ram[25440] = {-9'd10,-10'd10};
ram[25441] = {-9'd7,-10'd7};
ram[25442] = {-9'd4,-10'd4};
ram[25443] = {9'd0,10'd0};
ram[25444] = {9'd3,10'd3};
ram[25445] = {9'd6,10'd6};
ram[25446] = {9'd9,10'd9};
ram[25447] = {9'd12,10'd12};
ram[25448] = {9'd15,10'd15};
ram[25449] = {9'd18,10'd18};
ram[25450] = {9'd21,10'd21};
ram[25451] = {9'd25,10'd25};
ram[25452] = {9'd28,10'd28};
ram[25453] = {9'd31,10'd31};
ram[25454] = {9'd34,10'd34};
ram[25455] = {9'd37,10'd37};
ram[25456] = {9'd40,10'd40};
ram[25457] = {9'd43,10'd43};
ram[25458] = {9'd47,10'd47};
ram[25459] = {9'd50,10'd50};
ram[25460] = {9'd53,10'd53};
ram[25461] = {9'd56,10'd56};
ram[25462] = {9'd59,10'd59};
ram[25463] = {9'd62,10'd62};
ram[25464] = {9'd65,10'd65};
ram[25465] = {9'd69,10'd69};
ram[25466] = {9'd72,10'd72};
ram[25467] = {9'd75,10'd75};
ram[25468] = {9'd78,10'd78};
ram[25469] = {9'd81,10'd81};
ram[25470] = {9'd84,10'd84};
ram[25471] = {9'd87,10'd87};
ram[25472] = {9'd87,10'd87};
ram[25473] = {9'd91,10'd91};
ram[25474] = {9'd94,10'd94};
ram[25475] = {9'd97,10'd97};
ram[25476] = {-9'd100,10'd100};
ram[25477] = {-9'd97,10'd103};
ram[25478] = {-9'd94,10'd106};
ram[25479] = {-9'd91,10'd109};
ram[25480] = {-9'd88,10'd113};
ram[25481] = {-9'd85,10'd116};
ram[25482] = {-9'd81,10'd119};
ram[25483] = {-9'd78,10'd122};
ram[25484] = {-9'd75,10'd125};
ram[25485] = {-9'd72,10'd128};
ram[25486] = {-9'd69,10'd131};
ram[25487] = {-9'd66,10'd135};
ram[25488] = {-9'd63,10'd138};
ram[25489] = {-9'd59,10'd141};
ram[25490] = {-9'd56,10'd144};
ram[25491] = {-9'd53,10'd147};
ram[25492] = {-9'd50,10'd150};
ram[25493] = {-9'd47,10'd153};
ram[25494] = {-9'd44,10'd157};
ram[25495] = {-9'd41,10'd160};
ram[25496] = {-9'd37,10'd163};
ram[25497] = {-9'd34,10'd166};
ram[25498] = {-9'd31,10'd169};
ram[25499] = {-9'd28,10'd172};
ram[25500] = {-9'd25,10'd175};
ram[25501] = {-9'd22,10'd179};
ram[25502] = {-9'd19,10'd182};
ram[25503] = {-9'd15,10'd185};
ram[25504] = {-9'd12,10'd188};
ram[25505] = {-9'd9,10'd191};
ram[25506] = {-9'd6,10'd194};
ram[25507] = {-9'd3,10'd197};
ram[25508] = {9'd0,10'd201};
ram[25509] = {9'd3,10'd204};
ram[25510] = {9'd7,10'd207};
ram[25511] = {9'd10,10'd210};
ram[25512] = {9'd13,10'd213};
ram[25513] = {9'd16,10'd216};
ram[25514] = {9'd19,10'd219};
ram[25515] = {9'd22,10'd223};
ram[25516] = {9'd25,10'd226};
ram[25517] = {9'd29,10'd229};
ram[25518] = {9'd32,10'd232};
ram[25519] = {9'd35,10'd235};
ram[25520] = {9'd38,10'd238};
ram[25521] = {9'd41,10'd241};
ram[25522] = {9'd44,10'd245};
ram[25523] = {9'd47,10'd248};
ram[25524] = {9'd51,10'd251};
ram[25525] = {9'd54,10'd254};
ram[25526] = {9'd57,10'd257};
ram[25527] = {9'd60,10'd260};
ram[25528] = {9'd63,10'd263};
ram[25529] = {9'd66,10'd267};
ram[25530] = {9'd69,10'd270};
ram[25531] = {9'd73,10'd273};
ram[25532] = {9'd76,10'd276};
ram[25533] = {9'd79,10'd279};
ram[25534] = {9'd82,10'd282};
ram[25535] = {9'd85,10'd285};
ram[25536] = {9'd88,10'd289};
ram[25537] = {9'd91,10'd292};
ram[25538] = {9'd95,10'd295};
ram[25539] = {9'd98,10'd298};
ram[25540] = {-9'd99,10'd301};
ram[25541] = {-9'd96,10'd304};
ram[25542] = {-9'd93,10'd307};
ram[25543] = {-9'd90,10'd311};
ram[25544] = {-9'd87,10'd314};
ram[25545] = {-9'd84,10'd317};
ram[25546] = {-9'd81,10'd320};
ram[25547] = {-9'd77,10'd323};
ram[25548] = {-9'd74,10'd326};
ram[25549] = {-9'd71,10'd329};
ram[25550] = {-9'd68,10'd333};
ram[25551] = {-9'd65,10'd336};
ram[25552] = {-9'd62,10'd339};
ram[25553] = {-9'd59,10'd342};
ram[25554] = {-9'd55,10'd345};
ram[25555] = {-9'd52,10'd348};
ram[25556] = {-9'd49,10'd351};
ram[25557] = {-9'd46,10'd354};
ram[25558] = {-9'd43,10'd358};
ram[25559] = {-9'd40,10'd361};
ram[25560] = {-9'd37,10'd364};
ram[25561] = {-9'd33,10'd367};
ram[25562] = {-9'd30,10'd370};
ram[25563] = {-9'd27,10'd373};
ram[25564] = {-9'd24,10'd376};
ram[25565] = {-9'd21,10'd380};
ram[25566] = {-9'd18,10'd383};
ram[25567] = {-9'd15,10'd386};
ram[25568] = {-9'd11,10'd389};
ram[25569] = {-9'd8,10'd392};
ram[25570] = {-9'd5,10'd395};
ram[25571] = {-9'd2,10'd398};
ram[25572] = {9'd1,-10'd399};
ram[25573] = {9'd4,-10'd396};
ram[25574] = {9'd7,-10'd393};
ram[25575] = {9'd10,-10'd390};
ram[25576] = {9'd14,-10'd387};
ram[25577] = {9'd17,-10'd384};
ram[25578] = {9'd20,-10'd381};
ram[25579] = {9'd23,-10'd377};
ram[25580] = {9'd26,-10'd374};
ram[25581] = {9'd29,-10'd371};
ram[25582] = {9'd32,-10'd368};
ram[25583] = {9'd36,-10'd365};
ram[25584] = {9'd39,-10'd362};
ram[25585] = {9'd42,-10'd359};
ram[25586] = {9'd45,-10'd355};
ram[25587] = {9'd48,-10'd352};
ram[25588] = {9'd51,-10'd349};
ram[25589] = {9'd54,-10'd346};
ram[25590] = {9'd58,-10'd343};
ram[25591] = {9'd61,-10'd340};
ram[25592] = {9'd64,-10'd337};
ram[25593] = {9'd67,-10'd334};
ram[25594] = {9'd70,-10'd330};
ram[25595] = {9'd73,-10'd327};
ram[25596] = {9'd76,-10'd324};
ram[25597] = {9'd80,-10'd321};
ram[25598] = {9'd83,-10'd318};
ram[25599] = {9'd86,-10'd315};
ram[25600] = {9'd86,-10'd315};
ram[25601] = {9'd89,-10'd312};
ram[25602] = {9'd92,-10'd308};
ram[25603] = {9'd95,-10'd305};
ram[25604] = {9'd98,-10'd302};
ram[25605] = {-9'd99,-10'd299};
ram[25606] = {-9'd96,-10'd296};
ram[25607] = {-9'd92,-10'd293};
ram[25608] = {-9'd89,-10'd290};
ram[25609] = {-9'd86,-10'd286};
ram[25610] = {-9'd83,-10'd283};
ram[25611] = {-9'd80,-10'd280};
ram[25612] = {-9'd77,-10'd277};
ram[25613] = {-9'd74,-10'd274};
ram[25614] = {-9'd70,-10'd271};
ram[25615] = {-9'd67,-10'd268};
ram[25616] = {-9'd64,-10'd264};
ram[25617] = {-9'd61,-10'd261};
ram[25618] = {-9'd58,-10'd258};
ram[25619] = {-9'd55,-10'd255};
ram[25620] = {-9'd52,-10'd252};
ram[25621] = {-9'd48,-10'd249};
ram[25622] = {-9'd45,-10'd246};
ram[25623] = {-9'd42,-10'd242};
ram[25624] = {-9'd39,-10'd239};
ram[25625] = {-9'd36,-10'd236};
ram[25626] = {-9'd33,-10'd233};
ram[25627] = {-9'd30,-10'd230};
ram[25628] = {-9'd26,-10'd227};
ram[25629] = {-9'd23,-10'd224};
ram[25630] = {-9'd20,-10'd220};
ram[25631] = {-9'd17,-10'd217};
ram[25632] = {-9'd14,-10'd214};
ram[25633] = {-9'd11,-10'd211};
ram[25634] = {-9'd8,-10'd208};
ram[25635] = {-9'd4,-10'd205};
ram[25636] = {-9'd1,-10'd202};
ram[25637] = {9'd2,-10'd198};
ram[25638] = {9'd5,-10'd195};
ram[25639] = {9'd8,-10'd192};
ram[25640] = {9'd11,-10'd189};
ram[25641] = {9'd14,-10'd186};
ram[25642] = {9'd18,-10'd183};
ram[25643] = {9'd21,-10'd180};
ram[25644] = {9'd24,-10'd176};
ram[25645] = {9'd27,-10'd173};
ram[25646] = {9'd30,-10'd170};
ram[25647] = {9'd33,-10'd167};
ram[25648] = {9'd36,-10'd164};
ram[25649] = {9'd40,-10'd161};
ram[25650] = {9'd43,-10'd158};
ram[25651] = {9'd46,-10'd154};
ram[25652] = {9'd49,-10'd151};
ram[25653] = {9'd52,-10'd148};
ram[25654] = {9'd55,-10'd145};
ram[25655] = {9'd58,-10'd142};
ram[25656] = {9'd62,-10'd139};
ram[25657] = {9'd65,-10'd136};
ram[25658] = {9'd68,-10'd132};
ram[25659] = {9'd71,-10'd129};
ram[25660] = {9'd74,-10'd126};
ram[25661] = {9'd77,-10'd123};
ram[25662] = {9'd80,-10'd120};
ram[25663] = {9'd84,-10'd117};
ram[25664] = {9'd87,-10'd114};
ram[25665] = {9'd90,-10'd110};
ram[25666] = {9'd93,-10'd107};
ram[25667] = {9'd96,-10'd104};
ram[25668] = {9'd99,-10'd101};
ram[25669] = {-9'd98,-10'd98};
ram[25670] = {-9'd95,-10'd95};
ram[25671] = {-9'd92,-10'd92};
ram[25672] = {-9'd88,-10'd88};
ram[25673] = {-9'd85,-10'd85};
ram[25674] = {-9'd82,-10'd82};
ram[25675] = {-9'd79,-10'd79};
ram[25676] = {-9'd76,-10'd76};
ram[25677] = {-9'd73,-10'd73};
ram[25678] = {-9'd70,-10'd70};
ram[25679] = {-9'd66,-10'd66};
ram[25680] = {-9'd63,-10'd63};
ram[25681] = {-9'd60,-10'd60};
ram[25682] = {-9'd57,-10'd57};
ram[25683] = {-9'd54,-10'd54};
ram[25684] = {-9'd51,-10'd51};
ram[25685] = {-9'd48,-10'd48};
ram[25686] = {-9'd44,-10'd44};
ram[25687] = {-9'd41,-10'd41};
ram[25688] = {-9'd38,-10'd38};
ram[25689] = {-9'd35,-10'd35};
ram[25690] = {-9'd32,-10'd32};
ram[25691] = {-9'd29,-10'd29};
ram[25692] = {-9'd26,-10'd26};
ram[25693] = {-9'd22,-10'd22};
ram[25694] = {-9'd19,-10'd19};
ram[25695] = {-9'd16,-10'd16};
ram[25696] = {-9'd13,-10'd13};
ram[25697] = {-9'd10,-10'd10};
ram[25698] = {-9'd7,-10'd7};
ram[25699] = {-9'd4,-10'd4};
ram[25700] = {9'd0,10'd0};
ram[25701] = {9'd3,10'd3};
ram[25702] = {9'd6,10'd6};
ram[25703] = {9'd9,10'd9};
ram[25704] = {9'd12,10'd12};
ram[25705] = {9'd15,10'd15};
ram[25706] = {9'd18,10'd18};
ram[25707] = {9'd21,10'd21};
ram[25708] = {9'd25,10'd25};
ram[25709] = {9'd28,10'd28};
ram[25710] = {9'd31,10'd31};
ram[25711] = {9'd34,10'd34};
ram[25712] = {9'd37,10'd37};
ram[25713] = {9'd40,10'd40};
ram[25714] = {9'd43,10'd43};
ram[25715] = {9'd47,10'd47};
ram[25716] = {9'd50,10'd50};
ram[25717] = {9'd53,10'd53};
ram[25718] = {9'd56,10'd56};
ram[25719] = {9'd59,10'd59};
ram[25720] = {9'd62,10'd62};
ram[25721] = {9'd65,10'd65};
ram[25722] = {9'd69,10'd69};
ram[25723] = {9'd72,10'd72};
ram[25724] = {9'd75,10'd75};
ram[25725] = {9'd78,10'd78};
ram[25726] = {9'd81,10'd81};
ram[25727] = {9'd84,10'd84};
ram[25728] = {9'd84,10'd84};
ram[25729] = {9'd87,10'd87};
ram[25730] = {9'd91,10'd91};
ram[25731] = {9'd94,10'd94};
ram[25732] = {9'd97,10'd97};
ram[25733] = {-9'd100,10'd100};
ram[25734] = {-9'd97,10'd103};
ram[25735] = {-9'd94,10'd106};
ram[25736] = {-9'd91,10'd109};
ram[25737] = {-9'd88,10'd113};
ram[25738] = {-9'd85,10'd116};
ram[25739] = {-9'd81,10'd119};
ram[25740] = {-9'd78,10'd122};
ram[25741] = {-9'd75,10'd125};
ram[25742] = {-9'd72,10'd128};
ram[25743] = {-9'd69,10'd131};
ram[25744] = {-9'd66,10'd135};
ram[25745] = {-9'd63,10'd138};
ram[25746] = {-9'd59,10'd141};
ram[25747] = {-9'd56,10'd144};
ram[25748] = {-9'd53,10'd147};
ram[25749] = {-9'd50,10'd150};
ram[25750] = {-9'd47,10'd153};
ram[25751] = {-9'd44,10'd157};
ram[25752] = {-9'd41,10'd160};
ram[25753] = {-9'd37,10'd163};
ram[25754] = {-9'd34,10'd166};
ram[25755] = {-9'd31,10'd169};
ram[25756] = {-9'd28,10'd172};
ram[25757] = {-9'd25,10'd175};
ram[25758] = {-9'd22,10'd179};
ram[25759] = {-9'd19,10'd182};
ram[25760] = {-9'd15,10'd185};
ram[25761] = {-9'd12,10'd188};
ram[25762] = {-9'd9,10'd191};
ram[25763] = {-9'd6,10'd194};
ram[25764] = {-9'd3,10'd197};
ram[25765] = {9'd0,10'd201};
ram[25766] = {9'd3,10'd204};
ram[25767] = {9'd7,10'd207};
ram[25768] = {9'd10,10'd210};
ram[25769] = {9'd13,10'd213};
ram[25770] = {9'd16,10'd216};
ram[25771] = {9'd19,10'd219};
ram[25772] = {9'd22,10'd223};
ram[25773] = {9'd25,10'd226};
ram[25774] = {9'd29,10'd229};
ram[25775] = {9'd32,10'd232};
ram[25776] = {9'd35,10'd235};
ram[25777] = {9'd38,10'd238};
ram[25778] = {9'd41,10'd241};
ram[25779] = {9'd44,10'd245};
ram[25780] = {9'd47,10'd248};
ram[25781] = {9'd51,10'd251};
ram[25782] = {9'd54,10'd254};
ram[25783] = {9'd57,10'd257};
ram[25784] = {9'd60,10'd260};
ram[25785] = {9'd63,10'd263};
ram[25786] = {9'd66,10'd267};
ram[25787] = {9'd69,10'd270};
ram[25788] = {9'd73,10'd273};
ram[25789] = {9'd76,10'd276};
ram[25790] = {9'd79,10'd279};
ram[25791] = {9'd82,10'd282};
ram[25792] = {9'd85,10'd285};
ram[25793] = {9'd88,10'd289};
ram[25794] = {9'd91,10'd292};
ram[25795] = {9'd95,10'd295};
ram[25796] = {9'd98,10'd298};
ram[25797] = {-9'd99,10'd301};
ram[25798] = {-9'd96,10'd304};
ram[25799] = {-9'd93,10'd307};
ram[25800] = {-9'd90,10'd311};
ram[25801] = {-9'd87,10'd314};
ram[25802] = {-9'd84,10'd317};
ram[25803] = {-9'd81,10'd320};
ram[25804] = {-9'd77,10'd323};
ram[25805] = {-9'd74,10'd326};
ram[25806] = {-9'd71,10'd329};
ram[25807] = {-9'd68,10'd333};
ram[25808] = {-9'd65,10'd336};
ram[25809] = {-9'd62,10'd339};
ram[25810] = {-9'd59,10'd342};
ram[25811] = {-9'd55,10'd345};
ram[25812] = {-9'd52,10'd348};
ram[25813] = {-9'd49,10'd351};
ram[25814] = {-9'd46,10'd354};
ram[25815] = {-9'd43,10'd358};
ram[25816] = {-9'd40,10'd361};
ram[25817] = {-9'd37,10'd364};
ram[25818] = {-9'd33,10'd367};
ram[25819] = {-9'd30,10'd370};
ram[25820] = {-9'd27,10'd373};
ram[25821] = {-9'd24,10'd376};
ram[25822] = {-9'd21,10'd380};
ram[25823] = {-9'd18,10'd383};
ram[25824] = {-9'd15,10'd386};
ram[25825] = {-9'd11,10'd389};
ram[25826] = {-9'd8,10'd392};
ram[25827] = {-9'd5,10'd395};
ram[25828] = {-9'd2,10'd398};
ram[25829] = {9'd1,-10'd399};
ram[25830] = {9'd4,-10'd396};
ram[25831] = {9'd7,-10'd393};
ram[25832] = {9'd10,-10'd390};
ram[25833] = {9'd14,-10'd387};
ram[25834] = {9'd17,-10'd384};
ram[25835] = {9'd20,-10'd381};
ram[25836] = {9'd23,-10'd377};
ram[25837] = {9'd26,-10'd374};
ram[25838] = {9'd29,-10'd371};
ram[25839] = {9'd32,-10'd368};
ram[25840] = {9'd36,-10'd365};
ram[25841] = {9'd39,-10'd362};
ram[25842] = {9'd42,-10'd359};
ram[25843] = {9'd45,-10'd355};
ram[25844] = {9'd48,-10'd352};
ram[25845] = {9'd51,-10'd349};
ram[25846] = {9'd54,-10'd346};
ram[25847] = {9'd58,-10'd343};
ram[25848] = {9'd61,-10'd340};
ram[25849] = {9'd64,-10'd337};
ram[25850] = {9'd67,-10'd334};
ram[25851] = {9'd70,-10'd330};
ram[25852] = {9'd73,-10'd327};
ram[25853] = {9'd76,-10'd324};
ram[25854] = {9'd80,-10'd321};
ram[25855] = {9'd83,-10'd318};
ram[25856] = {9'd83,-10'd318};
ram[25857] = {9'd86,-10'd315};
ram[25858] = {9'd89,-10'd312};
ram[25859] = {9'd92,-10'd308};
ram[25860] = {9'd95,-10'd305};
ram[25861] = {9'd98,-10'd302};
ram[25862] = {-9'd99,-10'd299};
ram[25863] = {-9'd96,-10'd296};
ram[25864] = {-9'd92,-10'd293};
ram[25865] = {-9'd89,-10'd290};
ram[25866] = {-9'd86,-10'd286};
ram[25867] = {-9'd83,-10'd283};
ram[25868] = {-9'd80,-10'd280};
ram[25869] = {-9'd77,-10'd277};
ram[25870] = {-9'd74,-10'd274};
ram[25871] = {-9'd70,-10'd271};
ram[25872] = {-9'd67,-10'd268};
ram[25873] = {-9'd64,-10'd264};
ram[25874] = {-9'd61,-10'd261};
ram[25875] = {-9'd58,-10'd258};
ram[25876] = {-9'd55,-10'd255};
ram[25877] = {-9'd52,-10'd252};
ram[25878] = {-9'd48,-10'd249};
ram[25879] = {-9'd45,-10'd246};
ram[25880] = {-9'd42,-10'd242};
ram[25881] = {-9'd39,-10'd239};
ram[25882] = {-9'd36,-10'd236};
ram[25883] = {-9'd33,-10'd233};
ram[25884] = {-9'd30,-10'd230};
ram[25885] = {-9'd26,-10'd227};
ram[25886] = {-9'd23,-10'd224};
ram[25887] = {-9'd20,-10'd220};
ram[25888] = {-9'd17,-10'd217};
ram[25889] = {-9'd14,-10'd214};
ram[25890] = {-9'd11,-10'd211};
ram[25891] = {-9'd8,-10'd208};
ram[25892] = {-9'd4,-10'd205};
ram[25893] = {-9'd1,-10'd202};
ram[25894] = {9'd2,-10'd198};
ram[25895] = {9'd5,-10'd195};
ram[25896] = {9'd8,-10'd192};
ram[25897] = {9'd11,-10'd189};
ram[25898] = {9'd14,-10'd186};
ram[25899] = {9'd18,-10'd183};
ram[25900] = {9'd21,-10'd180};
ram[25901] = {9'd24,-10'd176};
ram[25902] = {9'd27,-10'd173};
ram[25903] = {9'd30,-10'd170};
ram[25904] = {9'd33,-10'd167};
ram[25905] = {9'd36,-10'd164};
ram[25906] = {9'd40,-10'd161};
ram[25907] = {9'd43,-10'd158};
ram[25908] = {9'd46,-10'd154};
ram[25909] = {9'd49,-10'd151};
ram[25910] = {9'd52,-10'd148};
ram[25911] = {9'd55,-10'd145};
ram[25912] = {9'd58,-10'd142};
ram[25913] = {9'd62,-10'd139};
ram[25914] = {9'd65,-10'd136};
ram[25915] = {9'd68,-10'd132};
ram[25916] = {9'd71,-10'd129};
ram[25917] = {9'd74,-10'd126};
ram[25918] = {9'd77,-10'd123};
ram[25919] = {9'd80,-10'd120};
ram[25920] = {9'd84,-10'd117};
ram[25921] = {9'd87,-10'd114};
ram[25922] = {9'd90,-10'd110};
ram[25923] = {9'd93,-10'd107};
ram[25924] = {9'd96,-10'd104};
ram[25925] = {9'd99,-10'd101};
ram[25926] = {-9'd98,-10'd98};
ram[25927] = {-9'd95,-10'd95};
ram[25928] = {-9'd92,-10'd92};
ram[25929] = {-9'd88,-10'd88};
ram[25930] = {-9'd85,-10'd85};
ram[25931] = {-9'd82,-10'd82};
ram[25932] = {-9'd79,-10'd79};
ram[25933] = {-9'd76,-10'd76};
ram[25934] = {-9'd73,-10'd73};
ram[25935] = {-9'd70,-10'd70};
ram[25936] = {-9'd66,-10'd66};
ram[25937] = {-9'd63,-10'd63};
ram[25938] = {-9'd60,-10'd60};
ram[25939] = {-9'd57,-10'd57};
ram[25940] = {-9'd54,-10'd54};
ram[25941] = {-9'd51,-10'd51};
ram[25942] = {-9'd48,-10'd48};
ram[25943] = {-9'd44,-10'd44};
ram[25944] = {-9'd41,-10'd41};
ram[25945] = {-9'd38,-10'd38};
ram[25946] = {-9'd35,-10'd35};
ram[25947] = {-9'd32,-10'd32};
ram[25948] = {-9'd29,-10'd29};
ram[25949] = {-9'd26,-10'd26};
ram[25950] = {-9'd22,-10'd22};
ram[25951] = {-9'd19,-10'd19};
ram[25952] = {-9'd16,-10'd16};
ram[25953] = {-9'd13,-10'd13};
ram[25954] = {-9'd10,-10'd10};
ram[25955] = {-9'd7,-10'd7};
ram[25956] = {-9'd4,-10'd4};
ram[25957] = {9'd0,10'd0};
ram[25958] = {9'd3,10'd3};
ram[25959] = {9'd6,10'd6};
ram[25960] = {9'd9,10'd9};
ram[25961] = {9'd12,10'd12};
ram[25962] = {9'd15,10'd15};
ram[25963] = {9'd18,10'd18};
ram[25964] = {9'd21,10'd21};
ram[25965] = {9'd25,10'd25};
ram[25966] = {9'd28,10'd28};
ram[25967] = {9'd31,10'd31};
ram[25968] = {9'd34,10'd34};
ram[25969] = {9'd37,10'd37};
ram[25970] = {9'd40,10'd40};
ram[25971] = {9'd43,10'd43};
ram[25972] = {9'd47,10'd47};
ram[25973] = {9'd50,10'd50};
ram[25974] = {9'd53,10'd53};
ram[25975] = {9'd56,10'd56};
ram[25976] = {9'd59,10'd59};
ram[25977] = {9'd62,10'd62};
ram[25978] = {9'd65,10'd65};
ram[25979] = {9'd69,10'd69};
ram[25980] = {9'd72,10'd72};
ram[25981] = {9'd75,10'd75};
ram[25982] = {9'd78,10'd78};
ram[25983] = {9'd81,10'd81};
ram[25984] = {9'd81,10'd81};
ram[25985] = {9'd84,10'd84};
ram[25986] = {9'd87,10'd87};
ram[25987] = {9'd91,10'd91};
ram[25988] = {9'd94,10'd94};
ram[25989] = {9'd97,10'd97};
ram[25990] = {-9'd100,10'd100};
ram[25991] = {-9'd97,10'd103};
ram[25992] = {-9'd94,10'd106};
ram[25993] = {-9'd91,10'd109};
ram[25994] = {-9'd88,10'd113};
ram[25995] = {-9'd85,10'd116};
ram[25996] = {-9'd81,10'd119};
ram[25997] = {-9'd78,10'd122};
ram[25998] = {-9'd75,10'd125};
ram[25999] = {-9'd72,10'd128};
ram[26000] = {-9'd69,10'd131};
ram[26001] = {-9'd66,10'd135};
ram[26002] = {-9'd63,10'd138};
ram[26003] = {-9'd59,10'd141};
ram[26004] = {-9'd56,10'd144};
ram[26005] = {-9'd53,10'd147};
ram[26006] = {-9'd50,10'd150};
ram[26007] = {-9'd47,10'd153};
ram[26008] = {-9'd44,10'd157};
ram[26009] = {-9'd41,10'd160};
ram[26010] = {-9'd37,10'd163};
ram[26011] = {-9'd34,10'd166};
ram[26012] = {-9'd31,10'd169};
ram[26013] = {-9'd28,10'd172};
ram[26014] = {-9'd25,10'd175};
ram[26015] = {-9'd22,10'd179};
ram[26016] = {-9'd19,10'd182};
ram[26017] = {-9'd15,10'd185};
ram[26018] = {-9'd12,10'd188};
ram[26019] = {-9'd9,10'd191};
ram[26020] = {-9'd6,10'd194};
ram[26021] = {-9'd3,10'd197};
ram[26022] = {9'd0,10'd201};
ram[26023] = {9'd3,10'd204};
ram[26024] = {9'd7,10'd207};
ram[26025] = {9'd10,10'd210};
ram[26026] = {9'd13,10'd213};
ram[26027] = {9'd16,10'd216};
ram[26028] = {9'd19,10'd219};
ram[26029] = {9'd22,10'd223};
ram[26030] = {9'd25,10'd226};
ram[26031] = {9'd29,10'd229};
ram[26032] = {9'd32,10'd232};
ram[26033] = {9'd35,10'd235};
ram[26034] = {9'd38,10'd238};
ram[26035] = {9'd41,10'd241};
ram[26036] = {9'd44,10'd245};
ram[26037] = {9'd47,10'd248};
ram[26038] = {9'd51,10'd251};
ram[26039] = {9'd54,10'd254};
ram[26040] = {9'd57,10'd257};
ram[26041] = {9'd60,10'd260};
ram[26042] = {9'd63,10'd263};
ram[26043] = {9'd66,10'd267};
ram[26044] = {9'd69,10'd270};
ram[26045] = {9'd73,10'd273};
ram[26046] = {9'd76,10'd276};
ram[26047] = {9'd79,10'd279};
ram[26048] = {9'd82,10'd282};
ram[26049] = {9'd85,10'd285};
ram[26050] = {9'd88,10'd289};
ram[26051] = {9'd91,10'd292};
ram[26052] = {9'd95,10'd295};
ram[26053] = {9'd98,10'd298};
ram[26054] = {-9'd99,10'd301};
ram[26055] = {-9'd96,10'd304};
ram[26056] = {-9'd93,10'd307};
ram[26057] = {-9'd90,10'd311};
ram[26058] = {-9'd87,10'd314};
ram[26059] = {-9'd84,10'd317};
ram[26060] = {-9'd81,10'd320};
ram[26061] = {-9'd77,10'd323};
ram[26062] = {-9'd74,10'd326};
ram[26063] = {-9'd71,10'd329};
ram[26064] = {-9'd68,10'd333};
ram[26065] = {-9'd65,10'd336};
ram[26066] = {-9'd62,10'd339};
ram[26067] = {-9'd59,10'd342};
ram[26068] = {-9'd55,10'd345};
ram[26069] = {-9'd52,10'd348};
ram[26070] = {-9'd49,10'd351};
ram[26071] = {-9'd46,10'd354};
ram[26072] = {-9'd43,10'd358};
ram[26073] = {-9'd40,10'd361};
ram[26074] = {-9'd37,10'd364};
ram[26075] = {-9'd33,10'd367};
ram[26076] = {-9'd30,10'd370};
ram[26077] = {-9'd27,10'd373};
ram[26078] = {-9'd24,10'd376};
ram[26079] = {-9'd21,10'd380};
ram[26080] = {-9'd18,10'd383};
ram[26081] = {-9'd15,10'd386};
ram[26082] = {-9'd11,10'd389};
ram[26083] = {-9'd8,10'd392};
ram[26084] = {-9'd5,10'd395};
ram[26085] = {-9'd2,10'd398};
ram[26086] = {9'd1,-10'd399};
ram[26087] = {9'd4,-10'd396};
ram[26088] = {9'd7,-10'd393};
ram[26089] = {9'd10,-10'd390};
ram[26090] = {9'd14,-10'd387};
ram[26091] = {9'd17,-10'd384};
ram[26092] = {9'd20,-10'd381};
ram[26093] = {9'd23,-10'd377};
ram[26094] = {9'd26,-10'd374};
ram[26095] = {9'd29,-10'd371};
ram[26096] = {9'd32,-10'd368};
ram[26097] = {9'd36,-10'd365};
ram[26098] = {9'd39,-10'd362};
ram[26099] = {9'd42,-10'd359};
ram[26100] = {9'd45,-10'd355};
ram[26101] = {9'd48,-10'd352};
ram[26102] = {9'd51,-10'd349};
ram[26103] = {9'd54,-10'd346};
ram[26104] = {9'd58,-10'd343};
ram[26105] = {9'd61,-10'd340};
ram[26106] = {9'd64,-10'd337};
ram[26107] = {9'd67,-10'd334};
ram[26108] = {9'd70,-10'd330};
ram[26109] = {9'd73,-10'd327};
ram[26110] = {9'd76,-10'd324};
ram[26111] = {9'd80,-10'd321};
ram[26112] = {9'd80,-10'd321};
ram[26113] = {9'd83,-10'd318};
ram[26114] = {9'd86,-10'd315};
ram[26115] = {9'd89,-10'd312};
ram[26116] = {9'd92,-10'd308};
ram[26117] = {9'd95,-10'd305};
ram[26118] = {9'd98,-10'd302};
ram[26119] = {-9'd99,-10'd299};
ram[26120] = {-9'd96,-10'd296};
ram[26121] = {-9'd92,-10'd293};
ram[26122] = {-9'd89,-10'd290};
ram[26123] = {-9'd86,-10'd286};
ram[26124] = {-9'd83,-10'd283};
ram[26125] = {-9'd80,-10'd280};
ram[26126] = {-9'd77,-10'd277};
ram[26127] = {-9'd74,-10'd274};
ram[26128] = {-9'd70,-10'd271};
ram[26129] = {-9'd67,-10'd268};
ram[26130] = {-9'd64,-10'd264};
ram[26131] = {-9'd61,-10'd261};
ram[26132] = {-9'd58,-10'd258};
ram[26133] = {-9'd55,-10'd255};
ram[26134] = {-9'd52,-10'd252};
ram[26135] = {-9'd48,-10'd249};
ram[26136] = {-9'd45,-10'd246};
ram[26137] = {-9'd42,-10'd242};
ram[26138] = {-9'd39,-10'd239};
ram[26139] = {-9'd36,-10'd236};
ram[26140] = {-9'd33,-10'd233};
ram[26141] = {-9'd30,-10'd230};
ram[26142] = {-9'd26,-10'd227};
ram[26143] = {-9'd23,-10'd224};
ram[26144] = {-9'd20,-10'd220};
ram[26145] = {-9'd17,-10'd217};
ram[26146] = {-9'd14,-10'd214};
ram[26147] = {-9'd11,-10'd211};
ram[26148] = {-9'd8,-10'd208};
ram[26149] = {-9'd4,-10'd205};
ram[26150] = {-9'd1,-10'd202};
ram[26151] = {9'd2,-10'd198};
ram[26152] = {9'd5,-10'd195};
ram[26153] = {9'd8,-10'd192};
ram[26154] = {9'd11,-10'd189};
ram[26155] = {9'd14,-10'd186};
ram[26156] = {9'd18,-10'd183};
ram[26157] = {9'd21,-10'd180};
ram[26158] = {9'd24,-10'd176};
ram[26159] = {9'd27,-10'd173};
ram[26160] = {9'd30,-10'd170};
ram[26161] = {9'd33,-10'd167};
ram[26162] = {9'd36,-10'd164};
ram[26163] = {9'd40,-10'd161};
ram[26164] = {9'd43,-10'd158};
ram[26165] = {9'd46,-10'd154};
ram[26166] = {9'd49,-10'd151};
ram[26167] = {9'd52,-10'd148};
ram[26168] = {9'd55,-10'd145};
ram[26169] = {9'd58,-10'd142};
ram[26170] = {9'd62,-10'd139};
ram[26171] = {9'd65,-10'd136};
ram[26172] = {9'd68,-10'd132};
ram[26173] = {9'd71,-10'd129};
ram[26174] = {9'd74,-10'd126};
ram[26175] = {9'd77,-10'd123};
ram[26176] = {9'd80,-10'd120};
ram[26177] = {9'd84,-10'd117};
ram[26178] = {9'd87,-10'd114};
ram[26179] = {9'd90,-10'd110};
ram[26180] = {9'd93,-10'd107};
ram[26181] = {9'd96,-10'd104};
ram[26182] = {9'd99,-10'd101};
ram[26183] = {-9'd98,-10'd98};
ram[26184] = {-9'd95,-10'd95};
ram[26185] = {-9'd92,-10'd92};
ram[26186] = {-9'd88,-10'd88};
ram[26187] = {-9'd85,-10'd85};
ram[26188] = {-9'd82,-10'd82};
ram[26189] = {-9'd79,-10'd79};
ram[26190] = {-9'd76,-10'd76};
ram[26191] = {-9'd73,-10'd73};
ram[26192] = {-9'd70,-10'd70};
ram[26193] = {-9'd66,-10'd66};
ram[26194] = {-9'd63,-10'd63};
ram[26195] = {-9'd60,-10'd60};
ram[26196] = {-9'd57,-10'd57};
ram[26197] = {-9'd54,-10'd54};
ram[26198] = {-9'd51,-10'd51};
ram[26199] = {-9'd48,-10'd48};
ram[26200] = {-9'd44,-10'd44};
ram[26201] = {-9'd41,-10'd41};
ram[26202] = {-9'd38,-10'd38};
ram[26203] = {-9'd35,-10'd35};
ram[26204] = {-9'd32,-10'd32};
ram[26205] = {-9'd29,-10'd29};
ram[26206] = {-9'd26,-10'd26};
ram[26207] = {-9'd22,-10'd22};
ram[26208] = {-9'd19,-10'd19};
ram[26209] = {-9'd16,-10'd16};
ram[26210] = {-9'd13,-10'd13};
ram[26211] = {-9'd10,-10'd10};
ram[26212] = {-9'd7,-10'd7};
ram[26213] = {-9'd4,-10'd4};
ram[26214] = {9'd0,10'd0};
ram[26215] = {9'd3,10'd3};
ram[26216] = {9'd6,10'd6};
ram[26217] = {9'd9,10'd9};
ram[26218] = {9'd12,10'd12};
ram[26219] = {9'd15,10'd15};
ram[26220] = {9'd18,10'd18};
ram[26221] = {9'd21,10'd21};
ram[26222] = {9'd25,10'd25};
ram[26223] = {9'd28,10'd28};
ram[26224] = {9'd31,10'd31};
ram[26225] = {9'd34,10'd34};
ram[26226] = {9'd37,10'd37};
ram[26227] = {9'd40,10'd40};
ram[26228] = {9'd43,10'd43};
ram[26229] = {9'd47,10'd47};
ram[26230] = {9'd50,10'd50};
ram[26231] = {9'd53,10'd53};
ram[26232] = {9'd56,10'd56};
ram[26233] = {9'd59,10'd59};
ram[26234] = {9'd62,10'd62};
ram[26235] = {9'd65,10'd65};
ram[26236] = {9'd69,10'd69};
ram[26237] = {9'd72,10'd72};
ram[26238] = {9'd75,10'd75};
ram[26239] = {9'd78,10'd78};
ram[26240] = {9'd78,10'd78};
ram[26241] = {9'd81,10'd81};
ram[26242] = {9'd84,10'd84};
ram[26243] = {9'd87,10'd87};
ram[26244] = {9'd91,10'd91};
ram[26245] = {9'd94,10'd94};
ram[26246] = {9'd97,10'd97};
ram[26247] = {-9'd100,10'd100};
ram[26248] = {-9'd97,10'd103};
ram[26249] = {-9'd94,10'd106};
ram[26250] = {-9'd91,10'd109};
ram[26251] = {-9'd88,10'd113};
ram[26252] = {-9'd85,10'd116};
ram[26253] = {-9'd81,10'd119};
ram[26254] = {-9'd78,10'd122};
ram[26255] = {-9'd75,10'd125};
ram[26256] = {-9'd72,10'd128};
ram[26257] = {-9'd69,10'd131};
ram[26258] = {-9'd66,10'd135};
ram[26259] = {-9'd63,10'd138};
ram[26260] = {-9'd59,10'd141};
ram[26261] = {-9'd56,10'd144};
ram[26262] = {-9'd53,10'd147};
ram[26263] = {-9'd50,10'd150};
ram[26264] = {-9'd47,10'd153};
ram[26265] = {-9'd44,10'd157};
ram[26266] = {-9'd41,10'd160};
ram[26267] = {-9'd37,10'd163};
ram[26268] = {-9'd34,10'd166};
ram[26269] = {-9'd31,10'd169};
ram[26270] = {-9'd28,10'd172};
ram[26271] = {-9'd25,10'd175};
ram[26272] = {-9'd22,10'd179};
ram[26273] = {-9'd19,10'd182};
ram[26274] = {-9'd15,10'd185};
ram[26275] = {-9'd12,10'd188};
ram[26276] = {-9'd9,10'd191};
ram[26277] = {-9'd6,10'd194};
ram[26278] = {-9'd3,10'd197};
ram[26279] = {9'd0,10'd201};
ram[26280] = {9'd3,10'd204};
ram[26281] = {9'd7,10'd207};
ram[26282] = {9'd10,10'd210};
ram[26283] = {9'd13,10'd213};
ram[26284] = {9'd16,10'd216};
ram[26285] = {9'd19,10'd219};
ram[26286] = {9'd22,10'd223};
ram[26287] = {9'd25,10'd226};
ram[26288] = {9'd29,10'd229};
ram[26289] = {9'd32,10'd232};
ram[26290] = {9'd35,10'd235};
ram[26291] = {9'd38,10'd238};
ram[26292] = {9'd41,10'd241};
ram[26293] = {9'd44,10'd245};
ram[26294] = {9'd47,10'd248};
ram[26295] = {9'd51,10'd251};
ram[26296] = {9'd54,10'd254};
ram[26297] = {9'd57,10'd257};
ram[26298] = {9'd60,10'd260};
ram[26299] = {9'd63,10'd263};
ram[26300] = {9'd66,10'd267};
ram[26301] = {9'd69,10'd270};
ram[26302] = {9'd73,10'd273};
ram[26303] = {9'd76,10'd276};
ram[26304] = {9'd79,10'd279};
ram[26305] = {9'd82,10'd282};
ram[26306] = {9'd85,10'd285};
ram[26307] = {9'd88,10'd289};
ram[26308] = {9'd91,10'd292};
ram[26309] = {9'd95,10'd295};
ram[26310] = {9'd98,10'd298};
ram[26311] = {-9'd99,10'd301};
ram[26312] = {-9'd96,10'd304};
ram[26313] = {-9'd93,10'd307};
ram[26314] = {-9'd90,10'd311};
ram[26315] = {-9'd87,10'd314};
ram[26316] = {-9'd84,10'd317};
ram[26317] = {-9'd81,10'd320};
ram[26318] = {-9'd77,10'd323};
ram[26319] = {-9'd74,10'd326};
ram[26320] = {-9'd71,10'd329};
ram[26321] = {-9'd68,10'd333};
ram[26322] = {-9'd65,10'd336};
ram[26323] = {-9'd62,10'd339};
ram[26324] = {-9'd59,10'd342};
ram[26325] = {-9'd55,10'd345};
ram[26326] = {-9'd52,10'd348};
ram[26327] = {-9'd49,10'd351};
ram[26328] = {-9'd46,10'd354};
ram[26329] = {-9'd43,10'd358};
ram[26330] = {-9'd40,10'd361};
ram[26331] = {-9'd37,10'd364};
ram[26332] = {-9'd33,10'd367};
ram[26333] = {-9'd30,10'd370};
ram[26334] = {-9'd27,10'd373};
ram[26335] = {-9'd24,10'd376};
ram[26336] = {-9'd21,10'd380};
ram[26337] = {-9'd18,10'd383};
ram[26338] = {-9'd15,10'd386};
ram[26339] = {-9'd11,10'd389};
ram[26340] = {-9'd8,10'd392};
ram[26341] = {-9'd5,10'd395};
ram[26342] = {-9'd2,10'd398};
ram[26343] = {9'd1,-10'd399};
ram[26344] = {9'd4,-10'd396};
ram[26345] = {9'd7,-10'd393};
ram[26346] = {9'd10,-10'd390};
ram[26347] = {9'd14,-10'd387};
ram[26348] = {9'd17,-10'd384};
ram[26349] = {9'd20,-10'd381};
ram[26350] = {9'd23,-10'd377};
ram[26351] = {9'd26,-10'd374};
ram[26352] = {9'd29,-10'd371};
ram[26353] = {9'd32,-10'd368};
ram[26354] = {9'd36,-10'd365};
ram[26355] = {9'd39,-10'd362};
ram[26356] = {9'd42,-10'd359};
ram[26357] = {9'd45,-10'd355};
ram[26358] = {9'd48,-10'd352};
ram[26359] = {9'd51,-10'd349};
ram[26360] = {9'd54,-10'd346};
ram[26361] = {9'd58,-10'd343};
ram[26362] = {9'd61,-10'd340};
ram[26363] = {9'd64,-10'd337};
ram[26364] = {9'd67,-10'd334};
ram[26365] = {9'd70,-10'd330};
ram[26366] = {9'd73,-10'd327};
ram[26367] = {9'd76,-10'd324};
ram[26368] = {9'd76,-10'd324};
ram[26369] = {9'd80,-10'd321};
ram[26370] = {9'd83,-10'd318};
ram[26371] = {9'd86,-10'd315};
ram[26372] = {9'd89,-10'd312};
ram[26373] = {9'd92,-10'd308};
ram[26374] = {9'd95,-10'd305};
ram[26375] = {9'd98,-10'd302};
ram[26376] = {-9'd99,-10'd299};
ram[26377] = {-9'd96,-10'd296};
ram[26378] = {-9'd92,-10'd293};
ram[26379] = {-9'd89,-10'd290};
ram[26380] = {-9'd86,-10'd286};
ram[26381] = {-9'd83,-10'd283};
ram[26382] = {-9'd80,-10'd280};
ram[26383] = {-9'd77,-10'd277};
ram[26384] = {-9'd74,-10'd274};
ram[26385] = {-9'd70,-10'd271};
ram[26386] = {-9'd67,-10'd268};
ram[26387] = {-9'd64,-10'd264};
ram[26388] = {-9'd61,-10'd261};
ram[26389] = {-9'd58,-10'd258};
ram[26390] = {-9'd55,-10'd255};
ram[26391] = {-9'd52,-10'd252};
ram[26392] = {-9'd48,-10'd249};
ram[26393] = {-9'd45,-10'd246};
ram[26394] = {-9'd42,-10'd242};
ram[26395] = {-9'd39,-10'd239};
ram[26396] = {-9'd36,-10'd236};
ram[26397] = {-9'd33,-10'd233};
ram[26398] = {-9'd30,-10'd230};
ram[26399] = {-9'd26,-10'd227};
ram[26400] = {-9'd23,-10'd224};
ram[26401] = {-9'd20,-10'd220};
ram[26402] = {-9'd17,-10'd217};
ram[26403] = {-9'd14,-10'd214};
ram[26404] = {-9'd11,-10'd211};
ram[26405] = {-9'd8,-10'd208};
ram[26406] = {-9'd4,-10'd205};
ram[26407] = {-9'd1,-10'd202};
ram[26408] = {9'd2,-10'd198};
ram[26409] = {9'd5,-10'd195};
ram[26410] = {9'd8,-10'd192};
ram[26411] = {9'd11,-10'd189};
ram[26412] = {9'd14,-10'd186};
ram[26413] = {9'd18,-10'd183};
ram[26414] = {9'd21,-10'd180};
ram[26415] = {9'd24,-10'd176};
ram[26416] = {9'd27,-10'd173};
ram[26417] = {9'd30,-10'd170};
ram[26418] = {9'd33,-10'd167};
ram[26419] = {9'd36,-10'd164};
ram[26420] = {9'd40,-10'd161};
ram[26421] = {9'd43,-10'd158};
ram[26422] = {9'd46,-10'd154};
ram[26423] = {9'd49,-10'd151};
ram[26424] = {9'd52,-10'd148};
ram[26425] = {9'd55,-10'd145};
ram[26426] = {9'd58,-10'd142};
ram[26427] = {9'd62,-10'd139};
ram[26428] = {9'd65,-10'd136};
ram[26429] = {9'd68,-10'd132};
ram[26430] = {9'd71,-10'd129};
ram[26431] = {9'd74,-10'd126};
ram[26432] = {9'd77,-10'd123};
ram[26433] = {9'd80,-10'd120};
ram[26434] = {9'd84,-10'd117};
ram[26435] = {9'd87,-10'd114};
ram[26436] = {9'd90,-10'd110};
ram[26437] = {9'd93,-10'd107};
ram[26438] = {9'd96,-10'd104};
ram[26439] = {9'd99,-10'd101};
ram[26440] = {-9'd98,-10'd98};
ram[26441] = {-9'd95,-10'd95};
ram[26442] = {-9'd92,-10'd92};
ram[26443] = {-9'd88,-10'd88};
ram[26444] = {-9'd85,-10'd85};
ram[26445] = {-9'd82,-10'd82};
ram[26446] = {-9'd79,-10'd79};
ram[26447] = {-9'd76,-10'd76};
ram[26448] = {-9'd73,-10'd73};
ram[26449] = {-9'd70,-10'd70};
ram[26450] = {-9'd66,-10'd66};
ram[26451] = {-9'd63,-10'd63};
ram[26452] = {-9'd60,-10'd60};
ram[26453] = {-9'd57,-10'd57};
ram[26454] = {-9'd54,-10'd54};
ram[26455] = {-9'd51,-10'd51};
ram[26456] = {-9'd48,-10'd48};
ram[26457] = {-9'd44,-10'd44};
ram[26458] = {-9'd41,-10'd41};
ram[26459] = {-9'd38,-10'd38};
ram[26460] = {-9'd35,-10'd35};
ram[26461] = {-9'd32,-10'd32};
ram[26462] = {-9'd29,-10'd29};
ram[26463] = {-9'd26,-10'd26};
ram[26464] = {-9'd22,-10'd22};
ram[26465] = {-9'd19,-10'd19};
ram[26466] = {-9'd16,-10'd16};
ram[26467] = {-9'd13,-10'd13};
ram[26468] = {-9'd10,-10'd10};
ram[26469] = {-9'd7,-10'd7};
ram[26470] = {-9'd4,-10'd4};
ram[26471] = {9'd0,10'd0};
ram[26472] = {9'd3,10'd3};
ram[26473] = {9'd6,10'd6};
ram[26474] = {9'd9,10'd9};
ram[26475] = {9'd12,10'd12};
ram[26476] = {9'd15,10'd15};
ram[26477] = {9'd18,10'd18};
ram[26478] = {9'd21,10'd21};
ram[26479] = {9'd25,10'd25};
ram[26480] = {9'd28,10'd28};
ram[26481] = {9'd31,10'd31};
ram[26482] = {9'd34,10'd34};
ram[26483] = {9'd37,10'd37};
ram[26484] = {9'd40,10'd40};
ram[26485] = {9'd43,10'd43};
ram[26486] = {9'd47,10'd47};
ram[26487] = {9'd50,10'd50};
ram[26488] = {9'd53,10'd53};
ram[26489] = {9'd56,10'd56};
ram[26490] = {9'd59,10'd59};
ram[26491] = {9'd62,10'd62};
ram[26492] = {9'd65,10'd65};
ram[26493] = {9'd69,10'd69};
ram[26494] = {9'd72,10'd72};
ram[26495] = {9'd75,10'd75};
ram[26496] = {9'd75,10'd75};
ram[26497] = {9'd78,10'd78};
ram[26498] = {9'd81,10'd81};
ram[26499] = {9'd84,10'd84};
ram[26500] = {9'd87,10'd87};
ram[26501] = {9'd91,10'd91};
ram[26502] = {9'd94,10'd94};
ram[26503] = {9'd97,10'd97};
ram[26504] = {-9'd100,10'd100};
ram[26505] = {-9'd97,10'd103};
ram[26506] = {-9'd94,10'd106};
ram[26507] = {-9'd91,10'd109};
ram[26508] = {-9'd88,10'd113};
ram[26509] = {-9'd85,10'd116};
ram[26510] = {-9'd81,10'd119};
ram[26511] = {-9'd78,10'd122};
ram[26512] = {-9'd75,10'd125};
ram[26513] = {-9'd72,10'd128};
ram[26514] = {-9'd69,10'd131};
ram[26515] = {-9'd66,10'd135};
ram[26516] = {-9'd63,10'd138};
ram[26517] = {-9'd59,10'd141};
ram[26518] = {-9'd56,10'd144};
ram[26519] = {-9'd53,10'd147};
ram[26520] = {-9'd50,10'd150};
ram[26521] = {-9'd47,10'd153};
ram[26522] = {-9'd44,10'd157};
ram[26523] = {-9'd41,10'd160};
ram[26524] = {-9'd37,10'd163};
ram[26525] = {-9'd34,10'd166};
ram[26526] = {-9'd31,10'd169};
ram[26527] = {-9'd28,10'd172};
ram[26528] = {-9'd25,10'd175};
ram[26529] = {-9'd22,10'd179};
ram[26530] = {-9'd19,10'd182};
ram[26531] = {-9'd15,10'd185};
ram[26532] = {-9'd12,10'd188};
ram[26533] = {-9'd9,10'd191};
ram[26534] = {-9'd6,10'd194};
ram[26535] = {-9'd3,10'd197};
ram[26536] = {9'd0,10'd201};
ram[26537] = {9'd3,10'd204};
ram[26538] = {9'd7,10'd207};
ram[26539] = {9'd10,10'd210};
ram[26540] = {9'd13,10'd213};
ram[26541] = {9'd16,10'd216};
ram[26542] = {9'd19,10'd219};
ram[26543] = {9'd22,10'd223};
ram[26544] = {9'd25,10'd226};
ram[26545] = {9'd29,10'd229};
ram[26546] = {9'd32,10'd232};
ram[26547] = {9'd35,10'd235};
ram[26548] = {9'd38,10'd238};
ram[26549] = {9'd41,10'd241};
ram[26550] = {9'd44,10'd245};
ram[26551] = {9'd47,10'd248};
ram[26552] = {9'd51,10'd251};
ram[26553] = {9'd54,10'd254};
ram[26554] = {9'd57,10'd257};
ram[26555] = {9'd60,10'd260};
ram[26556] = {9'd63,10'd263};
ram[26557] = {9'd66,10'd267};
ram[26558] = {9'd69,10'd270};
ram[26559] = {9'd73,10'd273};
ram[26560] = {9'd76,10'd276};
ram[26561] = {9'd79,10'd279};
ram[26562] = {9'd82,10'd282};
ram[26563] = {9'd85,10'd285};
ram[26564] = {9'd88,10'd289};
ram[26565] = {9'd91,10'd292};
ram[26566] = {9'd95,10'd295};
ram[26567] = {9'd98,10'd298};
ram[26568] = {-9'd99,10'd301};
ram[26569] = {-9'd96,10'd304};
ram[26570] = {-9'd93,10'd307};
ram[26571] = {-9'd90,10'd311};
ram[26572] = {-9'd87,10'd314};
ram[26573] = {-9'd84,10'd317};
ram[26574] = {-9'd81,10'd320};
ram[26575] = {-9'd77,10'd323};
ram[26576] = {-9'd74,10'd326};
ram[26577] = {-9'd71,10'd329};
ram[26578] = {-9'd68,10'd333};
ram[26579] = {-9'd65,10'd336};
ram[26580] = {-9'd62,10'd339};
ram[26581] = {-9'd59,10'd342};
ram[26582] = {-9'd55,10'd345};
ram[26583] = {-9'd52,10'd348};
ram[26584] = {-9'd49,10'd351};
ram[26585] = {-9'd46,10'd354};
ram[26586] = {-9'd43,10'd358};
ram[26587] = {-9'd40,10'd361};
ram[26588] = {-9'd37,10'd364};
ram[26589] = {-9'd33,10'd367};
ram[26590] = {-9'd30,10'd370};
ram[26591] = {-9'd27,10'd373};
ram[26592] = {-9'd24,10'd376};
ram[26593] = {-9'd21,10'd380};
ram[26594] = {-9'd18,10'd383};
ram[26595] = {-9'd15,10'd386};
ram[26596] = {-9'd11,10'd389};
ram[26597] = {-9'd8,10'd392};
ram[26598] = {-9'd5,10'd395};
ram[26599] = {-9'd2,10'd398};
ram[26600] = {9'd1,-10'd399};
ram[26601] = {9'd4,-10'd396};
ram[26602] = {9'd7,-10'd393};
ram[26603] = {9'd10,-10'd390};
ram[26604] = {9'd14,-10'd387};
ram[26605] = {9'd17,-10'd384};
ram[26606] = {9'd20,-10'd381};
ram[26607] = {9'd23,-10'd377};
ram[26608] = {9'd26,-10'd374};
ram[26609] = {9'd29,-10'd371};
ram[26610] = {9'd32,-10'd368};
ram[26611] = {9'd36,-10'd365};
ram[26612] = {9'd39,-10'd362};
ram[26613] = {9'd42,-10'd359};
ram[26614] = {9'd45,-10'd355};
ram[26615] = {9'd48,-10'd352};
ram[26616] = {9'd51,-10'd349};
ram[26617] = {9'd54,-10'd346};
ram[26618] = {9'd58,-10'd343};
ram[26619] = {9'd61,-10'd340};
ram[26620] = {9'd64,-10'd337};
ram[26621] = {9'd67,-10'd334};
ram[26622] = {9'd70,-10'd330};
ram[26623] = {9'd73,-10'd327};
ram[26624] = {9'd73,-10'd327};
ram[26625] = {9'd76,-10'd324};
ram[26626] = {9'd80,-10'd321};
ram[26627] = {9'd83,-10'd318};
ram[26628] = {9'd86,-10'd315};
ram[26629] = {9'd89,-10'd312};
ram[26630] = {9'd92,-10'd308};
ram[26631] = {9'd95,-10'd305};
ram[26632] = {9'd98,-10'd302};
ram[26633] = {-9'd99,-10'd299};
ram[26634] = {-9'd96,-10'd296};
ram[26635] = {-9'd92,-10'd293};
ram[26636] = {-9'd89,-10'd290};
ram[26637] = {-9'd86,-10'd286};
ram[26638] = {-9'd83,-10'd283};
ram[26639] = {-9'd80,-10'd280};
ram[26640] = {-9'd77,-10'd277};
ram[26641] = {-9'd74,-10'd274};
ram[26642] = {-9'd70,-10'd271};
ram[26643] = {-9'd67,-10'd268};
ram[26644] = {-9'd64,-10'd264};
ram[26645] = {-9'd61,-10'd261};
ram[26646] = {-9'd58,-10'd258};
ram[26647] = {-9'd55,-10'd255};
ram[26648] = {-9'd52,-10'd252};
ram[26649] = {-9'd48,-10'd249};
ram[26650] = {-9'd45,-10'd246};
ram[26651] = {-9'd42,-10'd242};
ram[26652] = {-9'd39,-10'd239};
ram[26653] = {-9'd36,-10'd236};
ram[26654] = {-9'd33,-10'd233};
ram[26655] = {-9'd30,-10'd230};
ram[26656] = {-9'd26,-10'd227};
ram[26657] = {-9'd23,-10'd224};
ram[26658] = {-9'd20,-10'd220};
ram[26659] = {-9'd17,-10'd217};
ram[26660] = {-9'd14,-10'd214};
ram[26661] = {-9'd11,-10'd211};
ram[26662] = {-9'd8,-10'd208};
ram[26663] = {-9'd4,-10'd205};
ram[26664] = {-9'd1,-10'd202};
ram[26665] = {9'd2,-10'd198};
ram[26666] = {9'd5,-10'd195};
ram[26667] = {9'd8,-10'd192};
ram[26668] = {9'd11,-10'd189};
ram[26669] = {9'd14,-10'd186};
ram[26670] = {9'd18,-10'd183};
ram[26671] = {9'd21,-10'd180};
ram[26672] = {9'd24,-10'd176};
ram[26673] = {9'd27,-10'd173};
ram[26674] = {9'd30,-10'd170};
ram[26675] = {9'd33,-10'd167};
ram[26676] = {9'd36,-10'd164};
ram[26677] = {9'd40,-10'd161};
ram[26678] = {9'd43,-10'd158};
ram[26679] = {9'd46,-10'd154};
ram[26680] = {9'd49,-10'd151};
ram[26681] = {9'd52,-10'd148};
ram[26682] = {9'd55,-10'd145};
ram[26683] = {9'd58,-10'd142};
ram[26684] = {9'd62,-10'd139};
ram[26685] = {9'd65,-10'd136};
ram[26686] = {9'd68,-10'd132};
ram[26687] = {9'd71,-10'd129};
ram[26688] = {9'd74,-10'd126};
ram[26689] = {9'd77,-10'd123};
ram[26690] = {9'd80,-10'd120};
ram[26691] = {9'd84,-10'd117};
ram[26692] = {9'd87,-10'd114};
ram[26693] = {9'd90,-10'd110};
ram[26694] = {9'd93,-10'd107};
ram[26695] = {9'd96,-10'd104};
ram[26696] = {9'd99,-10'd101};
ram[26697] = {-9'd98,-10'd98};
ram[26698] = {-9'd95,-10'd95};
ram[26699] = {-9'd92,-10'd92};
ram[26700] = {-9'd88,-10'd88};
ram[26701] = {-9'd85,-10'd85};
ram[26702] = {-9'd82,-10'd82};
ram[26703] = {-9'd79,-10'd79};
ram[26704] = {-9'd76,-10'd76};
ram[26705] = {-9'd73,-10'd73};
ram[26706] = {-9'd70,-10'd70};
ram[26707] = {-9'd66,-10'd66};
ram[26708] = {-9'd63,-10'd63};
ram[26709] = {-9'd60,-10'd60};
ram[26710] = {-9'd57,-10'd57};
ram[26711] = {-9'd54,-10'd54};
ram[26712] = {-9'd51,-10'd51};
ram[26713] = {-9'd48,-10'd48};
ram[26714] = {-9'd44,-10'd44};
ram[26715] = {-9'd41,-10'd41};
ram[26716] = {-9'd38,-10'd38};
ram[26717] = {-9'd35,-10'd35};
ram[26718] = {-9'd32,-10'd32};
ram[26719] = {-9'd29,-10'd29};
ram[26720] = {-9'd26,-10'd26};
ram[26721] = {-9'd22,-10'd22};
ram[26722] = {-9'd19,-10'd19};
ram[26723] = {-9'd16,-10'd16};
ram[26724] = {-9'd13,-10'd13};
ram[26725] = {-9'd10,-10'd10};
ram[26726] = {-9'd7,-10'd7};
ram[26727] = {-9'd4,-10'd4};
ram[26728] = {9'd0,10'd0};
ram[26729] = {9'd3,10'd3};
ram[26730] = {9'd6,10'd6};
ram[26731] = {9'd9,10'd9};
ram[26732] = {9'd12,10'd12};
ram[26733] = {9'd15,10'd15};
ram[26734] = {9'd18,10'd18};
ram[26735] = {9'd21,10'd21};
ram[26736] = {9'd25,10'd25};
ram[26737] = {9'd28,10'd28};
ram[26738] = {9'd31,10'd31};
ram[26739] = {9'd34,10'd34};
ram[26740] = {9'd37,10'd37};
ram[26741] = {9'd40,10'd40};
ram[26742] = {9'd43,10'd43};
ram[26743] = {9'd47,10'd47};
ram[26744] = {9'd50,10'd50};
ram[26745] = {9'd53,10'd53};
ram[26746] = {9'd56,10'd56};
ram[26747] = {9'd59,10'd59};
ram[26748] = {9'd62,10'd62};
ram[26749] = {9'd65,10'd65};
ram[26750] = {9'd69,10'd69};
ram[26751] = {9'd72,10'd72};
ram[26752] = {9'd72,10'd72};
ram[26753] = {9'd75,10'd75};
ram[26754] = {9'd78,10'd78};
ram[26755] = {9'd81,10'd81};
ram[26756] = {9'd84,10'd84};
ram[26757] = {9'd87,10'd87};
ram[26758] = {9'd91,10'd91};
ram[26759] = {9'd94,10'd94};
ram[26760] = {9'd97,10'd97};
ram[26761] = {-9'd100,10'd100};
ram[26762] = {-9'd97,10'd103};
ram[26763] = {-9'd94,10'd106};
ram[26764] = {-9'd91,10'd109};
ram[26765] = {-9'd88,10'd113};
ram[26766] = {-9'd85,10'd116};
ram[26767] = {-9'd81,10'd119};
ram[26768] = {-9'd78,10'd122};
ram[26769] = {-9'd75,10'd125};
ram[26770] = {-9'd72,10'd128};
ram[26771] = {-9'd69,10'd131};
ram[26772] = {-9'd66,10'd135};
ram[26773] = {-9'd63,10'd138};
ram[26774] = {-9'd59,10'd141};
ram[26775] = {-9'd56,10'd144};
ram[26776] = {-9'd53,10'd147};
ram[26777] = {-9'd50,10'd150};
ram[26778] = {-9'd47,10'd153};
ram[26779] = {-9'd44,10'd157};
ram[26780] = {-9'd41,10'd160};
ram[26781] = {-9'd37,10'd163};
ram[26782] = {-9'd34,10'd166};
ram[26783] = {-9'd31,10'd169};
ram[26784] = {-9'd28,10'd172};
ram[26785] = {-9'd25,10'd175};
ram[26786] = {-9'd22,10'd179};
ram[26787] = {-9'd19,10'd182};
ram[26788] = {-9'd15,10'd185};
ram[26789] = {-9'd12,10'd188};
ram[26790] = {-9'd9,10'd191};
ram[26791] = {-9'd6,10'd194};
ram[26792] = {-9'd3,10'd197};
ram[26793] = {9'd0,10'd201};
ram[26794] = {9'd3,10'd204};
ram[26795] = {9'd7,10'd207};
ram[26796] = {9'd10,10'd210};
ram[26797] = {9'd13,10'd213};
ram[26798] = {9'd16,10'd216};
ram[26799] = {9'd19,10'd219};
ram[26800] = {9'd22,10'd223};
ram[26801] = {9'd25,10'd226};
ram[26802] = {9'd29,10'd229};
ram[26803] = {9'd32,10'd232};
ram[26804] = {9'd35,10'd235};
ram[26805] = {9'd38,10'd238};
ram[26806] = {9'd41,10'd241};
ram[26807] = {9'd44,10'd245};
ram[26808] = {9'd47,10'd248};
ram[26809] = {9'd51,10'd251};
ram[26810] = {9'd54,10'd254};
ram[26811] = {9'd57,10'd257};
ram[26812] = {9'd60,10'd260};
ram[26813] = {9'd63,10'd263};
ram[26814] = {9'd66,10'd267};
ram[26815] = {9'd69,10'd270};
ram[26816] = {9'd73,10'd273};
ram[26817] = {9'd76,10'd276};
ram[26818] = {9'd79,10'd279};
ram[26819] = {9'd82,10'd282};
ram[26820] = {9'd85,10'd285};
ram[26821] = {9'd88,10'd289};
ram[26822] = {9'd91,10'd292};
ram[26823] = {9'd95,10'd295};
ram[26824] = {9'd98,10'd298};
ram[26825] = {-9'd99,10'd301};
ram[26826] = {-9'd96,10'd304};
ram[26827] = {-9'd93,10'd307};
ram[26828] = {-9'd90,10'd311};
ram[26829] = {-9'd87,10'd314};
ram[26830] = {-9'd84,10'd317};
ram[26831] = {-9'd81,10'd320};
ram[26832] = {-9'd77,10'd323};
ram[26833] = {-9'd74,10'd326};
ram[26834] = {-9'd71,10'd329};
ram[26835] = {-9'd68,10'd333};
ram[26836] = {-9'd65,10'd336};
ram[26837] = {-9'd62,10'd339};
ram[26838] = {-9'd59,10'd342};
ram[26839] = {-9'd55,10'd345};
ram[26840] = {-9'd52,10'd348};
ram[26841] = {-9'd49,10'd351};
ram[26842] = {-9'd46,10'd354};
ram[26843] = {-9'd43,10'd358};
ram[26844] = {-9'd40,10'd361};
ram[26845] = {-9'd37,10'd364};
ram[26846] = {-9'd33,10'd367};
ram[26847] = {-9'd30,10'd370};
ram[26848] = {-9'd27,10'd373};
ram[26849] = {-9'd24,10'd376};
ram[26850] = {-9'd21,10'd380};
ram[26851] = {-9'd18,10'd383};
ram[26852] = {-9'd15,10'd386};
ram[26853] = {-9'd11,10'd389};
ram[26854] = {-9'd8,10'd392};
ram[26855] = {-9'd5,10'd395};
ram[26856] = {-9'd2,10'd398};
ram[26857] = {9'd1,-10'd399};
ram[26858] = {9'd4,-10'd396};
ram[26859] = {9'd7,-10'd393};
ram[26860] = {9'd10,-10'd390};
ram[26861] = {9'd14,-10'd387};
ram[26862] = {9'd17,-10'd384};
ram[26863] = {9'd20,-10'd381};
ram[26864] = {9'd23,-10'd377};
ram[26865] = {9'd26,-10'd374};
ram[26866] = {9'd29,-10'd371};
ram[26867] = {9'd32,-10'd368};
ram[26868] = {9'd36,-10'd365};
ram[26869] = {9'd39,-10'd362};
ram[26870] = {9'd42,-10'd359};
ram[26871] = {9'd45,-10'd355};
ram[26872] = {9'd48,-10'd352};
ram[26873] = {9'd51,-10'd349};
ram[26874] = {9'd54,-10'd346};
ram[26875] = {9'd58,-10'd343};
ram[26876] = {9'd61,-10'd340};
ram[26877] = {9'd64,-10'd337};
ram[26878] = {9'd67,-10'd334};
ram[26879] = {9'd70,-10'd330};
ram[26880] = {9'd70,-10'd330};
ram[26881] = {9'd73,-10'd327};
ram[26882] = {9'd76,-10'd324};
ram[26883] = {9'd80,-10'd321};
ram[26884] = {9'd83,-10'd318};
ram[26885] = {9'd86,-10'd315};
ram[26886] = {9'd89,-10'd312};
ram[26887] = {9'd92,-10'd308};
ram[26888] = {9'd95,-10'd305};
ram[26889] = {9'd98,-10'd302};
ram[26890] = {-9'd99,-10'd299};
ram[26891] = {-9'd96,-10'd296};
ram[26892] = {-9'd92,-10'd293};
ram[26893] = {-9'd89,-10'd290};
ram[26894] = {-9'd86,-10'd286};
ram[26895] = {-9'd83,-10'd283};
ram[26896] = {-9'd80,-10'd280};
ram[26897] = {-9'd77,-10'd277};
ram[26898] = {-9'd74,-10'd274};
ram[26899] = {-9'd70,-10'd271};
ram[26900] = {-9'd67,-10'd268};
ram[26901] = {-9'd64,-10'd264};
ram[26902] = {-9'd61,-10'd261};
ram[26903] = {-9'd58,-10'd258};
ram[26904] = {-9'd55,-10'd255};
ram[26905] = {-9'd52,-10'd252};
ram[26906] = {-9'd48,-10'd249};
ram[26907] = {-9'd45,-10'd246};
ram[26908] = {-9'd42,-10'd242};
ram[26909] = {-9'd39,-10'd239};
ram[26910] = {-9'd36,-10'd236};
ram[26911] = {-9'd33,-10'd233};
ram[26912] = {-9'd30,-10'd230};
ram[26913] = {-9'd26,-10'd227};
ram[26914] = {-9'd23,-10'd224};
ram[26915] = {-9'd20,-10'd220};
ram[26916] = {-9'd17,-10'd217};
ram[26917] = {-9'd14,-10'd214};
ram[26918] = {-9'd11,-10'd211};
ram[26919] = {-9'd8,-10'd208};
ram[26920] = {-9'd4,-10'd205};
ram[26921] = {-9'd1,-10'd202};
ram[26922] = {9'd2,-10'd198};
ram[26923] = {9'd5,-10'd195};
ram[26924] = {9'd8,-10'd192};
ram[26925] = {9'd11,-10'd189};
ram[26926] = {9'd14,-10'd186};
ram[26927] = {9'd18,-10'd183};
ram[26928] = {9'd21,-10'd180};
ram[26929] = {9'd24,-10'd176};
ram[26930] = {9'd27,-10'd173};
ram[26931] = {9'd30,-10'd170};
ram[26932] = {9'd33,-10'd167};
ram[26933] = {9'd36,-10'd164};
ram[26934] = {9'd40,-10'd161};
ram[26935] = {9'd43,-10'd158};
ram[26936] = {9'd46,-10'd154};
ram[26937] = {9'd49,-10'd151};
ram[26938] = {9'd52,-10'd148};
ram[26939] = {9'd55,-10'd145};
ram[26940] = {9'd58,-10'd142};
ram[26941] = {9'd62,-10'd139};
ram[26942] = {9'd65,-10'd136};
ram[26943] = {9'd68,-10'd132};
ram[26944] = {9'd71,-10'd129};
ram[26945] = {9'd74,-10'd126};
ram[26946] = {9'd77,-10'd123};
ram[26947] = {9'd80,-10'd120};
ram[26948] = {9'd84,-10'd117};
ram[26949] = {9'd87,-10'd114};
ram[26950] = {9'd90,-10'd110};
ram[26951] = {9'd93,-10'd107};
ram[26952] = {9'd96,-10'd104};
ram[26953] = {9'd99,-10'd101};
ram[26954] = {-9'd98,-10'd98};
ram[26955] = {-9'd95,-10'd95};
ram[26956] = {-9'd92,-10'd92};
ram[26957] = {-9'd88,-10'd88};
ram[26958] = {-9'd85,-10'd85};
ram[26959] = {-9'd82,-10'd82};
ram[26960] = {-9'd79,-10'd79};
ram[26961] = {-9'd76,-10'd76};
ram[26962] = {-9'd73,-10'd73};
ram[26963] = {-9'd70,-10'd70};
ram[26964] = {-9'd66,-10'd66};
ram[26965] = {-9'd63,-10'd63};
ram[26966] = {-9'd60,-10'd60};
ram[26967] = {-9'd57,-10'd57};
ram[26968] = {-9'd54,-10'd54};
ram[26969] = {-9'd51,-10'd51};
ram[26970] = {-9'd48,-10'd48};
ram[26971] = {-9'd44,-10'd44};
ram[26972] = {-9'd41,-10'd41};
ram[26973] = {-9'd38,-10'd38};
ram[26974] = {-9'd35,-10'd35};
ram[26975] = {-9'd32,-10'd32};
ram[26976] = {-9'd29,-10'd29};
ram[26977] = {-9'd26,-10'd26};
ram[26978] = {-9'd22,-10'd22};
ram[26979] = {-9'd19,-10'd19};
ram[26980] = {-9'd16,-10'd16};
ram[26981] = {-9'd13,-10'd13};
ram[26982] = {-9'd10,-10'd10};
ram[26983] = {-9'd7,-10'd7};
ram[26984] = {-9'd4,-10'd4};
ram[26985] = {9'd0,10'd0};
ram[26986] = {9'd3,10'd3};
ram[26987] = {9'd6,10'd6};
ram[26988] = {9'd9,10'd9};
ram[26989] = {9'd12,10'd12};
ram[26990] = {9'd15,10'd15};
ram[26991] = {9'd18,10'd18};
ram[26992] = {9'd21,10'd21};
ram[26993] = {9'd25,10'd25};
ram[26994] = {9'd28,10'd28};
ram[26995] = {9'd31,10'd31};
ram[26996] = {9'd34,10'd34};
ram[26997] = {9'd37,10'd37};
ram[26998] = {9'd40,10'd40};
ram[26999] = {9'd43,10'd43};
ram[27000] = {9'd47,10'd47};
ram[27001] = {9'd50,10'd50};
ram[27002] = {9'd53,10'd53};
ram[27003] = {9'd56,10'd56};
ram[27004] = {9'd59,10'd59};
ram[27005] = {9'd62,10'd62};
ram[27006] = {9'd65,10'd65};
ram[27007] = {9'd69,10'd69};
ram[27008] = {9'd69,10'd69};
ram[27009] = {9'd72,10'd72};
ram[27010] = {9'd75,10'd75};
ram[27011] = {9'd78,10'd78};
ram[27012] = {9'd81,10'd81};
ram[27013] = {9'd84,10'd84};
ram[27014] = {9'd87,10'd87};
ram[27015] = {9'd91,10'd91};
ram[27016] = {9'd94,10'd94};
ram[27017] = {9'd97,10'd97};
ram[27018] = {-9'd100,10'd100};
ram[27019] = {-9'd97,10'd103};
ram[27020] = {-9'd94,10'd106};
ram[27021] = {-9'd91,10'd109};
ram[27022] = {-9'd88,10'd113};
ram[27023] = {-9'd85,10'd116};
ram[27024] = {-9'd81,10'd119};
ram[27025] = {-9'd78,10'd122};
ram[27026] = {-9'd75,10'd125};
ram[27027] = {-9'd72,10'd128};
ram[27028] = {-9'd69,10'd131};
ram[27029] = {-9'd66,10'd135};
ram[27030] = {-9'd63,10'd138};
ram[27031] = {-9'd59,10'd141};
ram[27032] = {-9'd56,10'd144};
ram[27033] = {-9'd53,10'd147};
ram[27034] = {-9'd50,10'd150};
ram[27035] = {-9'd47,10'd153};
ram[27036] = {-9'd44,10'd157};
ram[27037] = {-9'd41,10'd160};
ram[27038] = {-9'd37,10'd163};
ram[27039] = {-9'd34,10'd166};
ram[27040] = {-9'd31,10'd169};
ram[27041] = {-9'd28,10'd172};
ram[27042] = {-9'd25,10'd175};
ram[27043] = {-9'd22,10'd179};
ram[27044] = {-9'd19,10'd182};
ram[27045] = {-9'd15,10'd185};
ram[27046] = {-9'd12,10'd188};
ram[27047] = {-9'd9,10'd191};
ram[27048] = {-9'd6,10'd194};
ram[27049] = {-9'd3,10'd197};
ram[27050] = {9'd0,10'd201};
ram[27051] = {9'd3,10'd204};
ram[27052] = {9'd7,10'd207};
ram[27053] = {9'd10,10'd210};
ram[27054] = {9'd13,10'd213};
ram[27055] = {9'd16,10'd216};
ram[27056] = {9'd19,10'd219};
ram[27057] = {9'd22,10'd223};
ram[27058] = {9'd25,10'd226};
ram[27059] = {9'd29,10'd229};
ram[27060] = {9'd32,10'd232};
ram[27061] = {9'd35,10'd235};
ram[27062] = {9'd38,10'd238};
ram[27063] = {9'd41,10'd241};
ram[27064] = {9'd44,10'd245};
ram[27065] = {9'd47,10'd248};
ram[27066] = {9'd51,10'd251};
ram[27067] = {9'd54,10'd254};
ram[27068] = {9'd57,10'd257};
ram[27069] = {9'd60,10'd260};
ram[27070] = {9'd63,10'd263};
ram[27071] = {9'd66,10'd267};
ram[27072] = {9'd69,10'd270};
ram[27073] = {9'd73,10'd273};
ram[27074] = {9'd76,10'd276};
ram[27075] = {9'd79,10'd279};
ram[27076] = {9'd82,10'd282};
ram[27077] = {9'd85,10'd285};
ram[27078] = {9'd88,10'd289};
ram[27079] = {9'd91,10'd292};
ram[27080] = {9'd95,10'd295};
ram[27081] = {9'd98,10'd298};
ram[27082] = {-9'd99,10'd301};
ram[27083] = {-9'd96,10'd304};
ram[27084] = {-9'd93,10'd307};
ram[27085] = {-9'd90,10'd311};
ram[27086] = {-9'd87,10'd314};
ram[27087] = {-9'd84,10'd317};
ram[27088] = {-9'd81,10'd320};
ram[27089] = {-9'd77,10'd323};
ram[27090] = {-9'd74,10'd326};
ram[27091] = {-9'd71,10'd329};
ram[27092] = {-9'd68,10'd333};
ram[27093] = {-9'd65,10'd336};
ram[27094] = {-9'd62,10'd339};
ram[27095] = {-9'd59,10'd342};
ram[27096] = {-9'd55,10'd345};
ram[27097] = {-9'd52,10'd348};
ram[27098] = {-9'd49,10'd351};
ram[27099] = {-9'd46,10'd354};
ram[27100] = {-9'd43,10'd358};
ram[27101] = {-9'd40,10'd361};
ram[27102] = {-9'd37,10'd364};
ram[27103] = {-9'd33,10'd367};
ram[27104] = {-9'd30,10'd370};
ram[27105] = {-9'd27,10'd373};
ram[27106] = {-9'd24,10'd376};
ram[27107] = {-9'd21,10'd380};
ram[27108] = {-9'd18,10'd383};
ram[27109] = {-9'd15,10'd386};
ram[27110] = {-9'd11,10'd389};
ram[27111] = {-9'd8,10'd392};
ram[27112] = {-9'd5,10'd395};
ram[27113] = {-9'd2,10'd398};
ram[27114] = {9'd1,-10'd399};
ram[27115] = {9'd4,-10'd396};
ram[27116] = {9'd7,-10'd393};
ram[27117] = {9'd10,-10'd390};
ram[27118] = {9'd14,-10'd387};
ram[27119] = {9'd17,-10'd384};
ram[27120] = {9'd20,-10'd381};
ram[27121] = {9'd23,-10'd377};
ram[27122] = {9'd26,-10'd374};
ram[27123] = {9'd29,-10'd371};
ram[27124] = {9'd32,-10'd368};
ram[27125] = {9'd36,-10'd365};
ram[27126] = {9'd39,-10'd362};
ram[27127] = {9'd42,-10'd359};
ram[27128] = {9'd45,-10'd355};
ram[27129] = {9'd48,-10'd352};
ram[27130] = {9'd51,-10'd349};
ram[27131] = {9'd54,-10'd346};
ram[27132] = {9'd58,-10'd343};
ram[27133] = {9'd61,-10'd340};
ram[27134] = {9'd64,-10'd337};
ram[27135] = {9'd67,-10'd334};
ram[27136] = {9'd67,-10'd334};
ram[27137] = {9'd70,-10'd330};
ram[27138] = {9'd73,-10'd327};
ram[27139] = {9'd76,-10'd324};
ram[27140] = {9'd80,-10'd321};
ram[27141] = {9'd83,-10'd318};
ram[27142] = {9'd86,-10'd315};
ram[27143] = {9'd89,-10'd312};
ram[27144] = {9'd92,-10'd308};
ram[27145] = {9'd95,-10'd305};
ram[27146] = {9'd98,-10'd302};
ram[27147] = {-9'd99,-10'd299};
ram[27148] = {-9'd96,-10'd296};
ram[27149] = {-9'd92,-10'd293};
ram[27150] = {-9'd89,-10'd290};
ram[27151] = {-9'd86,-10'd286};
ram[27152] = {-9'd83,-10'd283};
ram[27153] = {-9'd80,-10'd280};
ram[27154] = {-9'd77,-10'd277};
ram[27155] = {-9'd74,-10'd274};
ram[27156] = {-9'd70,-10'd271};
ram[27157] = {-9'd67,-10'd268};
ram[27158] = {-9'd64,-10'd264};
ram[27159] = {-9'd61,-10'd261};
ram[27160] = {-9'd58,-10'd258};
ram[27161] = {-9'd55,-10'd255};
ram[27162] = {-9'd52,-10'd252};
ram[27163] = {-9'd48,-10'd249};
ram[27164] = {-9'd45,-10'd246};
ram[27165] = {-9'd42,-10'd242};
ram[27166] = {-9'd39,-10'd239};
ram[27167] = {-9'd36,-10'd236};
ram[27168] = {-9'd33,-10'd233};
ram[27169] = {-9'd30,-10'd230};
ram[27170] = {-9'd26,-10'd227};
ram[27171] = {-9'd23,-10'd224};
ram[27172] = {-9'd20,-10'd220};
ram[27173] = {-9'd17,-10'd217};
ram[27174] = {-9'd14,-10'd214};
ram[27175] = {-9'd11,-10'd211};
ram[27176] = {-9'd8,-10'd208};
ram[27177] = {-9'd4,-10'd205};
ram[27178] = {-9'd1,-10'd202};
ram[27179] = {9'd2,-10'd198};
ram[27180] = {9'd5,-10'd195};
ram[27181] = {9'd8,-10'd192};
ram[27182] = {9'd11,-10'd189};
ram[27183] = {9'd14,-10'd186};
ram[27184] = {9'd18,-10'd183};
ram[27185] = {9'd21,-10'd180};
ram[27186] = {9'd24,-10'd176};
ram[27187] = {9'd27,-10'd173};
ram[27188] = {9'd30,-10'd170};
ram[27189] = {9'd33,-10'd167};
ram[27190] = {9'd36,-10'd164};
ram[27191] = {9'd40,-10'd161};
ram[27192] = {9'd43,-10'd158};
ram[27193] = {9'd46,-10'd154};
ram[27194] = {9'd49,-10'd151};
ram[27195] = {9'd52,-10'd148};
ram[27196] = {9'd55,-10'd145};
ram[27197] = {9'd58,-10'd142};
ram[27198] = {9'd62,-10'd139};
ram[27199] = {9'd65,-10'd136};
ram[27200] = {9'd68,-10'd132};
ram[27201] = {9'd71,-10'd129};
ram[27202] = {9'd74,-10'd126};
ram[27203] = {9'd77,-10'd123};
ram[27204] = {9'd80,-10'd120};
ram[27205] = {9'd84,-10'd117};
ram[27206] = {9'd87,-10'd114};
ram[27207] = {9'd90,-10'd110};
ram[27208] = {9'd93,-10'd107};
ram[27209] = {9'd96,-10'd104};
ram[27210] = {9'd99,-10'd101};
ram[27211] = {-9'd98,-10'd98};
ram[27212] = {-9'd95,-10'd95};
ram[27213] = {-9'd92,-10'd92};
ram[27214] = {-9'd88,-10'd88};
ram[27215] = {-9'd85,-10'd85};
ram[27216] = {-9'd82,-10'd82};
ram[27217] = {-9'd79,-10'd79};
ram[27218] = {-9'd76,-10'd76};
ram[27219] = {-9'd73,-10'd73};
ram[27220] = {-9'd70,-10'd70};
ram[27221] = {-9'd66,-10'd66};
ram[27222] = {-9'd63,-10'd63};
ram[27223] = {-9'd60,-10'd60};
ram[27224] = {-9'd57,-10'd57};
ram[27225] = {-9'd54,-10'd54};
ram[27226] = {-9'd51,-10'd51};
ram[27227] = {-9'd48,-10'd48};
ram[27228] = {-9'd44,-10'd44};
ram[27229] = {-9'd41,-10'd41};
ram[27230] = {-9'd38,-10'd38};
ram[27231] = {-9'd35,-10'd35};
ram[27232] = {-9'd32,-10'd32};
ram[27233] = {-9'd29,-10'd29};
ram[27234] = {-9'd26,-10'd26};
ram[27235] = {-9'd22,-10'd22};
ram[27236] = {-9'd19,-10'd19};
ram[27237] = {-9'd16,-10'd16};
ram[27238] = {-9'd13,-10'd13};
ram[27239] = {-9'd10,-10'd10};
ram[27240] = {-9'd7,-10'd7};
ram[27241] = {-9'd4,-10'd4};
ram[27242] = {9'd0,10'd0};
ram[27243] = {9'd3,10'd3};
ram[27244] = {9'd6,10'd6};
ram[27245] = {9'd9,10'd9};
ram[27246] = {9'd12,10'd12};
ram[27247] = {9'd15,10'd15};
ram[27248] = {9'd18,10'd18};
ram[27249] = {9'd21,10'd21};
ram[27250] = {9'd25,10'd25};
ram[27251] = {9'd28,10'd28};
ram[27252] = {9'd31,10'd31};
ram[27253] = {9'd34,10'd34};
ram[27254] = {9'd37,10'd37};
ram[27255] = {9'd40,10'd40};
ram[27256] = {9'd43,10'd43};
ram[27257] = {9'd47,10'd47};
ram[27258] = {9'd50,10'd50};
ram[27259] = {9'd53,10'd53};
ram[27260] = {9'd56,10'd56};
ram[27261] = {9'd59,10'd59};
ram[27262] = {9'd62,10'd62};
ram[27263] = {9'd65,10'd65};
ram[27264] = {9'd65,10'd65};
ram[27265] = {9'd69,10'd69};
ram[27266] = {9'd72,10'd72};
ram[27267] = {9'd75,10'd75};
ram[27268] = {9'd78,10'd78};
ram[27269] = {9'd81,10'd81};
ram[27270] = {9'd84,10'd84};
ram[27271] = {9'd87,10'd87};
ram[27272] = {9'd91,10'd91};
ram[27273] = {9'd94,10'd94};
ram[27274] = {9'd97,10'd97};
ram[27275] = {-9'd100,10'd100};
ram[27276] = {-9'd97,10'd103};
ram[27277] = {-9'd94,10'd106};
ram[27278] = {-9'd91,10'd109};
ram[27279] = {-9'd88,10'd113};
ram[27280] = {-9'd85,10'd116};
ram[27281] = {-9'd81,10'd119};
ram[27282] = {-9'd78,10'd122};
ram[27283] = {-9'd75,10'd125};
ram[27284] = {-9'd72,10'd128};
ram[27285] = {-9'd69,10'd131};
ram[27286] = {-9'd66,10'd135};
ram[27287] = {-9'd63,10'd138};
ram[27288] = {-9'd59,10'd141};
ram[27289] = {-9'd56,10'd144};
ram[27290] = {-9'd53,10'd147};
ram[27291] = {-9'd50,10'd150};
ram[27292] = {-9'd47,10'd153};
ram[27293] = {-9'd44,10'd157};
ram[27294] = {-9'd41,10'd160};
ram[27295] = {-9'd37,10'd163};
ram[27296] = {-9'd34,10'd166};
ram[27297] = {-9'd31,10'd169};
ram[27298] = {-9'd28,10'd172};
ram[27299] = {-9'd25,10'd175};
ram[27300] = {-9'd22,10'd179};
ram[27301] = {-9'd19,10'd182};
ram[27302] = {-9'd15,10'd185};
ram[27303] = {-9'd12,10'd188};
ram[27304] = {-9'd9,10'd191};
ram[27305] = {-9'd6,10'd194};
ram[27306] = {-9'd3,10'd197};
ram[27307] = {9'd0,10'd201};
ram[27308] = {9'd3,10'd204};
ram[27309] = {9'd7,10'd207};
ram[27310] = {9'd10,10'd210};
ram[27311] = {9'd13,10'd213};
ram[27312] = {9'd16,10'd216};
ram[27313] = {9'd19,10'd219};
ram[27314] = {9'd22,10'd223};
ram[27315] = {9'd25,10'd226};
ram[27316] = {9'd29,10'd229};
ram[27317] = {9'd32,10'd232};
ram[27318] = {9'd35,10'd235};
ram[27319] = {9'd38,10'd238};
ram[27320] = {9'd41,10'd241};
ram[27321] = {9'd44,10'd245};
ram[27322] = {9'd47,10'd248};
ram[27323] = {9'd51,10'd251};
ram[27324] = {9'd54,10'd254};
ram[27325] = {9'd57,10'd257};
ram[27326] = {9'd60,10'd260};
ram[27327] = {9'd63,10'd263};
ram[27328] = {9'd66,10'd267};
ram[27329] = {9'd69,10'd270};
ram[27330] = {9'd73,10'd273};
ram[27331] = {9'd76,10'd276};
ram[27332] = {9'd79,10'd279};
ram[27333] = {9'd82,10'd282};
ram[27334] = {9'd85,10'd285};
ram[27335] = {9'd88,10'd289};
ram[27336] = {9'd91,10'd292};
ram[27337] = {9'd95,10'd295};
ram[27338] = {9'd98,10'd298};
ram[27339] = {-9'd99,10'd301};
ram[27340] = {-9'd96,10'd304};
ram[27341] = {-9'd93,10'd307};
ram[27342] = {-9'd90,10'd311};
ram[27343] = {-9'd87,10'd314};
ram[27344] = {-9'd84,10'd317};
ram[27345] = {-9'd81,10'd320};
ram[27346] = {-9'd77,10'd323};
ram[27347] = {-9'd74,10'd326};
ram[27348] = {-9'd71,10'd329};
ram[27349] = {-9'd68,10'd333};
ram[27350] = {-9'd65,10'd336};
ram[27351] = {-9'd62,10'd339};
ram[27352] = {-9'd59,10'd342};
ram[27353] = {-9'd55,10'd345};
ram[27354] = {-9'd52,10'd348};
ram[27355] = {-9'd49,10'd351};
ram[27356] = {-9'd46,10'd354};
ram[27357] = {-9'd43,10'd358};
ram[27358] = {-9'd40,10'd361};
ram[27359] = {-9'd37,10'd364};
ram[27360] = {-9'd33,10'd367};
ram[27361] = {-9'd30,10'd370};
ram[27362] = {-9'd27,10'd373};
ram[27363] = {-9'd24,10'd376};
ram[27364] = {-9'd21,10'd380};
ram[27365] = {-9'd18,10'd383};
ram[27366] = {-9'd15,10'd386};
ram[27367] = {-9'd11,10'd389};
ram[27368] = {-9'd8,10'd392};
ram[27369] = {-9'd5,10'd395};
ram[27370] = {-9'd2,10'd398};
ram[27371] = {9'd1,-10'd399};
ram[27372] = {9'd4,-10'd396};
ram[27373] = {9'd7,-10'd393};
ram[27374] = {9'd10,-10'd390};
ram[27375] = {9'd14,-10'd387};
ram[27376] = {9'd17,-10'd384};
ram[27377] = {9'd20,-10'd381};
ram[27378] = {9'd23,-10'd377};
ram[27379] = {9'd26,-10'd374};
ram[27380] = {9'd29,-10'd371};
ram[27381] = {9'd32,-10'd368};
ram[27382] = {9'd36,-10'd365};
ram[27383] = {9'd39,-10'd362};
ram[27384] = {9'd42,-10'd359};
ram[27385] = {9'd45,-10'd355};
ram[27386] = {9'd48,-10'd352};
ram[27387] = {9'd51,-10'd349};
ram[27388] = {9'd54,-10'd346};
ram[27389] = {9'd58,-10'd343};
ram[27390] = {9'd61,-10'd340};
ram[27391] = {9'd64,-10'd337};
ram[27392] = {9'd64,-10'd337};
ram[27393] = {9'd67,-10'd334};
ram[27394] = {9'd70,-10'd330};
ram[27395] = {9'd73,-10'd327};
ram[27396] = {9'd76,-10'd324};
ram[27397] = {9'd80,-10'd321};
ram[27398] = {9'd83,-10'd318};
ram[27399] = {9'd86,-10'd315};
ram[27400] = {9'd89,-10'd312};
ram[27401] = {9'd92,-10'd308};
ram[27402] = {9'd95,-10'd305};
ram[27403] = {9'd98,-10'd302};
ram[27404] = {-9'd99,-10'd299};
ram[27405] = {-9'd96,-10'd296};
ram[27406] = {-9'd92,-10'd293};
ram[27407] = {-9'd89,-10'd290};
ram[27408] = {-9'd86,-10'd286};
ram[27409] = {-9'd83,-10'd283};
ram[27410] = {-9'd80,-10'd280};
ram[27411] = {-9'd77,-10'd277};
ram[27412] = {-9'd74,-10'd274};
ram[27413] = {-9'd70,-10'd271};
ram[27414] = {-9'd67,-10'd268};
ram[27415] = {-9'd64,-10'd264};
ram[27416] = {-9'd61,-10'd261};
ram[27417] = {-9'd58,-10'd258};
ram[27418] = {-9'd55,-10'd255};
ram[27419] = {-9'd52,-10'd252};
ram[27420] = {-9'd48,-10'd249};
ram[27421] = {-9'd45,-10'd246};
ram[27422] = {-9'd42,-10'd242};
ram[27423] = {-9'd39,-10'd239};
ram[27424] = {-9'd36,-10'd236};
ram[27425] = {-9'd33,-10'd233};
ram[27426] = {-9'd30,-10'd230};
ram[27427] = {-9'd26,-10'd227};
ram[27428] = {-9'd23,-10'd224};
ram[27429] = {-9'd20,-10'd220};
ram[27430] = {-9'd17,-10'd217};
ram[27431] = {-9'd14,-10'd214};
ram[27432] = {-9'd11,-10'd211};
ram[27433] = {-9'd8,-10'd208};
ram[27434] = {-9'd4,-10'd205};
ram[27435] = {-9'd1,-10'd202};
ram[27436] = {9'd2,-10'd198};
ram[27437] = {9'd5,-10'd195};
ram[27438] = {9'd8,-10'd192};
ram[27439] = {9'd11,-10'd189};
ram[27440] = {9'd14,-10'd186};
ram[27441] = {9'd18,-10'd183};
ram[27442] = {9'd21,-10'd180};
ram[27443] = {9'd24,-10'd176};
ram[27444] = {9'd27,-10'd173};
ram[27445] = {9'd30,-10'd170};
ram[27446] = {9'd33,-10'd167};
ram[27447] = {9'd36,-10'd164};
ram[27448] = {9'd40,-10'd161};
ram[27449] = {9'd43,-10'd158};
ram[27450] = {9'd46,-10'd154};
ram[27451] = {9'd49,-10'd151};
ram[27452] = {9'd52,-10'd148};
ram[27453] = {9'd55,-10'd145};
ram[27454] = {9'd58,-10'd142};
ram[27455] = {9'd62,-10'd139};
ram[27456] = {9'd65,-10'd136};
ram[27457] = {9'd68,-10'd132};
ram[27458] = {9'd71,-10'd129};
ram[27459] = {9'd74,-10'd126};
ram[27460] = {9'd77,-10'd123};
ram[27461] = {9'd80,-10'd120};
ram[27462] = {9'd84,-10'd117};
ram[27463] = {9'd87,-10'd114};
ram[27464] = {9'd90,-10'd110};
ram[27465] = {9'd93,-10'd107};
ram[27466] = {9'd96,-10'd104};
ram[27467] = {9'd99,-10'd101};
ram[27468] = {-9'd98,-10'd98};
ram[27469] = {-9'd95,-10'd95};
ram[27470] = {-9'd92,-10'd92};
ram[27471] = {-9'd88,-10'd88};
ram[27472] = {-9'd85,-10'd85};
ram[27473] = {-9'd82,-10'd82};
ram[27474] = {-9'd79,-10'd79};
ram[27475] = {-9'd76,-10'd76};
ram[27476] = {-9'd73,-10'd73};
ram[27477] = {-9'd70,-10'd70};
ram[27478] = {-9'd66,-10'd66};
ram[27479] = {-9'd63,-10'd63};
ram[27480] = {-9'd60,-10'd60};
ram[27481] = {-9'd57,-10'd57};
ram[27482] = {-9'd54,-10'd54};
ram[27483] = {-9'd51,-10'd51};
ram[27484] = {-9'd48,-10'd48};
ram[27485] = {-9'd44,-10'd44};
ram[27486] = {-9'd41,-10'd41};
ram[27487] = {-9'd38,-10'd38};
ram[27488] = {-9'd35,-10'd35};
ram[27489] = {-9'd32,-10'd32};
ram[27490] = {-9'd29,-10'd29};
ram[27491] = {-9'd26,-10'd26};
ram[27492] = {-9'd22,-10'd22};
ram[27493] = {-9'd19,-10'd19};
ram[27494] = {-9'd16,-10'd16};
ram[27495] = {-9'd13,-10'd13};
ram[27496] = {-9'd10,-10'd10};
ram[27497] = {-9'd7,-10'd7};
ram[27498] = {-9'd4,-10'd4};
ram[27499] = {9'd0,10'd0};
ram[27500] = {9'd3,10'd3};
ram[27501] = {9'd6,10'd6};
ram[27502] = {9'd9,10'd9};
ram[27503] = {9'd12,10'd12};
ram[27504] = {9'd15,10'd15};
ram[27505] = {9'd18,10'd18};
ram[27506] = {9'd21,10'd21};
ram[27507] = {9'd25,10'd25};
ram[27508] = {9'd28,10'd28};
ram[27509] = {9'd31,10'd31};
ram[27510] = {9'd34,10'd34};
ram[27511] = {9'd37,10'd37};
ram[27512] = {9'd40,10'd40};
ram[27513] = {9'd43,10'd43};
ram[27514] = {9'd47,10'd47};
ram[27515] = {9'd50,10'd50};
ram[27516] = {9'd53,10'd53};
ram[27517] = {9'd56,10'd56};
ram[27518] = {9'd59,10'd59};
ram[27519] = {9'd62,10'd62};
ram[27520] = {9'd62,10'd62};
ram[27521] = {9'd65,10'd65};
ram[27522] = {9'd69,10'd69};
ram[27523] = {9'd72,10'd72};
ram[27524] = {9'd75,10'd75};
ram[27525] = {9'd78,10'd78};
ram[27526] = {9'd81,10'd81};
ram[27527] = {9'd84,10'd84};
ram[27528] = {9'd87,10'd87};
ram[27529] = {9'd91,10'd91};
ram[27530] = {9'd94,10'd94};
ram[27531] = {9'd97,10'd97};
ram[27532] = {-9'd100,10'd100};
ram[27533] = {-9'd97,10'd103};
ram[27534] = {-9'd94,10'd106};
ram[27535] = {-9'd91,10'd109};
ram[27536] = {-9'd88,10'd113};
ram[27537] = {-9'd85,10'd116};
ram[27538] = {-9'd81,10'd119};
ram[27539] = {-9'd78,10'd122};
ram[27540] = {-9'd75,10'd125};
ram[27541] = {-9'd72,10'd128};
ram[27542] = {-9'd69,10'd131};
ram[27543] = {-9'd66,10'd135};
ram[27544] = {-9'd63,10'd138};
ram[27545] = {-9'd59,10'd141};
ram[27546] = {-9'd56,10'd144};
ram[27547] = {-9'd53,10'd147};
ram[27548] = {-9'd50,10'd150};
ram[27549] = {-9'd47,10'd153};
ram[27550] = {-9'd44,10'd157};
ram[27551] = {-9'd41,10'd160};
ram[27552] = {-9'd37,10'd163};
ram[27553] = {-9'd34,10'd166};
ram[27554] = {-9'd31,10'd169};
ram[27555] = {-9'd28,10'd172};
ram[27556] = {-9'd25,10'd175};
ram[27557] = {-9'd22,10'd179};
ram[27558] = {-9'd19,10'd182};
ram[27559] = {-9'd15,10'd185};
ram[27560] = {-9'd12,10'd188};
ram[27561] = {-9'd9,10'd191};
ram[27562] = {-9'd6,10'd194};
ram[27563] = {-9'd3,10'd197};
ram[27564] = {9'd0,10'd201};
ram[27565] = {9'd3,10'd204};
ram[27566] = {9'd7,10'd207};
ram[27567] = {9'd10,10'd210};
ram[27568] = {9'd13,10'd213};
ram[27569] = {9'd16,10'd216};
ram[27570] = {9'd19,10'd219};
ram[27571] = {9'd22,10'd223};
ram[27572] = {9'd25,10'd226};
ram[27573] = {9'd29,10'd229};
ram[27574] = {9'd32,10'd232};
ram[27575] = {9'd35,10'd235};
ram[27576] = {9'd38,10'd238};
ram[27577] = {9'd41,10'd241};
ram[27578] = {9'd44,10'd245};
ram[27579] = {9'd47,10'd248};
ram[27580] = {9'd51,10'd251};
ram[27581] = {9'd54,10'd254};
ram[27582] = {9'd57,10'd257};
ram[27583] = {9'd60,10'd260};
ram[27584] = {9'd63,10'd263};
ram[27585] = {9'd66,10'd267};
ram[27586] = {9'd69,10'd270};
ram[27587] = {9'd73,10'd273};
ram[27588] = {9'd76,10'd276};
ram[27589] = {9'd79,10'd279};
ram[27590] = {9'd82,10'd282};
ram[27591] = {9'd85,10'd285};
ram[27592] = {9'd88,10'd289};
ram[27593] = {9'd91,10'd292};
ram[27594] = {9'd95,10'd295};
ram[27595] = {9'd98,10'd298};
ram[27596] = {-9'd99,10'd301};
ram[27597] = {-9'd96,10'd304};
ram[27598] = {-9'd93,10'd307};
ram[27599] = {-9'd90,10'd311};
ram[27600] = {-9'd87,10'd314};
ram[27601] = {-9'd84,10'd317};
ram[27602] = {-9'd81,10'd320};
ram[27603] = {-9'd77,10'd323};
ram[27604] = {-9'd74,10'd326};
ram[27605] = {-9'd71,10'd329};
ram[27606] = {-9'd68,10'd333};
ram[27607] = {-9'd65,10'd336};
ram[27608] = {-9'd62,10'd339};
ram[27609] = {-9'd59,10'd342};
ram[27610] = {-9'd55,10'd345};
ram[27611] = {-9'd52,10'd348};
ram[27612] = {-9'd49,10'd351};
ram[27613] = {-9'd46,10'd354};
ram[27614] = {-9'd43,10'd358};
ram[27615] = {-9'd40,10'd361};
ram[27616] = {-9'd37,10'd364};
ram[27617] = {-9'd33,10'd367};
ram[27618] = {-9'd30,10'd370};
ram[27619] = {-9'd27,10'd373};
ram[27620] = {-9'd24,10'd376};
ram[27621] = {-9'd21,10'd380};
ram[27622] = {-9'd18,10'd383};
ram[27623] = {-9'd15,10'd386};
ram[27624] = {-9'd11,10'd389};
ram[27625] = {-9'd8,10'd392};
ram[27626] = {-9'd5,10'd395};
ram[27627] = {-9'd2,10'd398};
ram[27628] = {9'd1,-10'd399};
ram[27629] = {9'd4,-10'd396};
ram[27630] = {9'd7,-10'd393};
ram[27631] = {9'd10,-10'd390};
ram[27632] = {9'd14,-10'd387};
ram[27633] = {9'd17,-10'd384};
ram[27634] = {9'd20,-10'd381};
ram[27635] = {9'd23,-10'd377};
ram[27636] = {9'd26,-10'd374};
ram[27637] = {9'd29,-10'd371};
ram[27638] = {9'd32,-10'd368};
ram[27639] = {9'd36,-10'd365};
ram[27640] = {9'd39,-10'd362};
ram[27641] = {9'd42,-10'd359};
ram[27642] = {9'd45,-10'd355};
ram[27643] = {9'd48,-10'd352};
ram[27644] = {9'd51,-10'd349};
ram[27645] = {9'd54,-10'd346};
ram[27646] = {9'd58,-10'd343};
ram[27647] = {9'd61,-10'd340};
ram[27648] = {9'd61,-10'd340};
ram[27649] = {9'd64,-10'd337};
ram[27650] = {9'd67,-10'd334};
ram[27651] = {9'd70,-10'd330};
ram[27652] = {9'd73,-10'd327};
ram[27653] = {9'd76,-10'd324};
ram[27654] = {9'd80,-10'd321};
ram[27655] = {9'd83,-10'd318};
ram[27656] = {9'd86,-10'd315};
ram[27657] = {9'd89,-10'd312};
ram[27658] = {9'd92,-10'd308};
ram[27659] = {9'd95,-10'd305};
ram[27660] = {9'd98,-10'd302};
ram[27661] = {-9'd99,-10'd299};
ram[27662] = {-9'd96,-10'd296};
ram[27663] = {-9'd92,-10'd293};
ram[27664] = {-9'd89,-10'd290};
ram[27665] = {-9'd86,-10'd286};
ram[27666] = {-9'd83,-10'd283};
ram[27667] = {-9'd80,-10'd280};
ram[27668] = {-9'd77,-10'd277};
ram[27669] = {-9'd74,-10'd274};
ram[27670] = {-9'd70,-10'd271};
ram[27671] = {-9'd67,-10'd268};
ram[27672] = {-9'd64,-10'd264};
ram[27673] = {-9'd61,-10'd261};
ram[27674] = {-9'd58,-10'd258};
ram[27675] = {-9'd55,-10'd255};
ram[27676] = {-9'd52,-10'd252};
ram[27677] = {-9'd48,-10'd249};
ram[27678] = {-9'd45,-10'd246};
ram[27679] = {-9'd42,-10'd242};
ram[27680] = {-9'd39,-10'd239};
ram[27681] = {-9'd36,-10'd236};
ram[27682] = {-9'd33,-10'd233};
ram[27683] = {-9'd30,-10'd230};
ram[27684] = {-9'd26,-10'd227};
ram[27685] = {-9'd23,-10'd224};
ram[27686] = {-9'd20,-10'd220};
ram[27687] = {-9'd17,-10'd217};
ram[27688] = {-9'd14,-10'd214};
ram[27689] = {-9'd11,-10'd211};
ram[27690] = {-9'd8,-10'd208};
ram[27691] = {-9'd4,-10'd205};
ram[27692] = {-9'd1,-10'd202};
ram[27693] = {9'd2,-10'd198};
ram[27694] = {9'd5,-10'd195};
ram[27695] = {9'd8,-10'd192};
ram[27696] = {9'd11,-10'd189};
ram[27697] = {9'd14,-10'd186};
ram[27698] = {9'd18,-10'd183};
ram[27699] = {9'd21,-10'd180};
ram[27700] = {9'd24,-10'd176};
ram[27701] = {9'd27,-10'd173};
ram[27702] = {9'd30,-10'd170};
ram[27703] = {9'd33,-10'd167};
ram[27704] = {9'd36,-10'd164};
ram[27705] = {9'd40,-10'd161};
ram[27706] = {9'd43,-10'd158};
ram[27707] = {9'd46,-10'd154};
ram[27708] = {9'd49,-10'd151};
ram[27709] = {9'd52,-10'd148};
ram[27710] = {9'd55,-10'd145};
ram[27711] = {9'd58,-10'd142};
ram[27712] = {9'd62,-10'd139};
ram[27713] = {9'd65,-10'd136};
ram[27714] = {9'd68,-10'd132};
ram[27715] = {9'd71,-10'd129};
ram[27716] = {9'd74,-10'd126};
ram[27717] = {9'd77,-10'd123};
ram[27718] = {9'd80,-10'd120};
ram[27719] = {9'd84,-10'd117};
ram[27720] = {9'd87,-10'd114};
ram[27721] = {9'd90,-10'd110};
ram[27722] = {9'd93,-10'd107};
ram[27723] = {9'd96,-10'd104};
ram[27724] = {9'd99,-10'd101};
ram[27725] = {-9'd98,-10'd98};
ram[27726] = {-9'd95,-10'd95};
ram[27727] = {-9'd92,-10'd92};
ram[27728] = {-9'd88,-10'd88};
ram[27729] = {-9'd85,-10'd85};
ram[27730] = {-9'd82,-10'd82};
ram[27731] = {-9'd79,-10'd79};
ram[27732] = {-9'd76,-10'd76};
ram[27733] = {-9'd73,-10'd73};
ram[27734] = {-9'd70,-10'd70};
ram[27735] = {-9'd66,-10'd66};
ram[27736] = {-9'd63,-10'd63};
ram[27737] = {-9'd60,-10'd60};
ram[27738] = {-9'd57,-10'd57};
ram[27739] = {-9'd54,-10'd54};
ram[27740] = {-9'd51,-10'd51};
ram[27741] = {-9'd48,-10'd48};
ram[27742] = {-9'd44,-10'd44};
ram[27743] = {-9'd41,-10'd41};
ram[27744] = {-9'd38,-10'd38};
ram[27745] = {-9'd35,-10'd35};
ram[27746] = {-9'd32,-10'd32};
ram[27747] = {-9'd29,-10'd29};
ram[27748] = {-9'd26,-10'd26};
ram[27749] = {-9'd22,-10'd22};
ram[27750] = {-9'd19,-10'd19};
ram[27751] = {-9'd16,-10'd16};
ram[27752] = {-9'd13,-10'd13};
ram[27753] = {-9'd10,-10'd10};
ram[27754] = {-9'd7,-10'd7};
ram[27755] = {-9'd4,-10'd4};
ram[27756] = {9'd0,10'd0};
ram[27757] = {9'd3,10'd3};
ram[27758] = {9'd6,10'd6};
ram[27759] = {9'd9,10'd9};
ram[27760] = {9'd12,10'd12};
ram[27761] = {9'd15,10'd15};
ram[27762] = {9'd18,10'd18};
ram[27763] = {9'd21,10'd21};
ram[27764] = {9'd25,10'd25};
ram[27765] = {9'd28,10'd28};
ram[27766] = {9'd31,10'd31};
ram[27767] = {9'd34,10'd34};
ram[27768] = {9'd37,10'd37};
ram[27769] = {9'd40,10'd40};
ram[27770] = {9'd43,10'd43};
ram[27771] = {9'd47,10'd47};
ram[27772] = {9'd50,10'd50};
ram[27773] = {9'd53,10'd53};
ram[27774] = {9'd56,10'd56};
ram[27775] = {9'd59,10'd59};
ram[27776] = {9'd59,10'd59};
ram[27777] = {9'd62,10'd62};
ram[27778] = {9'd65,10'd65};
ram[27779] = {9'd69,10'd69};
ram[27780] = {9'd72,10'd72};
ram[27781] = {9'd75,10'd75};
ram[27782] = {9'd78,10'd78};
ram[27783] = {9'd81,10'd81};
ram[27784] = {9'd84,10'd84};
ram[27785] = {9'd87,10'd87};
ram[27786] = {9'd91,10'd91};
ram[27787] = {9'd94,10'd94};
ram[27788] = {9'd97,10'd97};
ram[27789] = {-9'd100,10'd100};
ram[27790] = {-9'd97,10'd103};
ram[27791] = {-9'd94,10'd106};
ram[27792] = {-9'd91,10'd109};
ram[27793] = {-9'd88,10'd113};
ram[27794] = {-9'd85,10'd116};
ram[27795] = {-9'd81,10'd119};
ram[27796] = {-9'd78,10'd122};
ram[27797] = {-9'd75,10'd125};
ram[27798] = {-9'd72,10'd128};
ram[27799] = {-9'd69,10'd131};
ram[27800] = {-9'd66,10'd135};
ram[27801] = {-9'd63,10'd138};
ram[27802] = {-9'd59,10'd141};
ram[27803] = {-9'd56,10'd144};
ram[27804] = {-9'd53,10'd147};
ram[27805] = {-9'd50,10'd150};
ram[27806] = {-9'd47,10'd153};
ram[27807] = {-9'd44,10'd157};
ram[27808] = {-9'd41,10'd160};
ram[27809] = {-9'd37,10'd163};
ram[27810] = {-9'd34,10'd166};
ram[27811] = {-9'd31,10'd169};
ram[27812] = {-9'd28,10'd172};
ram[27813] = {-9'd25,10'd175};
ram[27814] = {-9'd22,10'd179};
ram[27815] = {-9'd19,10'd182};
ram[27816] = {-9'd15,10'd185};
ram[27817] = {-9'd12,10'd188};
ram[27818] = {-9'd9,10'd191};
ram[27819] = {-9'd6,10'd194};
ram[27820] = {-9'd3,10'd197};
ram[27821] = {9'd0,10'd201};
ram[27822] = {9'd3,10'd204};
ram[27823] = {9'd7,10'd207};
ram[27824] = {9'd10,10'd210};
ram[27825] = {9'd13,10'd213};
ram[27826] = {9'd16,10'd216};
ram[27827] = {9'd19,10'd219};
ram[27828] = {9'd22,10'd223};
ram[27829] = {9'd25,10'd226};
ram[27830] = {9'd29,10'd229};
ram[27831] = {9'd32,10'd232};
ram[27832] = {9'd35,10'd235};
ram[27833] = {9'd38,10'd238};
ram[27834] = {9'd41,10'd241};
ram[27835] = {9'd44,10'd245};
ram[27836] = {9'd47,10'd248};
ram[27837] = {9'd51,10'd251};
ram[27838] = {9'd54,10'd254};
ram[27839] = {9'd57,10'd257};
ram[27840] = {9'd60,10'd260};
ram[27841] = {9'd63,10'd263};
ram[27842] = {9'd66,10'd267};
ram[27843] = {9'd69,10'd270};
ram[27844] = {9'd73,10'd273};
ram[27845] = {9'd76,10'd276};
ram[27846] = {9'd79,10'd279};
ram[27847] = {9'd82,10'd282};
ram[27848] = {9'd85,10'd285};
ram[27849] = {9'd88,10'd289};
ram[27850] = {9'd91,10'd292};
ram[27851] = {9'd95,10'd295};
ram[27852] = {9'd98,10'd298};
ram[27853] = {-9'd99,10'd301};
ram[27854] = {-9'd96,10'd304};
ram[27855] = {-9'd93,10'd307};
ram[27856] = {-9'd90,10'd311};
ram[27857] = {-9'd87,10'd314};
ram[27858] = {-9'd84,10'd317};
ram[27859] = {-9'd81,10'd320};
ram[27860] = {-9'd77,10'd323};
ram[27861] = {-9'd74,10'd326};
ram[27862] = {-9'd71,10'd329};
ram[27863] = {-9'd68,10'd333};
ram[27864] = {-9'd65,10'd336};
ram[27865] = {-9'd62,10'd339};
ram[27866] = {-9'd59,10'd342};
ram[27867] = {-9'd55,10'd345};
ram[27868] = {-9'd52,10'd348};
ram[27869] = {-9'd49,10'd351};
ram[27870] = {-9'd46,10'd354};
ram[27871] = {-9'd43,10'd358};
ram[27872] = {-9'd40,10'd361};
ram[27873] = {-9'd37,10'd364};
ram[27874] = {-9'd33,10'd367};
ram[27875] = {-9'd30,10'd370};
ram[27876] = {-9'd27,10'd373};
ram[27877] = {-9'd24,10'd376};
ram[27878] = {-9'd21,10'd380};
ram[27879] = {-9'd18,10'd383};
ram[27880] = {-9'd15,10'd386};
ram[27881] = {-9'd11,10'd389};
ram[27882] = {-9'd8,10'd392};
ram[27883] = {-9'd5,10'd395};
ram[27884] = {-9'd2,10'd398};
ram[27885] = {9'd1,-10'd399};
ram[27886] = {9'd4,-10'd396};
ram[27887] = {9'd7,-10'd393};
ram[27888] = {9'd10,-10'd390};
ram[27889] = {9'd14,-10'd387};
ram[27890] = {9'd17,-10'd384};
ram[27891] = {9'd20,-10'd381};
ram[27892] = {9'd23,-10'd377};
ram[27893] = {9'd26,-10'd374};
ram[27894] = {9'd29,-10'd371};
ram[27895] = {9'd32,-10'd368};
ram[27896] = {9'd36,-10'd365};
ram[27897] = {9'd39,-10'd362};
ram[27898] = {9'd42,-10'd359};
ram[27899] = {9'd45,-10'd355};
ram[27900] = {9'd48,-10'd352};
ram[27901] = {9'd51,-10'd349};
ram[27902] = {9'd54,-10'd346};
ram[27903] = {9'd58,-10'd343};
ram[27904] = {9'd58,-10'd343};
ram[27905] = {9'd61,-10'd340};
ram[27906] = {9'd64,-10'd337};
ram[27907] = {9'd67,-10'd334};
ram[27908] = {9'd70,-10'd330};
ram[27909] = {9'd73,-10'd327};
ram[27910] = {9'd76,-10'd324};
ram[27911] = {9'd80,-10'd321};
ram[27912] = {9'd83,-10'd318};
ram[27913] = {9'd86,-10'd315};
ram[27914] = {9'd89,-10'd312};
ram[27915] = {9'd92,-10'd308};
ram[27916] = {9'd95,-10'd305};
ram[27917] = {9'd98,-10'd302};
ram[27918] = {-9'd99,-10'd299};
ram[27919] = {-9'd96,-10'd296};
ram[27920] = {-9'd92,-10'd293};
ram[27921] = {-9'd89,-10'd290};
ram[27922] = {-9'd86,-10'd286};
ram[27923] = {-9'd83,-10'd283};
ram[27924] = {-9'd80,-10'd280};
ram[27925] = {-9'd77,-10'd277};
ram[27926] = {-9'd74,-10'd274};
ram[27927] = {-9'd70,-10'd271};
ram[27928] = {-9'd67,-10'd268};
ram[27929] = {-9'd64,-10'd264};
ram[27930] = {-9'd61,-10'd261};
ram[27931] = {-9'd58,-10'd258};
ram[27932] = {-9'd55,-10'd255};
ram[27933] = {-9'd52,-10'd252};
ram[27934] = {-9'd48,-10'd249};
ram[27935] = {-9'd45,-10'd246};
ram[27936] = {-9'd42,-10'd242};
ram[27937] = {-9'd39,-10'd239};
ram[27938] = {-9'd36,-10'd236};
ram[27939] = {-9'd33,-10'd233};
ram[27940] = {-9'd30,-10'd230};
ram[27941] = {-9'd26,-10'd227};
ram[27942] = {-9'd23,-10'd224};
ram[27943] = {-9'd20,-10'd220};
ram[27944] = {-9'd17,-10'd217};
ram[27945] = {-9'd14,-10'd214};
ram[27946] = {-9'd11,-10'd211};
ram[27947] = {-9'd8,-10'd208};
ram[27948] = {-9'd4,-10'd205};
ram[27949] = {-9'd1,-10'd202};
ram[27950] = {9'd2,-10'd198};
ram[27951] = {9'd5,-10'd195};
ram[27952] = {9'd8,-10'd192};
ram[27953] = {9'd11,-10'd189};
ram[27954] = {9'd14,-10'd186};
ram[27955] = {9'd18,-10'd183};
ram[27956] = {9'd21,-10'd180};
ram[27957] = {9'd24,-10'd176};
ram[27958] = {9'd27,-10'd173};
ram[27959] = {9'd30,-10'd170};
ram[27960] = {9'd33,-10'd167};
ram[27961] = {9'd36,-10'd164};
ram[27962] = {9'd40,-10'd161};
ram[27963] = {9'd43,-10'd158};
ram[27964] = {9'd46,-10'd154};
ram[27965] = {9'd49,-10'd151};
ram[27966] = {9'd52,-10'd148};
ram[27967] = {9'd55,-10'd145};
ram[27968] = {9'd58,-10'd142};
ram[27969] = {9'd62,-10'd139};
ram[27970] = {9'd65,-10'd136};
ram[27971] = {9'd68,-10'd132};
ram[27972] = {9'd71,-10'd129};
ram[27973] = {9'd74,-10'd126};
ram[27974] = {9'd77,-10'd123};
ram[27975] = {9'd80,-10'd120};
ram[27976] = {9'd84,-10'd117};
ram[27977] = {9'd87,-10'd114};
ram[27978] = {9'd90,-10'd110};
ram[27979] = {9'd93,-10'd107};
ram[27980] = {9'd96,-10'd104};
ram[27981] = {9'd99,-10'd101};
ram[27982] = {-9'd98,-10'd98};
ram[27983] = {-9'd95,-10'd95};
ram[27984] = {-9'd92,-10'd92};
ram[27985] = {-9'd88,-10'd88};
ram[27986] = {-9'd85,-10'd85};
ram[27987] = {-9'd82,-10'd82};
ram[27988] = {-9'd79,-10'd79};
ram[27989] = {-9'd76,-10'd76};
ram[27990] = {-9'd73,-10'd73};
ram[27991] = {-9'd70,-10'd70};
ram[27992] = {-9'd66,-10'd66};
ram[27993] = {-9'd63,-10'd63};
ram[27994] = {-9'd60,-10'd60};
ram[27995] = {-9'd57,-10'd57};
ram[27996] = {-9'd54,-10'd54};
ram[27997] = {-9'd51,-10'd51};
ram[27998] = {-9'd48,-10'd48};
ram[27999] = {-9'd44,-10'd44};
ram[28000] = {-9'd41,-10'd41};
ram[28001] = {-9'd38,-10'd38};
ram[28002] = {-9'd35,-10'd35};
ram[28003] = {-9'd32,-10'd32};
ram[28004] = {-9'd29,-10'd29};
ram[28005] = {-9'd26,-10'd26};
ram[28006] = {-9'd22,-10'd22};
ram[28007] = {-9'd19,-10'd19};
ram[28008] = {-9'd16,-10'd16};
ram[28009] = {-9'd13,-10'd13};
ram[28010] = {-9'd10,-10'd10};
ram[28011] = {-9'd7,-10'd7};
ram[28012] = {-9'd4,-10'd4};
ram[28013] = {9'd0,10'd0};
ram[28014] = {9'd3,10'd3};
ram[28015] = {9'd6,10'd6};
ram[28016] = {9'd9,10'd9};
ram[28017] = {9'd12,10'd12};
ram[28018] = {9'd15,10'd15};
ram[28019] = {9'd18,10'd18};
ram[28020] = {9'd21,10'd21};
ram[28021] = {9'd25,10'd25};
ram[28022] = {9'd28,10'd28};
ram[28023] = {9'd31,10'd31};
ram[28024] = {9'd34,10'd34};
ram[28025] = {9'd37,10'd37};
ram[28026] = {9'd40,10'd40};
ram[28027] = {9'd43,10'd43};
ram[28028] = {9'd47,10'd47};
ram[28029] = {9'd50,10'd50};
ram[28030] = {9'd53,10'd53};
ram[28031] = {9'd56,10'd56};
ram[28032] = {9'd56,10'd56};
ram[28033] = {9'd59,10'd59};
ram[28034] = {9'd62,10'd62};
ram[28035] = {9'd65,10'd65};
ram[28036] = {9'd69,10'd69};
ram[28037] = {9'd72,10'd72};
ram[28038] = {9'd75,10'd75};
ram[28039] = {9'd78,10'd78};
ram[28040] = {9'd81,10'd81};
ram[28041] = {9'd84,10'd84};
ram[28042] = {9'd87,10'd87};
ram[28043] = {9'd91,10'd91};
ram[28044] = {9'd94,10'd94};
ram[28045] = {9'd97,10'd97};
ram[28046] = {-9'd100,10'd100};
ram[28047] = {-9'd97,10'd103};
ram[28048] = {-9'd94,10'd106};
ram[28049] = {-9'd91,10'd109};
ram[28050] = {-9'd88,10'd113};
ram[28051] = {-9'd85,10'd116};
ram[28052] = {-9'd81,10'd119};
ram[28053] = {-9'd78,10'd122};
ram[28054] = {-9'd75,10'd125};
ram[28055] = {-9'd72,10'd128};
ram[28056] = {-9'd69,10'd131};
ram[28057] = {-9'd66,10'd135};
ram[28058] = {-9'd63,10'd138};
ram[28059] = {-9'd59,10'd141};
ram[28060] = {-9'd56,10'd144};
ram[28061] = {-9'd53,10'd147};
ram[28062] = {-9'd50,10'd150};
ram[28063] = {-9'd47,10'd153};
ram[28064] = {-9'd44,10'd157};
ram[28065] = {-9'd41,10'd160};
ram[28066] = {-9'd37,10'd163};
ram[28067] = {-9'd34,10'd166};
ram[28068] = {-9'd31,10'd169};
ram[28069] = {-9'd28,10'd172};
ram[28070] = {-9'd25,10'd175};
ram[28071] = {-9'd22,10'd179};
ram[28072] = {-9'd19,10'd182};
ram[28073] = {-9'd15,10'd185};
ram[28074] = {-9'd12,10'd188};
ram[28075] = {-9'd9,10'd191};
ram[28076] = {-9'd6,10'd194};
ram[28077] = {-9'd3,10'd197};
ram[28078] = {9'd0,10'd201};
ram[28079] = {9'd3,10'd204};
ram[28080] = {9'd7,10'd207};
ram[28081] = {9'd10,10'd210};
ram[28082] = {9'd13,10'd213};
ram[28083] = {9'd16,10'd216};
ram[28084] = {9'd19,10'd219};
ram[28085] = {9'd22,10'd223};
ram[28086] = {9'd25,10'd226};
ram[28087] = {9'd29,10'd229};
ram[28088] = {9'd32,10'd232};
ram[28089] = {9'd35,10'd235};
ram[28090] = {9'd38,10'd238};
ram[28091] = {9'd41,10'd241};
ram[28092] = {9'd44,10'd245};
ram[28093] = {9'd47,10'd248};
ram[28094] = {9'd51,10'd251};
ram[28095] = {9'd54,10'd254};
ram[28096] = {9'd57,10'd257};
ram[28097] = {9'd60,10'd260};
ram[28098] = {9'd63,10'd263};
ram[28099] = {9'd66,10'd267};
ram[28100] = {9'd69,10'd270};
ram[28101] = {9'd73,10'd273};
ram[28102] = {9'd76,10'd276};
ram[28103] = {9'd79,10'd279};
ram[28104] = {9'd82,10'd282};
ram[28105] = {9'd85,10'd285};
ram[28106] = {9'd88,10'd289};
ram[28107] = {9'd91,10'd292};
ram[28108] = {9'd95,10'd295};
ram[28109] = {9'd98,10'd298};
ram[28110] = {-9'd99,10'd301};
ram[28111] = {-9'd96,10'd304};
ram[28112] = {-9'd93,10'd307};
ram[28113] = {-9'd90,10'd311};
ram[28114] = {-9'd87,10'd314};
ram[28115] = {-9'd84,10'd317};
ram[28116] = {-9'd81,10'd320};
ram[28117] = {-9'd77,10'd323};
ram[28118] = {-9'd74,10'd326};
ram[28119] = {-9'd71,10'd329};
ram[28120] = {-9'd68,10'd333};
ram[28121] = {-9'd65,10'd336};
ram[28122] = {-9'd62,10'd339};
ram[28123] = {-9'd59,10'd342};
ram[28124] = {-9'd55,10'd345};
ram[28125] = {-9'd52,10'd348};
ram[28126] = {-9'd49,10'd351};
ram[28127] = {-9'd46,10'd354};
ram[28128] = {-9'd43,10'd358};
ram[28129] = {-9'd40,10'd361};
ram[28130] = {-9'd37,10'd364};
ram[28131] = {-9'd33,10'd367};
ram[28132] = {-9'd30,10'd370};
ram[28133] = {-9'd27,10'd373};
ram[28134] = {-9'd24,10'd376};
ram[28135] = {-9'd21,10'd380};
ram[28136] = {-9'd18,10'd383};
ram[28137] = {-9'd15,10'd386};
ram[28138] = {-9'd11,10'd389};
ram[28139] = {-9'd8,10'd392};
ram[28140] = {-9'd5,10'd395};
ram[28141] = {-9'd2,10'd398};
ram[28142] = {9'd1,-10'd399};
ram[28143] = {9'd4,-10'd396};
ram[28144] = {9'd7,-10'd393};
ram[28145] = {9'd10,-10'd390};
ram[28146] = {9'd14,-10'd387};
ram[28147] = {9'd17,-10'd384};
ram[28148] = {9'd20,-10'd381};
ram[28149] = {9'd23,-10'd377};
ram[28150] = {9'd26,-10'd374};
ram[28151] = {9'd29,-10'd371};
ram[28152] = {9'd32,-10'd368};
ram[28153] = {9'd36,-10'd365};
ram[28154] = {9'd39,-10'd362};
ram[28155] = {9'd42,-10'd359};
ram[28156] = {9'd45,-10'd355};
ram[28157] = {9'd48,-10'd352};
ram[28158] = {9'd51,-10'd349};
ram[28159] = {9'd54,-10'd346};
ram[28160] = {9'd54,-10'd346};
ram[28161] = {9'd58,-10'd343};
ram[28162] = {9'd61,-10'd340};
ram[28163] = {9'd64,-10'd337};
ram[28164] = {9'd67,-10'd334};
ram[28165] = {9'd70,-10'd330};
ram[28166] = {9'd73,-10'd327};
ram[28167] = {9'd76,-10'd324};
ram[28168] = {9'd80,-10'd321};
ram[28169] = {9'd83,-10'd318};
ram[28170] = {9'd86,-10'd315};
ram[28171] = {9'd89,-10'd312};
ram[28172] = {9'd92,-10'd308};
ram[28173] = {9'd95,-10'd305};
ram[28174] = {9'd98,-10'd302};
ram[28175] = {-9'd99,-10'd299};
ram[28176] = {-9'd96,-10'd296};
ram[28177] = {-9'd92,-10'd293};
ram[28178] = {-9'd89,-10'd290};
ram[28179] = {-9'd86,-10'd286};
ram[28180] = {-9'd83,-10'd283};
ram[28181] = {-9'd80,-10'd280};
ram[28182] = {-9'd77,-10'd277};
ram[28183] = {-9'd74,-10'd274};
ram[28184] = {-9'd70,-10'd271};
ram[28185] = {-9'd67,-10'd268};
ram[28186] = {-9'd64,-10'd264};
ram[28187] = {-9'd61,-10'd261};
ram[28188] = {-9'd58,-10'd258};
ram[28189] = {-9'd55,-10'd255};
ram[28190] = {-9'd52,-10'd252};
ram[28191] = {-9'd48,-10'd249};
ram[28192] = {-9'd45,-10'd246};
ram[28193] = {-9'd42,-10'd242};
ram[28194] = {-9'd39,-10'd239};
ram[28195] = {-9'd36,-10'd236};
ram[28196] = {-9'd33,-10'd233};
ram[28197] = {-9'd30,-10'd230};
ram[28198] = {-9'd26,-10'd227};
ram[28199] = {-9'd23,-10'd224};
ram[28200] = {-9'd20,-10'd220};
ram[28201] = {-9'd17,-10'd217};
ram[28202] = {-9'd14,-10'd214};
ram[28203] = {-9'd11,-10'd211};
ram[28204] = {-9'd8,-10'd208};
ram[28205] = {-9'd4,-10'd205};
ram[28206] = {-9'd1,-10'd202};
ram[28207] = {9'd2,-10'd198};
ram[28208] = {9'd5,-10'd195};
ram[28209] = {9'd8,-10'd192};
ram[28210] = {9'd11,-10'd189};
ram[28211] = {9'd14,-10'd186};
ram[28212] = {9'd18,-10'd183};
ram[28213] = {9'd21,-10'd180};
ram[28214] = {9'd24,-10'd176};
ram[28215] = {9'd27,-10'd173};
ram[28216] = {9'd30,-10'd170};
ram[28217] = {9'd33,-10'd167};
ram[28218] = {9'd36,-10'd164};
ram[28219] = {9'd40,-10'd161};
ram[28220] = {9'd43,-10'd158};
ram[28221] = {9'd46,-10'd154};
ram[28222] = {9'd49,-10'd151};
ram[28223] = {9'd52,-10'd148};
ram[28224] = {9'd55,-10'd145};
ram[28225] = {9'd58,-10'd142};
ram[28226] = {9'd62,-10'd139};
ram[28227] = {9'd65,-10'd136};
ram[28228] = {9'd68,-10'd132};
ram[28229] = {9'd71,-10'd129};
ram[28230] = {9'd74,-10'd126};
ram[28231] = {9'd77,-10'd123};
ram[28232] = {9'd80,-10'd120};
ram[28233] = {9'd84,-10'd117};
ram[28234] = {9'd87,-10'd114};
ram[28235] = {9'd90,-10'd110};
ram[28236] = {9'd93,-10'd107};
ram[28237] = {9'd96,-10'd104};
ram[28238] = {9'd99,-10'd101};
ram[28239] = {-9'd98,-10'd98};
ram[28240] = {-9'd95,-10'd95};
ram[28241] = {-9'd92,-10'd92};
ram[28242] = {-9'd88,-10'd88};
ram[28243] = {-9'd85,-10'd85};
ram[28244] = {-9'd82,-10'd82};
ram[28245] = {-9'd79,-10'd79};
ram[28246] = {-9'd76,-10'd76};
ram[28247] = {-9'd73,-10'd73};
ram[28248] = {-9'd70,-10'd70};
ram[28249] = {-9'd66,-10'd66};
ram[28250] = {-9'd63,-10'd63};
ram[28251] = {-9'd60,-10'd60};
ram[28252] = {-9'd57,-10'd57};
ram[28253] = {-9'd54,-10'd54};
ram[28254] = {-9'd51,-10'd51};
ram[28255] = {-9'd48,-10'd48};
ram[28256] = {-9'd44,-10'd44};
ram[28257] = {-9'd41,-10'd41};
ram[28258] = {-9'd38,-10'd38};
ram[28259] = {-9'd35,-10'd35};
ram[28260] = {-9'd32,-10'd32};
ram[28261] = {-9'd29,-10'd29};
ram[28262] = {-9'd26,-10'd26};
ram[28263] = {-9'd22,-10'd22};
ram[28264] = {-9'd19,-10'd19};
ram[28265] = {-9'd16,-10'd16};
ram[28266] = {-9'd13,-10'd13};
ram[28267] = {-9'd10,-10'd10};
ram[28268] = {-9'd7,-10'd7};
ram[28269] = {-9'd4,-10'd4};
ram[28270] = {9'd0,10'd0};
ram[28271] = {9'd3,10'd3};
ram[28272] = {9'd6,10'd6};
ram[28273] = {9'd9,10'd9};
ram[28274] = {9'd12,10'd12};
ram[28275] = {9'd15,10'd15};
ram[28276] = {9'd18,10'd18};
ram[28277] = {9'd21,10'd21};
ram[28278] = {9'd25,10'd25};
ram[28279] = {9'd28,10'd28};
ram[28280] = {9'd31,10'd31};
ram[28281] = {9'd34,10'd34};
ram[28282] = {9'd37,10'd37};
ram[28283] = {9'd40,10'd40};
ram[28284] = {9'd43,10'd43};
ram[28285] = {9'd47,10'd47};
ram[28286] = {9'd50,10'd50};
ram[28287] = {9'd53,10'd53};
ram[28288] = {9'd53,10'd53};
ram[28289] = {9'd56,10'd56};
ram[28290] = {9'd59,10'd59};
ram[28291] = {9'd62,10'd62};
ram[28292] = {9'd65,10'd65};
ram[28293] = {9'd69,10'd69};
ram[28294] = {9'd72,10'd72};
ram[28295] = {9'd75,10'd75};
ram[28296] = {9'd78,10'd78};
ram[28297] = {9'd81,10'd81};
ram[28298] = {9'd84,10'd84};
ram[28299] = {9'd87,10'd87};
ram[28300] = {9'd91,10'd91};
ram[28301] = {9'd94,10'd94};
ram[28302] = {9'd97,10'd97};
ram[28303] = {-9'd100,10'd100};
ram[28304] = {-9'd97,10'd103};
ram[28305] = {-9'd94,10'd106};
ram[28306] = {-9'd91,10'd109};
ram[28307] = {-9'd88,10'd113};
ram[28308] = {-9'd85,10'd116};
ram[28309] = {-9'd81,10'd119};
ram[28310] = {-9'd78,10'd122};
ram[28311] = {-9'd75,10'd125};
ram[28312] = {-9'd72,10'd128};
ram[28313] = {-9'd69,10'd131};
ram[28314] = {-9'd66,10'd135};
ram[28315] = {-9'd63,10'd138};
ram[28316] = {-9'd59,10'd141};
ram[28317] = {-9'd56,10'd144};
ram[28318] = {-9'd53,10'd147};
ram[28319] = {-9'd50,10'd150};
ram[28320] = {-9'd47,10'd153};
ram[28321] = {-9'd44,10'd157};
ram[28322] = {-9'd41,10'd160};
ram[28323] = {-9'd37,10'd163};
ram[28324] = {-9'd34,10'd166};
ram[28325] = {-9'd31,10'd169};
ram[28326] = {-9'd28,10'd172};
ram[28327] = {-9'd25,10'd175};
ram[28328] = {-9'd22,10'd179};
ram[28329] = {-9'd19,10'd182};
ram[28330] = {-9'd15,10'd185};
ram[28331] = {-9'd12,10'd188};
ram[28332] = {-9'd9,10'd191};
ram[28333] = {-9'd6,10'd194};
ram[28334] = {-9'd3,10'd197};
ram[28335] = {9'd0,10'd201};
ram[28336] = {9'd3,10'd204};
ram[28337] = {9'd7,10'd207};
ram[28338] = {9'd10,10'd210};
ram[28339] = {9'd13,10'd213};
ram[28340] = {9'd16,10'd216};
ram[28341] = {9'd19,10'd219};
ram[28342] = {9'd22,10'd223};
ram[28343] = {9'd25,10'd226};
ram[28344] = {9'd29,10'd229};
ram[28345] = {9'd32,10'd232};
ram[28346] = {9'd35,10'd235};
ram[28347] = {9'd38,10'd238};
ram[28348] = {9'd41,10'd241};
ram[28349] = {9'd44,10'd245};
ram[28350] = {9'd47,10'd248};
ram[28351] = {9'd51,10'd251};
ram[28352] = {9'd54,10'd254};
ram[28353] = {9'd57,10'd257};
ram[28354] = {9'd60,10'd260};
ram[28355] = {9'd63,10'd263};
ram[28356] = {9'd66,10'd267};
ram[28357] = {9'd69,10'd270};
ram[28358] = {9'd73,10'd273};
ram[28359] = {9'd76,10'd276};
ram[28360] = {9'd79,10'd279};
ram[28361] = {9'd82,10'd282};
ram[28362] = {9'd85,10'd285};
ram[28363] = {9'd88,10'd289};
ram[28364] = {9'd91,10'd292};
ram[28365] = {9'd95,10'd295};
ram[28366] = {9'd98,10'd298};
ram[28367] = {-9'd99,10'd301};
ram[28368] = {-9'd96,10'd304};
ram[28369] = {-9'd93,10'd307};
ram[28370] = {-9'd90,10'd311};
ram[28371] = {-9'd87,10'd314};
ram[28372] = {-9'd84,10'd317};
ram[28373] = {-9'd81,10'd320};
ram[28374] = {-9'd77,10'd323};
ram[28375] = {-9'd74,10'd326};
ram[28376] = {-9'd71,10'd329};
ram[28377] = {-9'd68,10'd333};
ram[28378] = {-9'd65,10'd336};
ram[28379] = {-9'd62,10'd339};
ram[28380] = {-9'd59,10'd342};
ram[28381] = {-9'd55,10'd345};
ram[28382] = {-9'd52,10'd348};
ram[28383] = {-9'd49,10'd351};
ram[28384] = {-9'd46,10'd354};
ram[28385] = {-9'd43,10'd358};
ram[28386] = {-9'd40,10'd361};
ram[28387] = {-9'd37,10'd364};
ram[28388] = {-9'd33,10'd367};
ram[28389] = {-9'd30,10'd370};
ram[28390] = {-9'd27,10'd373};
ram[28391] = {-9'd24,10'd376};
ram[28392] = {-9'd21,10'd380};
ram[28393] = {-9'd18,10'd383};
ram[28394] = {-9'd15,10'd386};
ram[28395] = {-9'd11,10'd389};
ram[28396] = {-9'd8,10'd392};
ram[28397] = {-9'd5,10'd395};
ram[28398] = {-9'd2,10'd398};
ram[28399] = {9'd1,-10'd399};
ram[28400] = {9'd4,-10'd396};
ram[28401] = {9'd7,-10'd393};
ram[28402] = {9'd10,-10'd390};
ram[28403] = {9'd14,-10'd387};
ram[28404] = {9'd17,-10'd384};
ram[28405] = {9'd20,-10'd381};
ram[28406] = {9'd23,-10'd377};
ram[28407] = {9'd26,-10'd374};
ram[28408] = {9'd29,-10'd371};
ram[28409] = {9'd32,-10'd368};
ram[28410] = {9'd36,-10'd365};
ram[28411] = {9'd39,-10'd362};
ram[28412] = {9'd42,-10'd359};
ram[28413] = {9'd45,-10'd355};
ram[28414] = {9'd48,-10'd352};
ram[28415] = {9'd51,-10'd349};
ram[28416] = {9'd51,-10'd349};
ram[28417] = {9'd54,-10'd346};
ram[28418] = {9'd58,-10'd343};
ram[28419] = {9'd61,-10'd340};
ram[28420] = {9'd64,-10'd337};
ram[28421] = {9'd67,-10'd334};
ram[28422] = {9'd70,-10'd330};
ram[28423] = {9'd73,-10'd327};
ram[28424] = {9'd76,-10'd324};
ram[28425] = {9'd80,-10'd321};
ram[28426] = {9'd83,-10'd318};
ram[28427] = {9'd86,-10'd315};
ram[28428] = {9'd89,-10'd312};
ram[28429] = {9'd92,-10'd308};
ram[28430] = {9'd95,-10'd305};
ram[28431] = {9'd98,-10'd302};
ram[28432] = {-9'd99,-10'd299};
ram[28433] = {-9'd96,-10'd296};
ram[28434] = {-9'd92,-10'd293};
ram[28435] = {-9'd89,-10'd290};
ram[28436] = {-9'd86,-10'd286};
ram[28437] = {-9'd83,-10'd283};
ram[28438] = {-9'd80,-10'd280};
ram[28439] = {-9'd77,-10'd277};
ram[28440] = {-9'd74,-10'd274};
ram[28441] = {-9'd70,-10'd271};
ram[28442] = {-9'd67,-10'd268};
ram[28443] = {-9'd64,-10'd264};
ram[28444] = {-9'd61,-10'd261};
ram[28445] = {-9'd58,-10'd258};
ram[28446] = {-9'd55,-10'd255};
ram[28447] = {-9'd52,-10'd252};
ram[28448] = {-9'd48,-10'd249};
ram[28449] = {-9'd45,-10'd246};
ram[28450] = {-9'd42,-10'd242};
ram[28451] = {-9'd39,-10'd239};
ram[28452] = {-9'd36,-10'd236};
ram[28453] = {-9'd33,-10'd233};
ram[28454] = {-9'd30,-10'd230};
ram[28455] = {-9'd26,-10'd227};
ram[28456] = {-9'd23,-10'd224};
ram[28457] = {-9'd20,-10'd220};
ram[28458] = {-9'd17,-10'd217};
ram[28459] = {-9'd14,-10'd214};
ram[28460] = {-9'd11,-10'd211};
ram[28461] = {-9'd8,-10'd208};
ram[28462] = {-9'd4,-10'd205};
ram[28463] = {-9'd1,-10'd202};
ram[28464] = {9'd2,-10'd198};
ram[28465] = {9'd5,-10'd195};
ram[28466] = {9'd8,-10'd192};
ram[28467] = {9'd11,-10'd189};
ram[28468] = {9'd14,-10'd186};
ram[28469] = {9'd18,-10'd183};
ram[28470] = {9'd21,-10'd180};
ram[28471] = {9'd24,-10'd176};
ram[28472] = {9'd27,-10'd173};
ram[28473] = {9'd30,-10'd170};
ram[28474] = {9'd33,-10'd167};
ram[28475] = {9'd36,-10'd164};
ram[28476] = {9'd40,-10'd161};
ram[28477] = {9'd43,-10'd158};
ram[28478] = {9'd46,-10'd154};
ram[28479] = {9'd49,-10'd151};
ram[28480] = {9'd52,-10'd148};
ram[28481] = {9'd55,-10'd145};
ram[28482] = {9'd58,-10'd142};
ram[28483] = {9'd62,-10'd139};
ram[28484] = {9'd65,-10'd136};
ram[28485] = {9'd68,-10'd132};
ram[28486] = {9'd71,-10'd129};
ram[28487] = {9'd74,-10'd126};
ram[28488] = {9'd77,-10'd123};
ram[28489] = {9'd80,-10'd120};
ram[28490] = {9'd84,-10'd117};
ram[28491] = {9'd87,-10'd114};
ram[28492] = {9'd90,-10'd110};
ram[28493] = {9'd93,-10'd107};
ram[28494] = {9'd96,-10'd104};
ram[28495] = {9'd99,-10'd101};
ram[28496] = {-9'd98,-10'd98};
ram[28497] = {-9'd95,-10'd95};
ram[28498] = {-9'd92,-10'd92};
ram[28499] = {-9'd88,-10'd88};
ram[28500] = {-9'd85,-10'd85};
ram[28501] = {-9'd82,-10'd82};
ram[28502] = {-9'd79,-10'd79};
ram[28503] = {-9'd76,-10'd76};
ram[28504] = {-9'd73,-10'd73};
ram[28505] = {-9'd70,-10'd70};
ram[28506] = {-9'd66,-10'd66};
ram[28507] = {-9'd63,-10'd63};
ram[28508] = {-9'd60,-10'd60};
ram[28509] = {-9'd57,-10'd57};
ram[28510] = {-9'd54,-10'd54};
ram[28511] = {-9'd51,-10'd51};
ram[28512] = {-9'd48,-10'd48};
ram[28513] = {-9'd44,-10'd44};
ram[28514] = {-9'd41,-10'd41};
ram[28515] = {-9'd38,-10'd38};
ram[28516] = {-9'd35,-10'd35};
ram[28517] = {-9'd32,-10'd32};
ram[28518] = {-9'd29,-10'd29};
ram[28519] = {-9'd26,-10'd26};
ram[28520] = {-9'd22,-10'd22};
ram[28521] = {-9'd19,-10'd19};
ram[28522] = {-9'd16,-10'd16};
ram[28523] = {-9'd13,-10'd13};
ram[28524] = {-9'd10,-10'd10};
ram[28525] = {-9'd7,-10'd7};
ram[28526] = {-9'd4,-10'd4};
ram[28527] = {9'd0,10'd0};
ram[28528] = {9'd3,10'd3};
ram[28529] = {9'd6,10'd6};
ram[28530] = {9'd9,10'd9};
ram[28531] = {9'd12,10'd12};
ram[28532] = {9'd15,10'd15};
ram[28533] = {9'd18,10'd18};
ram[28534] = {9'd21,10'd21};
ram[28535] = {9'd25,10'd25};
ram[28536] = {9'd28,10'd28};
ram[28537] = {9'd31,10'd31};
ram[28538] = {9'd34,10'd34};
ram[28539] = {9'd37,10'd37};
ram[28540] = {9'd40,10'd40};
ram[28541] = {9'd43,10'd43};
ram[28542] = {9'd47,10'd47};
ram[28543] = {9'd50,10'd50};
ram[28544] = {9'd50,10'd50};
ram[28545] = {9'd53,10'd53};
ram[28546] = {9'd56,10'd56};
ram[28547] = {9'd59,10'd59};
ram[28548] = {9'd62,10'd62};
ram[28549] = {9'd65,10'd65};
ram[28550] = {9'd69,10'd69};
ram[28551] = {9'd72,10'd72};
ram[28552] = {9'd75,10'd75};
ram[28553] = {9'd78,10'd78};
ram[28554] = {9'd81,10'd81};
ram[28555] = {9'd84,10'd84};
ram[28556] = {9'd87,10'd87};
ram[28557] = {9'd91,10'd91};
ram[28558] = {9'd94,10'd94};
ram[28559] = {9'd97,10'd97};
ram[28560] = {-9'd100,10'd100};
ram[28561] = {-9'd97,10'd103};
ram[28562] = {-9'd94,10'd106};
ram[28563] = {-9'd91,10'd109};
ram[28564] = {-9'd88,10'd113};
ram[28565] = {-9'd85,10'd116};
ram[28566] = {-9'd81,10'd119};
ram[28567] = {-9'd78,10'd122};
ram[28568] = {-9'd75,10'd125};
ram[28569] = {-9'd72,10'd128};
ram[28570] = {-9'd69,10'd131};
ram[28571] = {-9'd66,10'd135};
ram[28572] = {-9'd63,10'd138};
ram[28573] = {-9'd59,10'd141};
ram[28574] = {-9'd56,10'd144};
ram[28575] = {-9'd53,10'd147};
ram[28576] = {-9'd50,10'd150};
ram[28577] = {-9'd47,10'd153};
ram[28578] = {-9'd44,10'd157};
ram[28579] = {-9'd41,10'd160};
ram[28580] = {-9'd37,10'd163};
ram[28581] = {-9'd34,10'd166};
ram[28582] = {-9'd31,10'd169};
ram[28583] = {-9'd28,10'd172};
ram[28584] = {-9'd25,10'd175};
ram[28585] = {-9'd22,10'd179};
ram[28586] = {-9'd19,10'd182};
ram[28587] = {-9'd15,10'd185};
ram[28588] = {-9'd12,10'd188};
ram[28589] = {-9'd9,10'd191};
ram[28590] = {-9'd6,10'd194};
ram[28591] = {-9'd3,10'd197};
ram[28592] = {9'd0,10'd201};
ram[28593] = {9'd3,10'd204};
ram[28594] = {9'd7,10'd207};
ram[28595] = {9'd10,10'd210};
ram[28596] = {9'd13,10'd213};
ram[28597] = {9'd16,10'd216};
ram[28598] = {9'd19,10'd219};
ram[28599] = {9'd22,10'd223};
ram[28600] = {9'd25,10'd226};
ram[28601] = {9'd29,10'd229};
ram[28602] = {9'd32,10'd232};
ram[28603] = {9'd35,10'd235};
ram[28604] = {9'd38,10'd238};
ram[28605] = {9'd41,10'd241};
ram[28606] = {9'd44,10'd245};
ram[28607] = {9'd47,10'd248};
ram[28608] = {9'd51,10'd251};
ram[28609] = {9'd54,10'd254};
ram[28610] = {9'd57,10'd257};
ram[28611] = {9'd60,10'd260};
ram[28612] = {9'd63,10'd263};
ram[28613] = {9'd66,10'd267};
ram[28614] = {9'd69,10'd270};
ram[28615] = {9'd73,10'd273};
ram[28616] = {9'd76,10'd276};
ram[28617] = {9'd79,10'd279};
ram[28618] = {9'd82,10'd282};
ram[28619] = {9'd85,10'd285};
ram[28620] = {9'd88,10'd289};
ram[28621] = {9'd91,10'd292};
ram[28622] = {9'd95,10'd295};
ram[28623] = {9'd98,10'd298};
ram[28624] = {-9'd99,10'd301};
ram[28625] = {-9'd96,10'd304};
ram[28626] = {-9'd93,10'd307};
ram[28627] = {-9'd90,10'd311};
ram[28628] = {-9'd87,10'd314};
ram[28629] = {-9'd84,10'd317};
ram[28630] = {-9'd81,10'd320};
ram[28631] = {-9'd77,10'd323};
ram[28632] = {-9'd74,10'd326};
ram[28633] = {-9'd71,10'd329};
ram[28634] = {-9'd68,10'd333};
ram[28635] = {-9'd65,10'd336};
ram[28636] = {-9'd62,10'd339};
ram[28637] = {-9'd59,10'd342};
ram[28638] = {-9'd55,10'd345};
ram[28639] = {-9'd52,10'd348};
ram[28640] = {-9'd49,10'd351};
ram[28641] = {-9'd46,10'd354};
ram[28642] = {-9'd43,10'd358};
ram[28643] = {-9'd40,10'd361};
ram[28644] = {-9'd37,10'd364};
ram[28645] = {-9'd33,10'd367};
ram[28646] = {-9'd30,10'd370};
ram[28647] = {-9'd27,10'd373};
ram[28648] = {-9'd24,10'd376};
ram[28649] = {-9'd21,10'd380};
ram[28650] = {-9'd18,10'd383};
ram[28651] = {-9'd15,10'd386};
ram[28652] = {-9'd11,10'd389};
ram[28653] = {-9'd8,10'd392};
ram[28654] = {-9'd5,10'd395};
ram[28655] = {-9'd2,10'd398};
ram[28656] = {9'd1,-10'd399};
ram[28657] = {9'd4,-10'd396};
ram[28658] = {9'd7,-10'd393};
ram[28659] = {9'd10,-10'd390};
ram[28660] = {9'd14,-10'd387};
ram[28661] = {9'd17,-10'd384};
ram[28662] = {9'd20,-10'd381};
ram[28663] = {9'd23,-10'd377};
ram[28664] = {9'd26,-10'd374};
ram[28665] = {9'd29,-10'd371};
ram[28666] = {9'd32,-10'd368};
ram[28667] = {9'd36,-10'd365};
ram[28668] = {9'd39,-10'd362};
ram[28669] = {9'd42,-10'd359};
ram[28670] = {9'd45,-10'd355};
ram[28671] = {9'd48,-10'd352};
ram[28672] = {9'd48,-10'd352};
ram[28673] = {9'd51,-10'd349};
ram[28674] = {9'd54,-10'd346};
ram[28675] = {9'd58,-10'd343};
ram[28676] = {9'd61,-10'd340};
ram[28677] = {9'd64,-10'd337};
ram[28678] = {9'd67,-10'd334};
ram[28679] = {9'd70,-10'd330};
ram[28680] = {9'd73,-10'd327};
ram[28681] = {9'd76,-10'd324};
ram[28682] = {9'd80,-10'd321};
ram[28683] = {9'd83,-10'd318};
ram[28684] = {9'd86,-10'd315};
ram[28685] = {9'd89,-10'd312};
ram[28686] = {9'd92,-10'd308};
ram[28687] = {9'd95,-10'd305};
ram[28688] = {9'd98,-10'd302};
ram[28689] = {-9'd99,-10'd299};
ram[28690] = {-9'd96,-10'd296};
ram[28691] = {-9'd92,-10'd293};
ram[28692] = {-9'd89,-10'd290};
ram[28693] = {-9'd86,-10'd286};
ram[28694] = {-9'd83,-10'd283};
ram[28695] = {-9'd80,-10'd280};
ram[28696] = {-9'd77,-10'd277};
ram[28697] = {-9'd74,-10'd274};
ram[28698] = {-9'd70,-10'd271};
ram[28699] = {-9'd67,-10'd268};
ram[28700] = {-9'd64,-10'd264};
ram[28701] = {-9'd61,-10'd261};
ram[28702] = {-9'd58,-10'd258};
ram[28703] = {-9'd55,-10'd255};
ram[28704] = {-9'd52,-10'd252};
ram[28705] = {-9'd48,-10'd249};
ram[28706] = {-9'd45,-10'd246};
ram[28707] = {-9'd42,-10'd242};
ram[28708] = {-9'd39,-10'd239};
ram[28709] = {-9'd36,-10'd236};
ram[28710] = {-9'd33,-10'd233};
ram[28711] = {-9'd30,-10'd230};
ram[28712] = {-9'd26,-10'd227};
ram[28713] = {-9'd23,-10'd224};
ram[28714] = {-9'd20,-10'd220};
ram[28715] = {-9'd17,-10'd217};
ram[28716] = {-9'd14,-10'd214};
ram[28717] = {-9'd11,-10'd211};
ram[28718] = {-9'd8,-10'd208};
ram[28719] = {-9'd4,-10'd205};
ram[28720] = {-9'd1,-10'd202};
ram[28721] = {9'd2,-10'd198};
ram[28722] = {9'd5,-10'd195};
ram[28723] = {9'd8,-10'd192};
ram[28724] = {9'd11,-10'd189};
ram[28725] = {9'd14,-10'd186};
ram[28726] = {9'd18,-10'd183};
ram[28727] = {9'd21,-10'd180};
ram[28728] = {9'd24,-10'd176};
ram[28729] = {9'd27,-10'd173};
ram[28730] = {9'd30,-10'd170};
ram[28731] = {9'd33,-10'd167};
ram[28732] = {9'd36,-10'd164};
ram[28733] = {9'd40,-10'd161};
ram[28734] = {9'd43,-10'd158};
ram[28735] = {9'd46,-10'd154};
ram[28736] = {9'd49,-10'd151};
ram[28737] = {9'd52,-10'd148};
ram[28738] = {9'd55,-10'd145};
ram[28739] = {9'd58,-10'd142};
ram[28740] = {9'd62,-10'd139};
ram[28741] = {9'd65,-10'd136};
ram[28742] = {9'd68,-10'd132};
ram[28743] = {9'd71,-10'd129};
ram[28744] = {9'd74,-10'd126};
ram[28745] = {9'd77,-10'd123};
ram[28746] = {9'd80,-10'd120};
ram[28747] = {9'd84,-10'd117};
ram[28748] = {9'd87,-10'd114};
ram[28749] = {9'd90,-10'd110};
ram[28750] = {9'd93,-10'd107};
ram[28751] = {9'd96,-10'd104};
ram[28752] = {9'd99,-10'd101};
ram[28753] = {-9'd98,-10'd98};
ram[28754] = {-9'd95,-10'd95};
ram[28755] = {-9'd92,-10'd92};
ram[28756] = {-9'd88,-10'd88};
ram[28757] = {-9'd85,-10'd85};
ram[28758] = {-9'd82,-10'd82};
ram[28759] = {-9'd79,-10'd79};
ram[28760] = {-9'd76,-10'd76};
ram[28761] = {-9'd73,-10'd73};
ram[28762] = {-9'd70,-10'd70};
ram[28763] = {-9'd66,-10'd66};
ram[28764] = {-9'd63,-10'd63};
ram[28765] = {-9'd60,-10'd60};
ram[28766] = {-9'd57,-10'd57};
ram[28767] = {-9'd54,-10'd54};
ram[28768] = {-9'd51,-10'd51};
ram[28769] = {-9'd48,-10'd48};
ram[28770] = {-9'd44,-10'd44};
ram[28771] = {-9'd41,-10'd41};
ram[28772] = {-9'd38,-10'd38};
ram[28773] = {-9'd35,-10'd35};
ram[28774] = {-9'd32,-10'd32};
ram[28775] = {-9'd29,-10'd29};
ram[28776] = {-9'd26,-10'd26};
ram[28777] = {-9'd22,-10'd22};
ram[28778] = {-9'd19,-10'd19};
ram[28779] = {-9'd16,-10'd16};
ram[28780] = {-9'd13,-10'd13};
ram[28781] = {-9'd10,-10'd10};
ram[28782] = {-9'd7,-10'd7};
ram[28783] = {-9'd4,-10'd4};
ram[28784] = {9'd0,10'd0};
ram[28785] = {9'd3,10'd3};
ram[28786] = {9'd6,10'd6};
ram[28787] = {9'd9,10'd9};
ram[28788] = {9'd12,10'd12};
ram[28789] = {9'd15,10'd15};
ram[28790] = {9'd18,10'd18};
ram[28791] = {9'd21,10'd21};
ram[28792] = {9'd25,10'd25};
ram[28793] = {9'd28,10'd28};
ram[28794] = {9'd31,10'd31};
ram[28795] = {9'd34,10'd34};
ram[28796] = {9'd37,10'd37};
ram[28797] = {9'd40,10'd40};
ram[28798] = {9'd43,10'd43};
ram[28799] = {9'd47,10'd47};
ram[28800] = {9'd47,10'd47};
ram[28801] = {9'd50,10'd50};
ram[28802] = {9'd53,10'd53};
ram[28803] = {9'd56,10'd56};
ram[28804] = {9'd59,10'd59};
ram[28805] = {9'd62,10'd62};
ram[28806] = {9'd65,10'd65};
ram[28807] = {9'd69,10'd69};
ram[28808] = {9'd72,10'd72};
ram[28809] = {9'd75,10'd75};
ram[28810] = {9'd78,10'd78};
ram[28811] = {9'd81,10'd81};
ram[28812] = {9'd84,10'd84};
ram[28813] = {9'd87,10'd87};
ram[28814] = {9'd91,10'd91};
ram[28815] = {9'd94,10'd94};
ram[28816] = {9'd97,10'd97};
ram[28817] = {-9'd100,10'd100};
ram[28818] = {-9'd97,10'd103};
ram[28819] = {-9'd94,10'd106};
ram[28820] = {-9'd91,10'd109};
ram[28821] = {-9'd88,10'd113};
ram[28822] = {-9'd85,10'd116};
ram[28823] = {-9'd81,10'd119};
ram[28824] = {-9'd78,10'd122};
ram[28825] = {-9'd75,10'd125};
ram[28826] = {-9'd72,10'd128};
ram[28827] = {-9'd69,10'd131};
ram[28828] = {-9'd66,10'd135};
ram[28829] = {-9'd63,10'd138};
ram[28830] = {-9'd59,10'd141};
ram[28831] = {-9'd56,10'd144};
ram[28832] = {-9'd53,10'd147};
ram[28833] = {-9'd50,10'd150};
ram[28834] = {-9'd47,10'd153};
ram[28835] = {-9'd44,10'd157};
ram[28836] = {-9'd41,10'd160};
ram[28837] = {-9'd37,10'd163};
ram[28838] = {-9'd34,10'd166};
ram[28839] = {-9'd31,10'd169};
ram[28840] = {-9'd28,10'd172};
ram[28841] = {-9'd25,10'd175};
ram[28842] = {-9'd22,10'd179};
ram[28843] = {-9'd19,10'd182};
ram[28844] = {-9'd15,10'd185};
ram[28845] = {-9'd12,10'd188};
ram[28846] = {-9'd9,10'd191};
ram[28847] = {-9'd6,10'd194};
ram[28848] = {-9'd3,10'd197};
ram[28849] = {9'd0,10'd201};
ram[28850] = {9'd3,10'd204};
ram[28851] = {9'd7,10'd207};
ram[28852] = {9'd10,10'd210};
ram[28853] = {9'd13,10'd213};
ram[28854] = {9'd16,10'd216};
ram[28855] = {9'd19,10'd219};
ram[28856] = {9'd22,10'd223};
ram[28857] = {9'd25,10'd226};
ram[28858] = {9'd29,10'd229};
ram[28859] = {9'd32,10'd232};
ram[28860] = {9'd35,10'd235};
ram[28861] = {9'd38,10'd238};
ram[28862] = {9'd41,10'd241};
ram[28863] = {9'd44,10'd245};
ram[28864] = {9'd47,10'd248};
ram[28865] = {9'd51,10'd251};
ram[28866] = {9'd54,10'd254};
ram[28867] = {9'd57,10'd257};
ram[28868] = {9'd60,10'd260};
ram[28869] = {9'd63,10'd263};
ram[28870] = {9'd66,10'd267};
ram[28871] = {9'd69,10'd270};
ram[28872] = {9'd73,10'd273};
ram[28873] = {9'd76,10'd276};
ram[28874] = {9'd79,10'd279};
ram[28875] = {9'd82,10'd282};
ram[28876] = {9'd85,10'd285};
ram[28877] = {9'd88,10'd289};
ram[28878] = {9'd91,10'd292};
ram[28879] = {9'd95,10'd295};
ram[28880] = {9'd98,10'd298};
ram[28881] = {-9'd99,10'd301};
ram[28882] = {-9'd96,10'd304};
ram[28883] = {-9'd93,10'd307};
ram[28884] = {-9'd90,10'd311};
ram[28885] = {-9'd87,10'd314};
ram[28886] = {-9'd84,10'd317};
ram[28887] = {-9'd81,10'd320};
ram[28888] = {-9'd77,10'd323};
ram[28889] = {-9'd74,10'd326};
ram[28890] = {-9'd71,10'd329};
ram[28891] = {-9'd68,10'd333};
ram[28892] = {-9'd65,10'd336};
ram[28893] = {-9'd62,10'd339};
ram[28894] = {-9'd59,10'd342};
ram[28895] = {-9'd55,10'd345};
ram[28896] = {-9'd52,10'd348};
ram[28897] = {-9'd49,10'd351};
ram[28898] = {-9'd46,10'd354};
ram[28899] = {-9'd43,10'd358};
ram[28900] = {-9'd40,10'd361};
ram[28901] = {-9'd37,10'd364};
ram[28902] = {-9'd33,10'd367};
ram[28903] = {-9'd30,10'd370};
ram[28904] = {-9'd27,10'd373};
ram[28905] = {-9'd24,10'd376};
ram[28906] = {-9'd21,10'd380};
ram[28907] = {-9'd18,10'd383};
ram[28908] = {-9'd15,10'd386};
ram[28909] = {-9'd11,10'd389};
ram[28910] = {-9'd8,10'd392};
ram[28911] = {-9'd5,10'd395};
ram[28912] = {-9'd2,10'd398};
ram[28913] = {9'd1,-10'd399};
ram[28914] = {9'd4,-10'd396};
ram[28915] = {9'd7,-10'd393};
ram[28916] = {9'd10,-10'd390};
ram[28917] = {9'd14,-10'd387};
ram[28918] = {9'd17,-10'd384};
ram[28919] = {9'd20,-10'd381};
ram[28920] = {9'd23,-10'd377};
ram[28921] = {9'd26,-10'd374};
ram[28922] = {9'd29,-10'd371};
ram[28923] = {9'd32,-10'd368};
ram[28924] = {9'd36,-10'd365};
ram[28925] = {9'd39,-10'd362};
ram[28926] = {9'd42,-10'd359};
ram[28927] = {9'd45,-10'd355};
ram[28928] = {9'd45,-10'd355};
ram[28929] = {9'd48,-10'd352};
ram[28930] = {9'd51,-10'd349};
ram[28931] = {9'd54,-10'd346};
ram[28932] = {9'd58,-10'd343};
ram[28933] = {9'd61,-10'd340};
ram[28934] = {9'd64,-10'd337};
ram[28935] = {9'd67,-10'd334};
ram[28936] = {9'd70,-10'd330};
ram[28937] = {9'd73,-10'd327};
ram[28938] = {9'd76,-10'd324};
ram[28939] = {9'd80,-10'd321};
ram[28940] = {9'd83,-10'd318};
ram[28941] = {9'd86,-10'd315};
ram[28942] = {9'd89,-10'd312};
ram[28943] = {9'd92,-10'd308};
ram[28944] = {9'd95,-10'd305};
ram[28945] = {9'd98,-10'd302};
ram[28946] = {-9'd99,-10'd299};
ram[28947] = {-9'd96,-10'd296};
ram[28948] = {-9'd92,-10'd293};
ram[28949] = {-9'd89,-10'd290};
ram[28950] = {-9'd86,-10'd286};
ram[28951] = {-9'd83,-10'd283};
ram[28952] = {-9'd80,-10'd280};
ram[28953] = {-9'd77,-10'd277};
ram[28954] = {-9'd74,-10'd274};
ram[28955] = {-9'd70,-10'd271};
ram[28956] = {-9'd67,-10'd268};
ram[28957] = {-9'd64,-10'd264};
ram[28958] = {-9'd61,-10'd261};
ram[28959] = {-9'd58,-10'd258};
ram[28960] = {-9'd55,-10'd255};
ram[28961] = {-9'd52,-10'd252};
ram[28962] = {-9'd48,-10'd249};
ram[28963] = {-9'd45,-10'd246};
ram[28964] = {-9'd42,-10'd242};
ram[28965] = {-9'd39,-10'd239};
ram[28966] = {-9'd36,-10'd236};
ram[28967] = {-9'd33,-10'd233};
ram[28968] = {-9'd30,-10'd230};
ram[28969] = {-9'd26,-10'd227};
ram[28970] = {-9'd23,-10'd224};
ram[28971] = {-9'd20,-10'd220};
ram[28972] = {-9'd17,-10'd217};
ram[28973] = {-9'd14,-10'd214};
ram[28974] = {-9'd11,-10'd211};
ram[28975] = {-9'd8,-10'd208};
ram[28976] = {-9'd4,-10'd205};
ram[28977] = {-9'd1,-10'd202};
ram[28978] = {9'd2,-10'd198};
ram[28979] = {9'd5,-10'd195};
ram[28980] = {9'd8,-10'd192};
ram[28981] = {9'd11,-10'd189};
ram[28982] = {9'd14,-10'd186};
ram[28983] = {9'd18,-10'd183};
ram[28984] = {9'd21,-10'd180};
ram[28985] = {9'd24,-10'd176};
ram[28986] = {9'd27,-10'd173};
ram[28987] = {9'd30,-10'd170};
ram[28988] = {9'd33,-10'd167};
ram[28989] = {9'd36,-10'd164};
ram[28990] = {9'd40,-10'd161};
ram[28991] = {9'd43,-10'd158};
ram[28992] = {9'd46,-10'd154};
ram[28993] = {9'd49,-10'd151};
ram[28994] = {9'd52,-10'd148};
ram[28995] = {9'd55,-10'd145};
ram[28996] = {9'd58,-10'd142};
ram[28997] = {9'd62,-10'd139};
ram[28998] = {9'd65,-10'd136};
ram[28999] = {9'd68,-10'd132};
ram[29000] = {9'd71,-10'd129};
ram[29001] = {9'd74,-10'd126};
ram[29002] = {9'd77,-10'd123};
ram[29003] = {9'd80,-10'd120};
ram[29004] = {9'd84,-10'd117};
ram[29005] = {9'd87,-10'd114};
ram[29006] = {9'd90,-10'd110};
ram[29007] = {9'd93,-10'd107};
ram[29008] = {9'd96,-10'd104};
ram[29009] = {9'd99,-10'd101};
ram[29010] = {-9'd98,-10'd98};
ram[29011] = {-9'd95,-10'd95};
ram[29012] = {-9'd92,-10'd92};
ram[29013] = {-9'd88,-10'd88};
ram[29014] = {-9'd85,-10'd85};
ram[29015] = {-9'd82,-10'd82};
ram[29016] = {-9'd79,-10'd79};
ram[29017] = {-9'd76,-10'd76};
ram[29018] = {-9'd73,-10'd73};
ram[29019] = {-9'd70,-10'd70};
ram[29020] = {-9'd66,-10'd66};
ram[29021] = {-9'd63,-10'd63};
ram[29022] = {-9'd60,-10'd60};
ram[29023] = {-9'd57,-10'd57};
ram[29024] = {-9'd54,-10'd54};
ram[29025] = {-9'd51,-10'd51};
ram[29026] = {-9'd48,-10'd48};
ram[29027] = {-9'd44,-10'd44};
ram[29028] = {-9'd41,-10'd41};
ram[29029] = {-9'd38,-10'd38};
ram[29030] = {-9'd35,-10'd35};
ram[29031] = {-9'd32,-10'd32};
ram[29032] = {-9'd29,-10'd29};
ram[29033] = {-9'd26,-10'd26};
ram[29034] = {-9'd22,-10'd22};
ram[29035] = {-9'd19,-10'd19};
ram[29036] = {-9'd16,-10'd16};
ram[29037] = {-9'd13,-10'd13};
ram[29038] = {-9'd10,-10'd10};
ram[29039] = {-9'd7,-10'd7};
ram[29040] = {-9'd4,-10'd4};
ram[29041] = {9'd0,10'd0};
ram[29042] = {9'd3,10'd3};
ram[29043] = {9'd6,10'd6};
ram[29044] = {9'd9,10'd9};
ram[29045] = {9'd12,10'd12};
ram[29046] = {9'd15,10'd15};
ram[29047] = {9'd18,10'd18};
ram[29048] = {9'd21,10'd21};
ram[29049] = {9'd25,10'd25};
ram[29050] = {9'd28,10'd28};
ram[29051] = {9'd31,10'd31};
ram[29052] = {9'd34,10'd34};
ram[29053] = {9'd37,10'd37};
ram[29054] = {9'd40,10'd40};
ram[29055] = {9'd43,10'd43};
ram[29056] = {9'd43,10'd43};
ram[29057] = {9'd47,10'd47};
ram[29058] = {9'd50,10'd50};
ram[29059] = {9'd53,10'd53};
ram[29060] = {9'd56,10'd56};
ram[29061] = {9'd59,10'd59};
ram[29062] = {9'd62,10'd62};
ram[29063] = {9'd65,10'd65};
ram[29064] = {9'd69,10'd69};
ram[29065] = {9'd72,10'd72};
ram[29066] = {9'd75,10'd75};
ram[29067] = {9'd78,10'd78};
ram[29068] = {9'd81,10'd81};
ram[29069] = {9'd84,10'd84};
ram[29070] = {9'd87,10'd87};
ram[29071] = {9'd91,10'd91};
ram[29072] = {9'd94,10'd94};
ram[29073] = {9'd97,10'd97};
ram[29074] = {-9'd100,10'd100};
ram[29075] = {-9'd97,10'd103};
ram[29076] = {-9'd94,10'd106};
ram[29077] = {-9'd91,10'd109};
ram[29078] = {-9'd88,10'd113};
ram[29079] = {-9'd85,10'd116};
ram[29080] = {-9'd81,10'd119};
ram[29081] = {-9'd78,10'd122};
ram[29082] = {-9'd75,10'd125};
ram[29083] = {-9'd72,10'd128};
ram[29084] = {-9'd69,10'd131};
ram[29085] = {-9'd66,10'd135};
ram[29086] = {-9'd63,10'd138};
ram[29087] = {-9'd59,10'd141};
ram[29088] = {-9'd56,10'd144};
ram[29089] = {-9'd53,10'd147};
ram[29090] = {-9'd50,10'd150};
ram[29091] = {-9'd47,10'd153};
ram[29092] = {-9'd44,10'd157};
ram[29093] = {-9'd41,10'd160};
ram[29094] = {-9'd37,10'd163};
ram[29095] = {-9'd34,10'd166};
ram[29096] = {-9'd31,10'd169};
ram[29097] = {-9'd28,10'd172};
ram[29098] = {-9'd25,10'd175};
ram[29099] = {-9'd22,10'd179};
ram[29100] = {-9'd19,10'd182};
ram[29101] = {-9'd15,10'd185};
ram[29102] = {-9'd12,10'd188};
ram[29103] = {-9'd9,10'd191};
ram[29104] = {-9'd6,10'd194};
ram[29105] = {-9'd3,10'd197};
ram[29106] = {9'd0,10'd201};
ram[29107] = {9'd3,10'd204};
ram[29108] = {9'd7,10'd207};
ram[29109] = {9'd10,10'd210};
ram[29110] = {9'd13,10'd213};
ram[29111] = {9'd16,10'd216};
ram[29112] = {9'd19,10'd219};
ram[29113] = {9'd22,10'd223};
ram[29114] = {9'd25,10'd226};
ram[29115] = {9'd29,10'd229};
ram[29116] = {9'd32,10'd232};
ram[29117] = {9'd35,10'd235};
ram[29118] = {9'd38,10'd238};
ram[29119] = {9'd41,10'd241};
ram[29120] = {9'd44,10'd245};
ram[29121] = {9'd47,10'd248};
ram[29122] = {9'd51,10'd251};
ram[29123] = {9'd54,10'd254};
ram[29124] = {9'd57,10'd257};
ram[29125] = {9'd60,10'd260};
ram[29126] = {9'd63,10'd263};
ram[29127] = {9'd66,10'd267};
ram[29128] = {9'd69,10'd270};
ram[29129] = {9'd73,10'd273};
ram[29130] = {9'd76,10'd276};
ram[29131] = {9'd79,10'd279};
ram[29132] = {9'd82,10'd282};
ram[29133] = {9'd85,10'd285};
ram[29134] = {9'd88,10'd289};
ram[29135] = {9'd91,10'd292};
ram[29136] = {9'd95,10'd295};
ram[29137] = {9'd98,10'd298};
ram[29138] = {-9'd99,10'd301};
ram[29139] = {-9'd96,10'd304};
ram[29140] = {-9'd93,10'd307};
ram[29141] = {-9'd90,10'd311};
ram[29142] = {-9'd87,10'd314};
ram[29143] = {-9'd84,10'd317};
ram[29144] = {-9'd81,10'd320};
ram[29145] = {-9'd77,10'd323};
ram[29146] = {-9'd74,10'd326};
ram[29147] = {-9'd71,10'd329};
ram[29148] = {-9'd68,10'd333};
ram[29149] = {-9'd65,10'd336};
ram[29150] = {-9'd62,10'd339};
ram[29151] = {-9'd59,10'd342};
ram[29152] = {-9'd55,10'd345};
ram[29153] = {-9'd52,10'd348};
ram[29154] = {-9'd49,10'd351};
ram[29155] = {-9'd46,10'd354};
ram[29156] = {-9'd43,10'd358};
ram[29157] = {-9'd40,10'd361};
ram[29158] = {-9'd37,10'd364};
ram[29159] = {-9'd33,10'd367};
ram[29160] = {-9'd30,10'd370};
ram[29161] = {-9'd27,10'd373};
ram[29162] = {-9'd24,10'd376};
ram[29163] = {-9'd21,10'd380};
ram[29164] = {-9'd18,10'd383};
ram[29165] = {-9'd15,10'd386};
ram[29166] = {-9'd11,10'd389};
ram[29167] = {-9'd8,10'd392};
ram[29168] = {-9'd5,10'd395};
ram[29169] = {-9'd2,10'd398};
ram[29170] = {9'd1,-10'd399};
ram[29171] = {9'd4,-10'd396};
ram[29172] = {9'd7,-10'd393};
ram[29173] = {9'd10,-10'd390};
ram[29174] = {9'd14,-10'd387};
ram[29175] = {9'd17,-10'd384};
ram[29176] = {9'd20,-10'd381};
ram[29177] = {9'd23,-10'd377};
ram[29178] = {9'd26,-10'd374};
ram[29179] = {9'd29,-10'd371};
ram[29180] = {9'd32,-10'd368};
ram[29181] = {9'd36,-10'd365};
ram[29182] = {9'd39,-10'd362};
ram[29183] = {9'd42,-10'd359};
ram[29184] = {9'd42,-10'd359};
ram[29185] = {9'd45,-10'd355};
ram[29186] = {9'd48,-10'd352};
ram[29187] = {9'd51,-10'd349};
ram[29188] = {9'd54,-10'd346};
ram[29189] = {9'd58,-10'd343};
ram[29190] = {9'd61,-10'd340};
ram[29191] = {9'd64,-10'd337};
ram[29192] = {9'd67,-10'd334};
ram[29193] = {9'd70,-10'd330};
ram[29194] = {9'd73,-10'd327};
ram[29195] = {9'd76,-10'd324};
ram[29196] = {9'd80,-10'd321};
ram[29197] = {9'd83,-10'd318};
ram[29198] = {9'd86,-10'd315};
ram[29199] = {9'd89,-10'd312};
ram[29200] = {9'd92,-10'd308};
ram[29201] = {9'd95,-10'd305};
ram[29202] = {9'd98,-10'd302};
ram[29203] = {-9'd99,-10'd299};
ram[29204] = {-9'd96,-10'd296};
ram[29205] = {-9'd92,-10'd293};
ram[29206] = {-9'd89,-10'd290};
ram[29207] = {-9'd86,-10'd286};
ram[29208] = {-9'd83,-10'd283};
ram[29209] = {-9'd80,-10'd280};
ram[29210] = {-9'd77,-10'd277};
ram[29211] = {-9'd74,-10'd274};
ram[29212] = {-9'd70,-10'd271};
ram[29213] = {-9'd67,-10'd268};
ram[29214] = {-9'd64,-10'd264};
ram[29215] = {-9'd61,-10'd261};
ram[29216] = {-9'd58,-10'd258};
ram[29217] = {-9'd55,-10'd255};
ram[29218] = {-9'd52,-10'd252};
ram[29219] = {-9'd48,-10'd249};
ram[29220] = {-9'd45,-10'd246};
ram[29221] = {-9'd42,-10'd242};
ram[29222] = {-9'd39,-10'd239};
ram[29223] = {-9'd36,-10'd236};
ram[29224] = {-9'd33,-10'd233};
ram[29225] = {-9'd30,-10'd230};
ram[29226] = {-9'd26,-10'd227};
ram[29227] = {-9'd23,-10'd224};
ram[29228] = {-9'd20,-10'd220};
ram[29229] = {-9'd17,-10'd217};
ram[29230] = {-9'd14,-10'd214};
ram[29231] = {-9'd11,-10'd211};
ram[29232] = {-9'd8,-10'd208};
ram[29233] = {-9'd4,-10'd205};
ram[29234] = {-9'd1,-10'd202};
ram[29235] = {9'd2,-10'd198};
ram[29236] = {9'd5,-10'd195};
ram[29237] = {9'd8,-10'd192};
ram[29238] = {9'd11,-10'd189};
ram[29239] = {9'd14,-10'd186};
ram[29240] = {9'd18,-10'd183};
ram[29241] = {9'd21,-10'd180};
ram[29242] = {9'd24,-10'd176};
ram[29243] = {9'd27,-10'd173};
ram[29244] = {9'd30,-10'd170};
ram[29245] = {9'd33,-10'd167};
ram[29246] = {9'd36,-10'd164};
ram[29247] = {9'd40,-10'd161};
ram[29248] = {9'd43,-10'd158};
ram[29249] = {9'd46,-10'd154};
ram[29250] = {9'd49,-10'd151};
ram[29251] = {9'd52,-10'd148};
ram[29252] = {9'd55,-10'd145};
ram[29253] = {9'd58,-10'd142};
ram[29254] = {9'd62,-10'd139};
ram[29255] = {9'd65,-10'd136};
ram[29256] = {9'd68,-10'd132};
ram[29257] = {9'd71,-10'd129};
ram[29258] = {9'd74,-10'd126};
ram[29259] = {9'd77,-10'd123};
ram[29260] = {9'd80,-10'd120};
ram[29261] = {9'd84,-10'd117};
ram[29262] = {9'd87,-10'd114};
ram[29263] = {9'd90,-10'd110};
ram[29264] = {9'd93,-10'd107};
ram[29265] = {9'd96,-10'd104};
ram[29266] = {9'd99,-10'd101};
ram[29267] = {-9'd98,-10'd98};
ram[29268] = {-9'd95,-10'd95};
ram[29269] = {-9'd92,-10'd92};
ram[29270] = {-9'd88,-10'd88};
ram[29271] = {-9'd85,-10'd85};
ram[29272] = {-9'd82,-10'd82};
ram[29273] = {-9'd79,-10'd79};
ram[29274] = {-9'd76,-10'd76};
ram[29275] = {-9'd73,-10'd73};
ram[29276] = {-9'd70,-10'd70};
ram[29277] = {-9'd66,-10'd66};
ram[29278] = {-9'd63,-10'd63};
ram[29279] = {-9'd60,-10'd60};
ram[29280] = {-9'd57,-10'd57};
ram[29281] = {-9'd54,-10'd54};
ram[29282] = {-9'd51,-10'd51};
ram[29283] = {-9'd48,-10'd48};
ram[29284] = {-9'd44,-10'd44};
ram[29285] = {-9'd41,-10'd41};
ram[29286] = {-9'd38,-10'd38};
ram[29287] = {-9'd35,-10'd35};
ram[29288] = {-9'd32,-10'd32};
ram[29289] = {-9'd29,-10'd29};
ram[29290] = {-9'd26,-10'd26};
ram[29291] = {-9'd22,-10'd22};
ram[29292] = {-9'd19,-10'd19};
ram[29293] = {-9'd16,-10'd16};
ram[29294] = {-9'd13,-10'd13};
ram[29295] = {-9'd10,-10'd10};
ram[29296] = {-9'd7,-10'd7};
ram[29297] = {-9'd4,-10'd4};
ram[29298] = {9'd0,10'd0};
ram[29299] = {9'd3,10'd3};
ram[29300] = {9'd6,10'd6};
ram[29301] = {9'd9,10'd9};
ram[29302] = {9'd12,10'd12};
ram[29303] = {9'd15,10'd15};
ram[29304] = {9'd18,10'd18};
ram[29305] = {9'd21,10'd21};
ram[29306] = {9'd25,10'd25};
ram[29307] = {9'd28,10'd28};
ram[29308] = {9'd31,10'd31};
ram[29309] = {9'd34,10'd34};
ram[29310] = {9'd37,10'd37};
ram[29311] = {9'd40,10'd40};
ram[29312] = {9'd40,10'd40};
ram[29313] = {9'd43,10'd43};
ram[29314] = {9'd47,10'd47};
ram[29315] = {9'd50,10'd50};
ram[29316] = {9'd53,10'd53};
ram[29317] = {9'd56,10'd56};
ram[29318] = {9'd59,10'd59};
ram[29319] = {9'd62,10'd62};
ram[29320] = {9'd65,10'd65};
ram[29321] = {9'd69,10'd69};
ram[29322] = {9'd72,10'd72};
ram[29323] = {9'd75,10'd75};
ram[29324] = {9'd78,10'd78};
ram[29325] = {9'd81,10'd81};
ram[29326] = {9'd84,10'd84};
ram[29327] = {9'd87,10'd87};
ram[29328] = {9'd91,10'd91};
ram[29329] = {9'd94,10'd94};
ram[29330] = {9'd97,10'd97};
ram[29331] = {-9'd100,10'd100};
ram[29332] = {-9'd97,10'd103};
ram[29333] = {-9'd94,10'd106};
ram[29334] = {-9'd91,10'd109};
ram[29335] = {-9'd88,10'd113};
ram[29336] = {-9'd85,10'd116};
ram[29337] = {-9'd81,10'd119};
ram[29338] = {-9'd78,10'd122};
ram[29339] = {-9'd75,10'd125};
ram[29340] = {-9'd72,10'd128};
ram[29341] = {-9'd69,10'd131};
ram[29342] = {-9'd66,10'd135};
ram[29343] = {-9'd63,10'd138};
ram[29344] = {-9'd59,10'd141};
ram[29345] = {-9'd56,10'd144};
ram[29346] = {-9'd53,10'd147};
ram[29347] = {-9'd50,10'd150};
ram[29348] = {-9'd47,10'd153};
ram[29349] = {-9'd44,10'd157};
ram[29350] = {-9'd41,10'd160};
ram[29351] = {-9'd37,10'd163};
ram[29352] = {-9'd34,10'd166};
ram[29353] = {-9'd31,10'd169};
ram[29354] = {-9'd28,10'd172};
ram[29355] = {-9'd25,10'd175};
ram[29356] = {-9'd22,10'd179};
ram[29357] = {-9'd19,10'd182};
ram[29358] = {-9'd15,10'd185};
ram[29359] = {-9'd12,10'd188};
ram[29360] = {-9'd9,10'd191};
ram[29361] = {-9'd6,10'd194};
ram[29362] = {-9'd3,10'd197};
ram[29363] = {9'd0,10'd201};
ram[29364] = {9'd3,10'd204};
ram[29365] = {9'd7,10'd207};
ram[29366] = {9'd10,10'd210};
ram[29367] = {9'd13,10'd213};
ram[29368] = {9'd16,10'd216};
ram[29369] = {9'd19,10'd219};
ram[29370] = {9'd22,10'd223};
ram[29371] = {9'd25,10'd226};
ram[29372] = {9'd29,10'd229};
ram[29373] = {9'd32,10'd232};
ram[29374] = {9'd35,10'd235};
ram[29375] = {9'd38,10'd238};
ram[29376] = {9'd41,10'd241};
ram[29377] = {9'd44,10'd245};
ram[29378] = {9'd47,10'd248};
ram[29379] = {9'd51,10'd251};
ram[29380] = {9'd54,10'd254};
ram[29381] = {9'd57,10'd257};
ram[29382] = {9'd60,10'd260};
ram[29383] = {9'd63,10'd263};
ram[29384] = {9'd66,10'd267};
ram[29385] = {9'd69,10'd270};
ram[29386] = {9'd73,10'd273};
ram[29387] = {9'd76,10'd276};
ram[29388] = {9'd79,10'd279};
ram[29389] = {9'd82,10'd282};
ram[29390] = {9'd85,10'd285};
ram[29391] = {9'd88,10'd289};
ram[29392] = {9'd91,10'd292};
ram[29393] = {9'd95,10'd295};
ram[29394] = {9'd98,10'd298};
ram[29395] = {-9'd99,10'd301};
ram[29396] = {-9'd96,10'd304};
ram[29397] = {-9'd93,10'd307};
ram[29398] = {-9'd90,10'd311};
ram[29399] = {-9'd87,10'd314};
ram[29400] = {-9'd84,10'd317};
ram[29401] = {-9'd81,10'd320};
ram[29402] = {-9'd77,10'd323};
ram[29403] = {-9'd74,10'd326};
ram[29404] = {-9'd71,10'd329};
ram[29405] = {-9'd68,10'd333};
ram[29406] = {-9'd65,10'd336};
ram[29407] = {-9'd62,10'd339};
ram[29408] = {-9'd59,10'd342};
ram[29409] = {-9'd55,10'd345};
ram[29410] = {-9'd52,10'd348};
ram[29411] = {-9'd49,10'd351};
ram[29412] = {-9'd46,10'd354};
ram[29413] = {-9'd43,10'd358};
ram[29414] = {-9'd40,10'd361};
ram[29415] = {-9'd37,10'd364};
ram[29416] = {-9'd33,10'd367};
ram[29417] = {-9'd30,10'd370};
ram[29418] = {-9'd27,10'd373};
ram[29419] = {-9'd24,10'd376};
ram[29420] = {-9'd21,10'd380};
ram[29421] = {-9'd18,10'd383};
ram[29422] = {-9'd15,10'd386};
ram[29423] = {-9'd11,10'd389};
ram[29424] = {-9'd8,10'd392};
ram[29425] = {-9'd5,10'd395};
ram[29426] = {-9'd2,10'd398};
ram[29427] = {9'd1,-10'd399};
ram[29428] = {9'd4,-10'd396};
ram[29429] = {9'd7,-10'd393};
ram[29430] = {9'd10,-10'd390};
ram[29431] = {9'd14,-10'd387};
ram[29432] = {9'd17,-10'd384};
ram[29433] = {9'd20,-10'd381};
ram[29434] = {9'd23,-10'd377};
ram[29435] = {9'd26,-10'd374};
ram[29436] = {9'd29,-10'd371};
ram[29437] = {9'd32,-10'd368};
ram[29438] = {9'd36,-10'd365};
ram[29439] = {9'd39,-10'd362};
ram[29440] = {9'd39,-10'd362};
ram[29441] = {9'd42,-10'd359};
ram[29442] = {9'd45,-10'd355};
ram[29443] = {9'd48,-10'd352};
ram[29444] = {9'd51,-10'd349};
ram[29445] = {9'd54,-10'd346};
ram[29446] = {9'd58,-10'd343};
ram[29447] = {9'd61,-10'd340};
ram[29448] = {9'd64,-10'd337};
ram[29449] = {9'd67,-10'd334};
ram[29450] = {9'd70,-10'd330};
ram[29451] = {9'd73,-10'd327};
ram[29452] = {9'd76,-10'd324};
ram[29453] = {9'd80,-10'd321};
ram[29454] = {9'd83,-10'd318};
ram[29455] = {9'd86,-10'd315};
ram[29456] = {9'd89,-10'd312};
ram[29457] = {9'd92,-10'd308};
ram[29458] = {9'd95,-10'd305};
ram[29459] = {9'd98,-10'd302};
ram[29460] = {-9'd99,-10'd299};
ram[29461] = {-9'd96,-10'd296};
ram[29462] = {-9'd92,-10'd293};
ram[29463] = {-9'd89,-10'd290};
ram[29464] = {-9'd86,-10'd286};
ram[29465] = {-9'd83,-10'd283};
ram[29466] = {-9'd80,-10'd280};
ram[29467] = {-9'd77,-10'd277};
ram[29468] = {-9'd74,-10'd274};
ram[29469] = {-9'd70,-10'd271};
ram[29470] = {-9'd67,-10'd268};
ram[29471] = {-9'd64,-10'd264};
ram[29472] = {-9'd61,-10'd261};
ram[29473] = {-9'd58,-10'd258};
ram[29474] = {-9'd55,-10'd255};
ram[29475] = {-9'd52,-10'd252};
ram[29476] = {-9'd48,-10'd249};
ram[29477] = {-9'd45,-10'd246};
ram[29478] = {-9'd42,-10'd242};
ram[29479] = {-9'd39,-10'd239};
ram[29480] = {-9'd36,-10'd236};
ram[29481] = {-9'd33,-10'd233};
ram[29482] = {-9'd30,-10'd230};
ram[29483] = {-9'd26,-10'd227};
ram[29484] = {-9'd23,-10'd224};
ram[29485] = {-9'd20,-10'd220};
ram[29486] = {-9'd17,-10'd217};
ram[29487] = {-9'd14,-10'd214};
ram[29488] = {-9'd11,-10'd211};
ram[29489] = {-9'd8,-10'd208};
ram[29490] = {-9'd4,-10'd205};
ram[29491] = {-9'd1,-10'd202};
ram[29492] = {9'd2,-10'd198};
ram[29493] = {9'd5,-10'd195};
ram[29494] = {9'd8,-10'd192};
ram[29495] = {9'd11,-10'd189};
ram[29496] = {9'd14,-10'd186};
ram[29497] = {9'd18,-10'd183};
ram[29498] = {9'd21,-10'd180};
ram[29499] = {9'd24,-10'd176};
ram[29500] = {9'd27,-10'd173};
ram[29501] = {9'd30,-10'd170};
ram[29502] = {9'd33,-10'd167};
ram[29503] = {9'd36,-10'd164};
ram[29504] = {9'd40,-10'd161};
ram[29505] = {9'd43,-10'd158};
ram[29506] = {9'd46,-10'd154};
ram[29507] = {9'd49,-10'd151};
ram[29508] = {9'd52,-10'd148};
ram[29509] = {9'd55,-10'd145};
ram[29510] = {9'd58,-10'd142};
ram[29511] = {9'd62,-10'd139};
ram[29512] = {9'd65,-10'd136};
ram[29513] = {9'd68,-10'd132};
ram[29514] = {9'd71,-10'd129};
ram[29515] = {9'd74,-10'd126};
ram[29516] = {9'd77,-10'd123};
ram[29517] = {9'd80,-10'd120};
ram[29518] = {9'd84,-10'd117};
ram[29519] = {9'd87,-10'd114};
ram[29520] = {9'd90,-10'd110};
ram[29521] = {9'd93,-10'd107};
ram[29522] = {9'd96,-10'd104};
ram[29523] = {9'd99,-10'd101};
ram[29524] = {-9'd98,-10'd98};
ram[29525] = {-9'd95,-10'd95};
ram[29526] = {-9'd92,-10'd92};
ram[29527] = {-9'd88,-10'd88};
ram[29528] = {-9'd85,-10'd85};
ram[29529] = {-9'd82,-10'd82};
ram[29530] = {-9'd79,-10'd79};
ram[29531] = {-9'd76,-10'd76};
ram[29532] = {-9'd73,-10'd73};
ram[29533] = {-9'd70,-10'd70};
ram[29534] = {-9'd66,-10'd66};
ram[29535] = {-9'd63,-10'd63};
ram[29536] = {-9'd60,-10'd60};
ram[29537] = {-9'd57,-10'd57};
ram[29538] = {-9'd54,-10'd54};
ram[29539] = {-9'd51,-10'd51};
ram[29540] = {-9'd48,-10'd48};
ram[29541] = {-9'd44,-10'd44};
ram[29542] = {-9'd41,-10'd41};
ram[29543] = {-9'd38,-10'd38};
ram[29544] = {-9'd35,-10'd35};
ram[29545] = {-9'd32,-10'd32};
ram[29546] = {-9'd29,-10'd29};
ram[29547] = {-9'd26,-10'd26};
ram[29548] = {-9'd22,-10'd22};
ram[29549] = {-9'd19,-10'd19};
ram[29550] = {-9'd16,-10'd16};
ram[29551] = {-9'd13,-10'd13};
ram[29552] = {-9'd10,-10'd10};
ram[29553] = {-9'd7,-10'd7};
ram[29554] = {-9'd4,-10'd4};
ram[29555] = {9'd0,10'd0};
ram[29556] = {9'd3,10'd3};
ram[29557] = {9'd6,10'd6};
ram[29558] = {9'd9,10'd9};
ram[29559] = {9'd12,10'd12};
ram[29560] = {9'd15,10'd15};
ram[29561] = {9'd18,10'd18};
ram[29562] = {9'd21,10'd21};
ram[29563] = {9'd25,10'd25};
ram[29564] = {9'd28,10'd28};
ram[29565] = {9'd31,10'd31};
ram[29566] = {9'd34,10'd34};
ram[29567] = {9'd37,10'd37};
ram[29568] = {9'd37,10'd37};
ram[29569] = {9'd40,10'd40};
ram[29570] = {9'd43,10'd43};
ram[29571] = {9'd47,10'd47};
ram[29572] = {9'd50,10'd50};
ram[29573] = {9'd53,10'd53};
ram[29574] = {9'd56,10'd56};
ram[29575] = {9'd59,10'd59};
ram[29576] = {9'd62,10'd62};
ram[29577] = {9'd65,10'd65};
ram[29578] = {9'd69,10'd69};
ram[29579] = {9'd72,10'd72};
ram[29580] = {9'd75,10'd75};
ram[29581] = {9'd78,10'd78};
ram[29582] = {9'd81,10'd81};
ram[29583] = {9'd84,10'd84};
ram[29584] = {9'd87,10'd87};
ram[29585] = {9'd91,10'd91};
ram[29586] = {9'd94,10'd94};
ram[29587] = {9'd97,10'd97};
ram[29588] = {-9'd100,10'd100};
ram[29589] = {-9'd97,10'd103};
ram[29590] = {-9'd94,10'd106};
ram[29591] = {-9'd91,10'd109};
ram[29592] = {-9'd88,10'd113};
ram[29593] = {-9'd85,10'd116};
ram[29594] = {-9'd81,10'd119};
ram[29595] = {-9'd78,10'd122};
ram[29596] = {-9'd75,10'd125};
ram[29597] = {-9'd72,10'd128};
ram[29598] = {-9'd69,10'd131};
ram[29599] = {-9'd66,10'd135};
ram[29600] = {-9'd63,10'd138};
ram[29601] = {-9'd59,10'd141};
ram[29602] = {-9'd56,10'd144};
ram[29603] = {-9'd53,10'd147};
ram[29604] = {-9'd50,10'd150};
ram[29605] = {-9'd47,10'd153};
ram[29606] = {-9'd44,10'd157};
ram[29607] = {-9'd41,10'd160};
ram[29608] = {-9'd37,10'd163};
ram[29609] = {-9'd34,10'd166};
ram[29610] = {-9'd31,10'd169};
ram[29611] = {-9'd28,10'd172};
ram[29612] = {-9'd25,10'd175};
ram[29613] = {-9'd22,10'd179};
ram[29614] = {-9'd19,10'd182};
ram[29615] = {-9'd15,10'd185};
ram[29616] = {-9'd12,10'd188};
ram[29617] = {-9'd9,10'd191};
ram[29618] = {-9'd6,10'd194};
ram[29619] = {-9'd3,10'd197};
ram[29620] = {9'd0,10'd201};
ram[29621] = {9'd3,10'd204};
ram[29622] = {9'd7,10'd207};
ram[29623] = {9'd10,10'd210};
ram[29624] = {9'd13,10'd213};
ram[29625] = {9'd16,10'd216};
ram[29626] = {9'd19,10'd219};
ram[29627] = {9'd22,10'd223};
ram[29628] = {9'd25,10'd226};
ram[29629] = {9'd29,10'd229};
ram[29630] = {9'd32,10'd232};
ram[29631] = {9'd35,10'd235};
ram[29632] = {9'd38,10'd238};
ram[29633] = {9'd41,10'd241};
ram[29634] = {9'd44,10'd245};
ram[29635] = {9'd47,10'd248};
ram[29636] = {9'd51,10'd251};
ram[29637] = {9'd54,10'd254};
ram[29638] = {9'd57,10'd257};
ram[29639] = {9'd60,10'd260};
ram[29640] = {9'd63,10'd263};
ram[29641] = {9'd66,10'd267};
ram[29642] = {9'd69,10'd270};
ram[29643] = {9'd73,10'd273};
ram[29644] = {9'd76,10'd276};
ram[29645] = {9'd79,10'd279};
ram[29646] = {9'd82,10'd282};
ram[29647] = {9'd85,10'd285};
ram[29648] = {9'd88,10'd289};
ram[29649] = {9'd91,10'd292};
ram[29650] = {9'd95,10'd295};
ram[29651] = {9'd98,10'd298};
ram[29652] = {-9'd99,10'd301};
ram[29653] = {-9'd96,10'd304};
ram[29654] = {-9'd93,10'd307};
ram[29655] = {-9'd90,10'd311};
ram[29656] = {-9'd87,10'd314};
ram[29657] = {-9'd84,10'd317};
ram[29658] = {-9'd81,10'd320};
ram[29659] = {-9'd77,10'd323};
ram[29660] = {-9'd74,10'd326};
ram[29661] = {-9'd71,10'd329};
ram[29662] = {-9'd68,10'd333};
ram[29663] = {-9'd65,10'd336};
ram[29664] = {-9'd62,10'd339};
ram[29665] = {-9'd59,10'd342};
ram[29666] = {-9'd55,10'd345};
ram[29667] = {-9'd52,10'd348};
ram[29668] = {-9'd49,10'd351};
ram[29669] = {-9'd46,10'd354};
ram[29670] = {-9'd43,10'd358};
ram[29671] = {-9'd40,10'd361};
ram[29672] = {-9'd37,10'd364};
ram[29673] = {-9'd33,10'd367};
ram[29674] = {-9'd30,10'd370};
ram[29675] = {-9'd27,10'd373};
ram[29676] = {-9'd24,10'd376};
ram[29677] = {-9'd21,10'd380};
ram[29678] = {-9'd18,10'd383};
ram[29679] = {-9'd15,10'd386};
ram[29680] = {-9'd11,10'd389};
ram[29681] = {-9'd8,10'd392};
ram[29682] = {-9'd5,10'd395};
ram[29683] = {-9'd2,10'd398};
ram[29684] = {9'd1,-10'd399};
ram[29685] = {9'd4,-10'd396};
ram[29686] = {9'd7,-10'd393};
ram[29687] = {9'd10,-10'd390};
ram[29688] = {9'd14,-10'd387};
ram[29689] = {9'd17,-10'd384};
ram[29690] = {9'd20,-10'd381};
ram[29691] = {9'd23,-10'd377};
ram[29692] = {9'd26,-10'd374};
ram[29693] = {9'd29,-10'd371};
ram[29694] = {9'd32,-10'd368};
ram[29695] = {9'd36,-10'd365};
ram[29696] = {9'd36,-10'd365};
ram[29697] = {9'd39,-10'd362};
ram[29698] = {9'd42,-10'd359};
ram[29699] = {9'd45,-10'd355};
ram[29700] = {9'd48,-10'd352};
ram[29701] = {9'd51,-10'd349};
ram[29702] = {9'd54,-10'd346};
ram[29703] = {9'd58,-10'd343};
ram[29704] = {9'd61,-10'd340};
ram[29705] = {9'd64,-10'd337};
ram[29706] = {9'd67,-10'd334};
ram[29707] = {9'd70,-10'd330};
ram[29708] = {9'd73,-10'd327};
ram[29709] = {9'd76,-10'd324};
ram[29710] = {9'd80,-10'd321};
ram[29711] = {9'd83,-10'd318};
ram[29712] = {9'd86,-10'd315};
ram[29713] = {9'd89,-10'd312};
ram[29714] = {9'd92,-10'd308};
ram[29715] = {9'd95,-10'd305};
ram[29716] = {9'd98,-10'd302};
ram[29717] = {-9'd99,-10'd299};
ram[29718] = {-9'd96,-10'd296};
ram[29719] = {-9'd92,-10'd293};
ram[29720] = {-9'd89,-10'd290};
ram[29721] = {-9'd86,-10'd286};
ram[29722] = {-9'd83,-10'd283};
ram[29723] = {-9'd80,-10'd280};
ram[29724] = {-9'd77,-10'd277};
ram[29725] = {-9'd74,-10'd274};
ram[29726] = {-9'd70,-10'd271};
ram[29727] = {-9'd67,-10'd268};
ram[29728] = {-9'd64,-10'd264};
ram[29729] = {-9'd61,-10'd261};
ram[29730] = {-9'd58,-10'd258};
ram[29731] = {-9'd55,-10'd255};
ram[29732] = {-9'd52,-10'd252};
ram[29733] = {-9'd48,-10'd249};
ram[29734] = {-9'd45,-10'd246};
ram[29735] = {-9'd42,-10'd242};
ram[29736] = {-9'd39,-10'd239};
ram[29737] = {-9'd36,-10'd236};
ram[29738] = {-9'd33,-10'd233};
ram[29739] = {-9'd30,-10'd230};
ram[29740] = {-9'd26,-10'd227};
ram[29741] = {-9'd23,-10'd224};
ram[29742] = {-9'd20,-10'd220};
ram[29743] = {-9'd17,-10'd217};
ram[29744] = {-9'd14,-10'd214};
ram[29745] = {-9'd11,-10'd211};
ram[29746] = {-9'd8,-10'd208};
ram[29747] = {-9'd4,-10'd205};
ram[29748] = {-9'd1,-10'd202};
ram[29749] = {9'd2,-10'd198};
ram[29750] = {9'd5,-10'd195};
ram[29751] = {9'd8,-10'd192};
ram[29752] = {9'd11,-10'd189};
ram[29753] = {9'd14,-10'd186};
ram[29754] = {9'd18,-10'd183};
ram[29755] = {9'd21,-10'd180};
ram[29756] = {9'd24,-10'd176};
ram[29757] = {9'd27,-10'd173};
ram[29758] = {9'd30,-10'd170};
ram[29759] = {9'd33,-10'd167};
ram[29760] = {9'd36,-10'd164};
ram[29761] = {9'd40,-10'd161};
ram[29762] = {9'd43,-10'd158};
ram[29763] = {9'd46,-10'd154};
ram[29764] = {9'd49,-10'd151};
ram[29765] = {9'd52,-10'd148};
ram[29766] = {9'd55,-10'd145};
ram[29767] = {9'd58,-10'd142};
ram[29768] = {9'd62,-10'd139};
ram[29769] = {9'd65,-10'd136};
ram[29770] = {9'd68,-10'd132};
ram[29771] = {9'd71,-10'd129};
ram[29772] = {9'd74,-10'd126};
ram[29773] = {9'd77,-10'd123};
ram[29774] = {9'd80,-10'd120};
ram[29775] = {9'd84,-10'd117};
ram[29776] = {9'd87,-10'd114};
ram[29777] = {9'd90,-10'd110};
ram[29778] = {9'd93,-10'd107};
ram[29779] = {9'd96,-10'd104};
ram[29780] = {9'd99,-10'd101};
ram[29781] = {-9'd98,-10'd98};
ram[29782] = {-9'd95,-10'd95};
ram[29783] = {-9'd92,-10'd92};
ram[29784] = {-9'd88,-10'd88};
ram[29785] = {-9'd85,-10'd85};
ram[29786] = {-9'd82,-10'd82};
ram[29787] = {-9'd79,-10'd79};
ram[29788] = {-9'd76,-10'd76};
ram[29789] = {-9'd73,-10'd73};
ram[29790] = {-9'd70,-10'd70};
ram[29791] = {-9'd66,-10'd66};
ram[29792] = {-9'd63,-10'd63};
ram[29793] = {-9'd60,-10'd60};
ram[29794] = {-9'd57,-10'd57};
ram[29795] = {-9'd54,-10'd54};
ram[29796] = {-9'd51,-10'd51};
ram[29797] = {-9'd48,-10'd48};
ram[29798] = {-9'd44,-10'd44};
ram[29799] = {-9'd41,-10'd41};
ram[29800] = {-9'd38,-10'd38};
ram[29801] = {-9'd35,-10'd35};
ram[29802] = {-9'd32,-10'd32};
ram[29803] = {-9'd29,-10'd29};
ram[29804] = {-9'd26,-10'd26};
ram[29805] = {-9'd22,-10'd22};
ram[29806] = {-9'd19,-10'd19};
ram[29807] = {-9'd16,-10'd16};
ram[29808] = {-9'd13,-10'd13};
ram[29809] = {-9'd10,-10'd10};
ram[29810] = {-9'd7,-10'd7};
ram[29811] = {-9'd4,-10'd4};
ram[29812] = {9'd0,10'd0};
ram[29813] = {9'd3,10'd3};
ram[29814] = {9'd6,10'd6};
ram[29815] = {9'd9,10'd9};
ram[29816] = {9'd12,10'd12};
ram[29817] = {9'd15,10'd15};
ram[29818] = {9'd18,10'd18};
ram[29819] = {9'd21,10'd21};
ram[29820] = {9'd25,10'd25};
ram[29821] = {9'd28,10'd28};
ram[29822] = {9'd31,10'd31};
ram[29823] = {9'd34,10'd34};
ram[29824] = {9'd34,10'd34};
ram[29825] = {9'd37,10'd37};
ram[29826] = {9'd40,10'd40};
ram[29827] = {9'd43,10'd43};
ram[29828] = {9'd47,10'd47};
ram[29829] = {9'd50,10'd50};
ram[29830] = {9'd53,10'd53};
ram[29831] = {9'd56,10'd56};
ram[29832] = {9'd59,10'd59};
ram[29833] = {9'd62,10'd62};
ram[29834] = {9'd65,10'd65};
ram[29835] = {9'd69,10'd69};
ram[29836] = {9'd72,10'd72};
ram[29837] = {9'd75,10'd75};
ram[29838] = {9'd78,10'd78};
ram[29839] = {9'd81,10'd81};
ram[29840] = {9'd84,10'd84};
ram[29841] = {9'd87,10'd87};
ram[29842] = {9'd91,10'd91};
ram[29843] = {9'd94,10'd94};
ram[29844] = {9'd97,10'd97};
ram[29845] = {-9'd100,10'd100};
ram[29846] = {-9'd97,10'd103};
ram[29847] = {-9'd94,10'd106};
ram[29848] = {-9'd91,10'd109};
ram[29849] = {-9'd88,10'd113};
ram[29850] = {-9'd85,10'd116};
ram[29851] = {-9'd81,10'd119};
ram[29852] = {-9'd78,10'd122};
ram[29853] = {-9'd75,10'd125};
ram[29854] = {-9'd72,10'd128};
ram[29855] = {-9'd69,10'd131};
ram[29856] = {-9'd66,10'd135};
ram[29857] = {-9'd63,10'd138};
ram[29858] = {-9'd59,10'd141};
ram[29859] = {-9'd56,10'd144};
ram[29860] = {-9'd53,10'd147};
ram[29861] = {-9'd50,10'd150};
ram[29862] = {-9'd47,10'd153};
ram[29863] = {-9'd44,10'd157};
ram[29864] = {-9'd41,10'd160};
ram[29865] = {-9'd37,10'd163};
ram[29866] = {-9'd34,10'd166};
ram[29867] = {-9'd31,10'd169};
ram[29868] = {-9'd28,10'd172};
ram[29869] = {-9'd25,10'd175};
ram[29870] = {-9'd22,10'd179};
ram[29871] = {-9'd19,10'd182};
ram[29872] = {-9'd15,10'd185};
ram[29873] = {-9'd12,10'd188};
ram[29874] = {-9'd9,10'd191};
ram[29875] = {-9'd6,10'd194};
ram[29876] = {-9'd3,10'd197};
ram[29877] = {9'd0,10'd201};
ram[29878] = {9'd3,10'd204};
ram[29879] = {9'd7,10'd207};
ram[29880] = {9'd10,10'd210};
ram[29881] = {9'd13,10'd213};
ram[29882] = {9'd16,10'd216};
ram[29883] = {9'd19,10'd219};
ram[29884] = {9'd22,10'd223};
ram[29885] = {9'd25,10'd226};
ram[29886] = {9'd29,10'd229};
ram[29887] = {9'd32,10'd232};
ram[29888] = {9'd35,10'd235};
ram[29889] = {9'd38,10'd238};
ram[29890] = {9'd41,10'd241};
ram[29891] = {9'd44,10'd245};
ram[29892] = {9'd47,10'd248};
ram[29893] = {9'd51,10'd251};
ram[29894] = {9'd54,10'd254};
ram[29895] = {9'd57,10'd257};
ram[29896] = {9'd60,10'd260};
ram[29897] = {9'd63,10'd263};
ram[29898] = {9'd66,10'd267};
ram[29899] = {9'd69,10'd270};
ram[29900] = {9'd73,10'd273};
ram[29901] = {9'd76,10'd276};
ram[29902] = {9'd79,10'd279};
ram[29903] = {9'd82,10'd282};
ram[29904] = {9'd85,10'd285};
ram[29905] = {9'd88,10'd289};
ram[29906] = {9'd91,10'd292};
ram[29907] = {9'd95,10'd295};
ram[29908] = {9'd98,10'd298};
ram[29909] = {-9'd99,10'd301};
ram[29910] = {-9'd96,10'd304};
ram[29911] = {-9'd93,10'd307};
ram[29912] = {-9'd90,10'd311};
ram[29913] = {-9'd87,10'd314};
ram[29914] = {-9'd84,10'd317};
ram[29915] = {-9'd81,10'd320};
ram[29916] = {-9'd77,10'd323};
ram[29917] = {-9'd74,10'd326};
ram[29918] = {-9'd71,10'd329};
ram[29919] = {-9'd68,10'd333};
ram[29920] = {-9'd65,10'd336};
ram[29921] = {-9'd62,10'd339};
ram[29922] = {-9'd59,10'd342};
ram[29923] = {-9'd55,10'd345};
ram[29924] = {-9'd52,10'd348};
ram[29925] = {-9'd49,10'd351};
ram[29926] = {-9'd46,10'd354};
ram[29927] = {-9'd43,10'd358};
ram[29928] = {-9'd40,10'd361};
ram[29929] = {-9'd37,10'd364};
ram[29930] = {-9'd33,10'd367};
ram[29931] = {-9'd30,10'd370};
ram[29932] = {-9'd27,10'd373};
ram[29933] = {-9'd24,10'd376};
ram[29934] = {-9'd21,10'd380};
ram[29935] = {-9'd18,10'd383};
ram[29936] = {-9'd15,10'd386};
ram[29937] = {-9'd11,10'd389};
ram[29938] = {-9'd8,10'd392};
ram[29939] = {-9'd5,10'd395};
ram[29940] = {-9'd2,10'd398};
ram[29941] = {9'd1,-10'd399};
ram[29942] = {9'd4,-10'd396};
ram[29943] = {9'd7,-10'd393};
ram[29944] = {9'd10,-10'd390};
ram[29945] = {9'd14,-10'd387};
ram[29946] = {9'd17,-10'd384};
ram[29947] = {9'd20,-10'd381};
ram[29948] = {9'd23,-10'd377};
ram[29949] = {9'd26,-10'd374};
ram[29950] = {9'd29,-10'd371};
ram[29951] = {9'd32,-10'd368};
ram[29952] = {9'd32,-10'd368};
ram[29953] = {9'd36,-10'd365};
ram[29954] = {9'd39,-10'd362};
ram[29955] = {9'd42,-10'd359};
ram[29956] = {9'd45,-10'd355};
ram[29957] = {9'd48,-10'd352};
ram[29958] = {9'd51,-10'd349};
ram[29959] = {9'd54,-10'd346};
ram[29960] = {9'd58,-10'd343};
ram[29961] = {9'd61,-10'd340};
ram[29962] = {9'd64,-10'd337};
ram[29963] = {9'd67,-10'd334};
ram[29964] = {9'd70,-10'd330};
ram[29965] = {9'd73,-10'd327};
ram[29966] = {9'd76,-10'd324};
ram[29967] = {9'd80,-10'd321};
ram[29968] = {9'd83,-10'd318};
ram[29969] = {9'd86,-10'd315};
ram[29970] = {9'd89,-10'd312};
ram[29971] = {9'd92,-10'd308};
ram[29972] = {9'd95,-10'd305};
ram[29973] = {9'd98,-10'd302};
ram[29974] = {-9'd99,-10'd299};
ram[29975] = {-9'd96,-10'd296};
ram[29976] = {-9'd92,-10'd293};
ram[29977] = {-9'd89,-10'd290};
ram[29978] = {-9'd86,-10'd286};
ram[29979] = {-9'd83,-10'd283};
ram[29980] = {-9'd80,-10'd280};
ram[29981] = {-9'd77,-10'd277};
ram[29982] = {-9'd74,-10'd274};
ram[29983] = {-9'd70,-10'd271};
ram[29984] = {-9'd67,-10'd268};
ram[29985] = {-9'd64,-10'd264};
ram[29986] = {-9'd61,-10'd261};
ram[29987] = {-9'd58,-10'd258};
ram[29988] = {-9'd55,-10'd255};
ram[29989] = {-9'd52,-10'd252};
ram[29990] = {-9'd48,-10'd249};
ram[29991] = {-9'd45,-10'd246};
ram[29992] = {-9'd42,-10'd242};
ram[29993] = {-9'd39,-10'd239};
ram[29994] = {-9'd36,-10'd236};
ram[29995] = {-9'd33,-10'd233};
ram[29996] = {-9'd30,-10'd230};
ram[29997] = {-9'd26,-10'd227};
ram[29998] = {-9'd23,-10'd224};
ram[29999] = {-9'd20,-10'd220};
ram[30000] = {-9'd17,-10'd217};
ram[30001] = {-9'd14,-10'd214};
ram[30002] = {-9'd11,-10'd211};
ram[30003] = {-9'd8,-10'd208};
ram[30004] = {-9'd4,-10'd205};
ram[30005] = {-9'd1,-10'd202};
ram[30006] = {9'd2,-10'd198};
ram[30007] = {9'd5,-10'd195};
ram[30008] = {9'd8,-10'd192};
ram[30009] = {9'd11,-10'd189};
ram[30010] = {9'd14,-10'd186};
ram[30011] = {9'd18,-10'd183};
ram[30012] = {9'd21,-10'd180};
ram[30013] = {9'd24,-10'd176};
ram[30014] = {9'd27,-10'd173};
ram[30015] = {9'd30,-10'd170};
ram[30016] = {9'd33,-10'd167};
ram[30017] = {9'd36,-10'd164};
ram[30018] = {9'd40,-10'd161};
ram[30019] = {9'd43,-10'd158};
ram[30020] = {9'd46,-10'd154};
ram[30021] = {9'd49,-10'd151};
ram[30022] = {9'd52,-10'd148};
ram[30023] = {9'd55,-10'd145};
ram[30024] = {9'd58,-10'd142};
ram[30025] = {9'd62,-10'd139};
ram[30026] = {9'd65,-10'd136};
ram[30027] = {9'd68,-10'd132};
ram[30028] = {9'd71,-10'd129};
ram[30029] = {9'd74,-10'd126};
ram[30030] = {9'd77,-10'd123};
ram[30031] = {9'd80,-10'd120};
ram[30032] = {9'd84,-10'd117};
ram[30033] = {9'd87,-10'd114};
ram[30034] = {9'd90,-10'd110};
ram[30035] = {9'd93,-10'd107};
ram[30036] = {9'd96,-10'd104};
ram[30037] = {9'd99,-10'd101};
ram[30038] = {-9'd98,-10'd98};
ram[30039] = {-9'd95,-10'd95};
ram[30040] = {-9'd92,-10'd92};
ram[30041] = {-9'd88,-10'd88};
ram[30042] = {-9'd85,-10'd85};
ram[30043] = {-9'd82,-10'd82};
ram[30044] = {-9'd79,-10'd79};
ram[30045] = {-9'd76,-10'd76};
ram[30046] = {-9'd73,-10'd73};
ram[30047] = {-9'd70,-10'd70};
ram[30048] = {-9'd66,-10'd66};
ram[30049] = {-9'd63,-10'd63};
ram[30050] = {-9'd60,-10'd60};
ram[30051] = {-9'd57,-10'd57};
ram[30052] = {-9'd54,-10'd54};
ram[30053] = {-9'd51,-10'd51};
ram[30054] = {-9'd48,-10'd48};
ram[30055] = {-9'd44,-10'd44};
ram[30056] = {-9'd41,-10'd41};
ram[30057] = {-9'd38,-10'd38};
ram[30058] = {-9'd35,-10'd35};
ram[30059] = {-9'd32,-10'd32};
ram[30060] = {-9'd29,-10'd29};
ram[30061] = {-9'd26,-10'd26};
ram[30062] = {-9'd22,-10'd22};
ram[30063] = {-9'd19,-10'd19};
ram[30064] = {-9'd16,-10'd16};
ram[30065] = {-9'd13,-10'd13};
ram[30066] = {-9'd10,-10'd10};
ram[30067] = {-9'd7,-10'd7};
ram[30068] = {-9'd4,-10'd4};
ram[30069] = {9'd0,10'd0};
ram[30070] = {9'd3,10'd3};
ram[30071] = {9'd6,10'd6};
ram[30072] = {9'd9,10'd9};
ram[30073] = {9'd12,10'd12};
ram[30074] = {9'd15,10'd15};
ram[30075] = {9'd18,10'd18};
ram[30076] = {9'd21,10'd21};
ram[30077] = {9'd25,10'd25};
ram[30078] = {9'd28,10'd28};
ram[30079] = {9'd31,10'd31};
ram[30080] = {9'd31,10'd31};
ram[30081] = {9'd34,10'd34};
ram[30082] = {9'd37,10'd37};
ram[30083] = {9'd40,10'd40};
ram[30084] = {9'd43,10'd43};
ram[30085] = {9'd47,10'd47};
ram[30086] = {9'd50,10'd50};
ram[30087] = {9'd53,10'd53};
ram[30088] = {9'd56,10'd56};
ram[30089] = {9'd59,10'd59};
ram[30090] = {9'd62,10'd62};
ram[30091] = {9'd65,10'd65};
ram[30092] = {9'd69,10'd69};
ram[30093] = {9'd72,10'd72};
ram[30094] = {9'd75,10'd75};
ram[30095] = {9'd78,10'd78};
ram[30096] = {9'd81,10'd81};
ram[30097] = {9'd84,10'd84};
ram[30098] = {9'd87,10'd87};
ram[30099] = {9'd91,10'd91};
ram[30100] = {9'd94,10'd94};
ram[30101] = {9'd97,10'd97};
ram[30102] = {-9'd100,10'd100};
ram[30103] = {-9'd97,10'd103};
ram[30104] = {-9'd94,10'd106};
ram[30105] = {-9'd91,10'd109};
ram[30106] = {-9'd88,10'd113};
ram[30107] = {-9'd85,10'd116};
ram[30108] = {-9'd81,10'd119};
ram[30109] = {-9'd78,10'd122};
ram[30110] = {-9'd75,10'd125};
ram[30111] = {-9'd72,10'd128};
ram[30112] = {-9'd69,10'd131};
ram[30113] = {-9'd66,10'd135};
ram[30114] = {-9'd63,10'd138};
ram[30115] = {-9'd59,10'd141};
ram[30116] = {-9'd56,10'd144};
ram[30117] = {-9'd53,10'd147};
ram[30118] = {-9'd50,10'd150};
ram[30119] = {-9'd47,10'd153};
ram[30120] = {-9'd44,10'd157};
ram[30121] = {-9'd41,10'd160};
ram[30122] = {-9'd37,10'd163};
ram[30123] = {-9'd34,10'd166};
ram[30124] = {-9'd31,10'd169};
ram[30125] = {-9'd28,10'd172};
ram[30126] = {-9'd25,10'd175};
ram[30127] = {-9'd22,10'd179};
ram[30128] = {-9'd19,10'd182};
ram[30129] = {-9'd15,10'd185};
ram[30130] = {-9'd12,10'd188};
ram[30131] = {-9'd9,10'd191};
ram[30132] = {-9'd6,10'd194};
ram[30133] = {-9'd3,10'd197};
ram[30134] = {9'd0,10'd201};
ram[30135] = {9'd3,10'd204};
ram[30136] = {9'd7,10'd207};
ram[30137] = {9'd10,10'd210};
ram[30138] = {9'd13,10'd213};
ram[30139] = {9'd16,10'd216};
ram[30140] = {9'd19,10'd219};
ram[30141] = {9'd22,10'd223};
ram[30142] = {9'd25,10'd226};
ram[30143] = {9'd29,10'd229};
ram[30144] = {9'd32,10'd232};
ram[30145] = {9'd35,10'd235};
ram[30146] = {9'd38,10'd238};
ram[30147] = {9'd41,10'd241};
ram[30148] = {9'd44,10'd245};
ram[30149] = {9'd47,10'd248};
ram[30150] = {9'd51,10'd251};
ram[30151] = {9'd54,10'd254};
ram[30152] = {9'd57,10'd257};
ram[30153] = {9'd60,10'd260};
ram[30154] = {9'd63,10'd263};
ram[30155] = {9'd66,10'd267};
ram[30156] = {9'd69,10'd270};
ram[30157] = {9'd73,10'd273};
ram[30158] = {9'd76,10'd276};
ram[30159] = {9'd79,10'd279};
ram[30160] = {9'd82,10'd282};
ram[30161] = {9'd85,10'd285};
ram[30162] = {9'd88,10'd289};
ram[30163] = {9'd91,10'd292};
ram[30164] = {9'd95,10'd295};
ram[30165] = {9'd98,10'd298};
ram[30166] = {-9'd99,10'd301};
ram[30167] = {-9'd96,10'd304};
ram[30168] = {-9'd93,10'd307};
ram[30169] = {-9'd90,10'd311};
ram[30170] = {-9'd87,10'd314};
ram[30171] = {-9'd84,10'd317};
ram[30172] = {-9'd81,10'd320};
ram[30173] = {-9'd77,10'd323};
ram[30174] = {-9'd74,10'd326};
ram[30175] = {-9'd71,10'd329};
ram[30176] = {-9'd68,10'd333};
ram[30177] = {-9'd65,10'd336};
ram[30178] = {-9'd62,10'd339};
ram[30179] = {-9'd59,10'd342};
ram[30180] = {-9'd55,10'd345};
ram[30181] = {-9'd52,10'd348};
ram[30182] = {-9'd49,10'd351};
ram[30183] = {-9'd46,10'd354};
ram[30184] = {-9'd43,10'd358};
ram[30185] = {-9'd40,10'd361};
ram[30186] = {-9'd37,10'd364};
ram[30187] = {-9'd33,10'd367};
ram[30188] = {-9'd30,10'd370};
ram[30189] = {-9'd27,10'd373};
ram[30190] = {-9'd24,10'd376};
ram[30191] = {-9'd21,10'd380};
ram[30192] = {-9'd18,10'd383};
ram[30193] = {-9'd15,10'd386};
ram[30194] = {-9'd11,10'd389};
ram[30195] = {-9'd8,10'd392};
ram[30196] = {-9'd5,10'd395};
ram[30197] = {-9'd2,10'd398};
ram[30198] = {9'd1,-10'd399};
ram[30199] = {9'd4,-10'd396};
ram[30200] = {9'd7,-10'd393};
ram[30201] = {9'd10,-10'd390};
ram[30202] = {9'd14,-10'd387};
ram[30203] = {9'd17,-10'd384};
ram[30204] = {9'd20,-10'd381};
ram[30205] = {9'd23,-10'd377};
ram[30206] = {9'd26,-10'd374};
ram[30207] = {9'd29,-10'd371};
ram[30208] = {9'd29,-10'd371};
ram[30209] = {9'd32,-10'd368};
ram[30210] = {9'd36,-10'd365};
ram[30211] = {9'd39,-10'd362};
ram[30212] = {9'd42,-10'd359};
ram[30213] = {9'd45,-10'd355};
ram[30214] = {9'd48,-10'd352};
ram[30215] = {9'd51,-10'd349};
ram[30216] = {9'd54,-10'd346};
ram[30217] = {9'd58,-10'd343};
ram[30218] = {9'd61,-10'd340};
ram[30219] = {9'd64,-10'd337};
ram[30220] = {9'd67,-10'd334};
ram[30221] = {9'd70,-10'd330};
ram[30222] = {9'd73,-10'd327};
ram[30223] = {9'd76,-10'd324};
ram[30224] = {9'd80,-10'd321};
ram[30225] = {9'd83,-10'd318};
ram[30226] = {9'd86,-10'd315};
ram[30227] = {9'd89,-10'd312};
ram[30228] = {9'd92,-10'd308};
ram[30229] = {9'd95,-10'd305};
ram[30230] = {9'd98,-10'd302};
ram[30231] = {-9'd99,-10'd299};
ram[30232] = {-9'd96,-10'd296};
ram[30233] = {-9'd92,-10'd293};
ram[30234] = {-9'd89,-10'd290};
ram[30235] = {-9'd86,-10'd286};
ram[30236] = {-9'd83,-10'd283};
ram[30237] = {-9'd80,-10'd280};
ram[30238] = {-9'd77,-10'd277};
ram[30239] = {-9'd74,-10'd274};
ram[30240] = {-9'd70,-10'd271};
ram[30241] = {-9'd67,-10'd268};
ram[30242] = {-9'd64,-10'd264};
ram[30243] = {-9'd61,-10'd261};
ram[30244] = {-9'd58,-10'd258};
ram[30245] = {-9'd55,-10'd255};
ram[30246] = {-9'd52,-10'd252};
ram[30247] = {-9'd48,-10'd249};
ram[30248] = {-9'd45,-10'd246};
ram[30249] = {-9'd42,-10'd242};
ram[30250] = {-9'd39,-10'd239};
ram[30251] = {-9'd36,-10'd236};
ram[30252] = {-9'd33,-10'd233};
ram[30253] = {-9'd30,-10'd230};
ram[30254] = {-9'd26,-10'd227};
ram[30255] = {-9'd23,-10'd224};
ram[30256] = {-9'd20,-10'd220};
ram[30257] = {-9'd17,-10'd217};
ram[30258] = {-9'd14,-10'd214};
ram[30259] = {-9'd11,-10'd211};
ram[30260] = {-9'd8,-10'd208};
ram[30261] = {-9'd4,-10'd205};
ram[30262] = {-9'd1,-10'd202};
ram[30263] = {9'd2,-10'd198};
ram[30264] = {9'd5,-10'd195};
ram[30265] = {9'd8,-10'd192};
ram[30266] = {9'd11,-10'd189};
ram[30267] = {9'd14,-10'd186};
ram[30268] = {9'd18,-10'd183};
ram[30269] = {9'd21,-10'd180};
ram[30270] = {9'd24,-10'd176};
ram[30271] = {9'd27,-10'd173};
ram[30272] = {9'd30,-10'd170};
ram[30273] = {9'd33,-10'd167};
ram[30274] = {9'd36,-10'd164};
ram[30275] = {9'd40,-10'd161};
ram[30276] = {9'd43,-10'd158};
ram[30277] = {9'd46,-10'd154};
ram[30278] = {9'd49,-10'd151};
ram[30279] = {9'd52,-10'd148};
ram[30280] = {9'd55,-10'd145};
ram[30281] = {9'd58,-10'd142};
ram[30282] = {9'd62,-10'd139};
ram[30283] = {9'd65,-10'd136};
ram[30284] = {9'd68,-10'd132};
ram[30285] = {9'd71,-10'd129};
ram[30286] = {9'd74,-10'd126};
ram[30287] = {9'd77,-10'd123};
ram[30288] = {9'd80,-10'd120};
ram[30289] = {9'd84,-10'd117};
ram[30290] = {9'd87,-10'd114};
ram[30291] = {9'd90,-10'd110};
ram[30292] = {9'd93,-10'd107};
ram[30293] = {9'd96,-10'd104};
ram[30294] = {9'd99,-10'd101};
ram[30295] = {-9'd98,-10'd98};
ram[30296] = {-9'd95,-10'd95};
ram[30297] = {-9'd92,-10'd92};
ram[30298] = {-9'd88,-10'd88};
ram[30299] = {-9'd85,-10'd85};
ram[30300] = {-9'd82,-10'd82};
ram[30301] = {-9'd79,-10'd79};
ram[30302] = {-9'd76,-10'd76};
ram[30303] = {-9'd73,-10'd73};
ram[30304] = {-9'd70,-10'd70};
ram[30305] = {-9'd66,-10'd66};
ram[30306] = {-9'd63,-10'd63};
ram[30307] = {-9'd60,-10'd60};
ram[30308] = {-9'd57,-10'd57};
ram[30309] = {-9'd54,-10'd54};
ram[30310] = {-9'd51,-10'd51};
ram[30311] = {-9'd48,-10'd48};
ram[30312] = {-9'd44,-10'd44};
ram[30313] = {-9'd41,-10'd41};
ram[30314] = {-9'd38,-10'd38};
ram[30315] = {-9'd35,-10'd35};
ram[30316] = {-9'd32,-10'd32};
ram[30317] = {-9'd29,-10'd29};
ram[30318] = {-9'd26,-10'd26};
ram[30319] = {-9'd22,-10'd22};
ram[30320] = {-9'd19,-10'd19};
ram[30321] = {-9'd16,-10'd16};
ram[30322] = {-9'd13,-10'd13};
ram[30323] = {-9'd10,-10'd10};
ram[30324] = {-9'd7,-10'd7};
ram[30325] = {-9'd4,-10'd4};
ram[30326] = {9'd0,10'd0};
ram[30327] = {9'd3,10'd3};
ram[30328] = {9'd6,10'd6};
ram[30329] = {9'd9,10'd9};
ram[30330] = {9'd12,10'd12};
ram[30331] = {9'd15,10'd15};
ram[30332] = {9'd18,10'd18};
ram[30333] = {9'd21,10'd21};
ram[30334] = {9'd25,10'd25};
ram[30335] = {9'd28,10'd28};
ram[30336] = {9'd28,10'd28};
ram[30337] = {9'd31,10'd31};
ram[30338] = {9'd34,10'd34};
ram[30339] = {9'd37,10'd37};
ram[30340] = {9'd40,10'd40};
ram[30341] = {9'd43,10'd43};
ram[30342] = {9'd47,10'd47};
ram[30343] = {9'd50,10'd50};
ram[30344] = {9'd53,10'd53};
ram[30345] = {9'd56,10'd56};
ram[30346] = {9'd59,10'd59};
ram[30347] = {9'd62,10'd62};
ram[30348] = {9'd65,10'd65};
ram[30349] = {9'd69,10'd69};
ram[30350] = {9'd72,10'd72};
ram[30351] = {9'd75,10'd75};
ram[30352] = {9'd78,10'd78};
ram[30353] = {9'd81,10'd81};
ram[30354] = {9'd84,10'd84};
ram[30355] = {9'd87,10'd87};
ram[30356] = {9'd91,10'd91};
ram[30357] = {9'd94,10'd94};
ram[30358] = {9'd97,10'd97};
ram[30359] = {-9'd100,10'd100};
ram[30360] = {-9'd97,10'd103};
ram[30361] = {-9'd94,10'd106};
ram[30362] = {-9'd91,10'd109};
ram[30363] = {-9'd88,10'd113};
ram[30364] = {-9'd85,10'd116};
ram[30365] = {-9'd81,10'd119};
ram[30366] = {-9'd78,10'd122};
ram[30367] = {-9'd75,10'd125};
ram[30368] = {-9'd72,10'd128};
ram[30369] = {-9'd69,10'd131};
ram[30370] = {-9'd66,10'd135};
ram[30371] = {-9'd63,10'd138};
ram[30372] = {-9'd59,10'd141};
ram[30373] = {-9'd56,10'd144};
ram[30374] = {-9'd53,10'd147};
ram[30375] = {-9'd50,10'd150};
ram[30376] = {-9'd47,10'd153};
ram[30377] = {-9'd44,10'd157};
ram[30378] = {-9'd41,10'd160};
ram[30379] = {-9'd37,10'd163};
ram[30380] = {-9'd34,10'd166};
ram[30381] = {-9'd31,10'd169};
ram[30382] = {-9'd28,10'd172};
ram[30383] = {-9'd25,10'd175};
ram[30384] = {-9'd22,10'd179};
ram[30385] = {-9'd19,10'd182};
ram[30386] = {-9'd15,10'd185};
ram[30387] = {-9'd12,10'd188};
ram[30388] = {-9'd9,10'd191};
ram[30389] = {-9'd6,10'd194};
ram[30390] = {-9'd3,10'd197};
ram[30391] = {9'd0,10'd201};
ram[30392] = {9'd3,10'd204};
ram[30393] = {9'd7,10'd207};
ram[30394] = {9'd10,10'd210};
ram[30395] = {9'd13,10'd213};
ram[30396] = {9'd16,10'd216};
ram[30397] = {9'd19,10'd219};
ram[30398] = {9'd22,10'd223};
ram[30399] = {9'd25,10'd226};
ram[30400] = {9'd29,10'd229};
ram[30401] = {9'd32,10'd232};
ram[30402] = {9'd35,10'd235};
ram[30403] = {9'd38,10'd238};
ram[30404] = {9'd41,10'd241};
ram[30405] = {9'd44,10'd245};
ram[30406] = {9'd47,10'd248};
ram[30407] = {9'd51,10'd251};
ram[30408] = {9'd54,10'd254};
ram[30409] = {9'd57,10'd257};
ram[30410] = {9'd60,10'd260};
ram[30411] = {9'd63,10'd263};
ram[30412] = {9'd66,10'd267};
ram[30413] = {9'd69,10'd270};
ram[30414] = {9'd73,10'd273};
ram[30415] = {9'd76,10'd276};
ram[30416] = {9'd79,10'd279};
ram[30417] = {9'd82,10'd282};
ram[30418] = {9'd85,10'd285};
ram[30419] = {9'd88,10'd289};
ram[30420] = {9'd91,10'd292};
ram[30421] = {9'd95,10'd295};
ram[30422] = {9'd98,10'd298};
ram[30423] = {-9'd99,10'd301};
ram[30424] = {-9'd96,10'd304};
ram[30425] = {-9'd93,10'd307};
ram[30426] = {-9'd90,10'd311};
ram[30427] = {-9'd87,10'd314};
ram[30428] = {-9'd84,10'd317};
ram[30429] = {-9'd81,10'd320};
ram[30430] = {-9'd77,10'd323};
ram[30431] = {-9'd74,10'd326};
ram[30432] = {-9'd71,10'd329};
ram[30433] = {-9'd68,10'd333};
ram[30434] = {-9'd65,10'd336};
ram[30435] = {-9'd62,10'd339};
ram[30436] = {-9'd59,10'd342};
ram[30437] = {-9'd55,10'd345};
ram[30438] = {-9'd52,10'd348};
ram[30439] = {-9'd49,10'd351};
ram[30440] = {-9'd46,10'd354};
ram[30441] = {-9'd43,10'd358};
ram[30442] = {-9'd40,10'd361};
ram[30443] = {-9'd37,10'd364};
ram[30444] = {-9'd33,10'd367};
ram[30445] = {-9'd30,10'd370};
ram[30446] = {-9'd27,10'd373};
ram[30447] = {-9'd24,10'd376};
ram[30448] = {-9'd21,10'd380};
ram[30449] = {-9'd18,10'd383};
ram[30450] = {-9'd15,10'd386};
ram[30451] = {-9'd11,10'd389};
ram[30452] = {-9'd8,10'd392};
ram[30453] = {-9'd5,10'd395};
ram[30454] = {-9'd2,10'd398};
ram[30455] = {9'd1,-10'd399};
ram[30456] = {9'd4,-10'd396};
ram[30457] = {9'd7,-10'd393};
ram[30458] = {9'd10,-10'd390};
ram[30459] = {9'd14,-10'd387};
ram[30460] = {9'd17,-10'd384};
ram[30461] = {9'd20,-10'd381};
ram[30462] = {9'd23,-10'd377};
ram[30463] = {9'd26,-10'd374};
ram[30464] = {9'd26,-10'd374};
ram[30465] = {9'd29,-10'd371};
ram[30466] = {9'd32,-10'd368};
ram[30467] = {9'd36,-10'd365};
ram[30468] = {9'd39,-10'd362};
ram[30469] = {9'd42,-10'd359};
ram[30470] = {9'd45,-10'd355};
ram[30471] = {9'd48,-10'd352};
ram[30472] = {9'd51,-10'd349};
ram[30473] = {9'd54,-10'd346};
ram[30474] = {9'd58,-10'd343};
ram[30475] = {9'd61,-10'd340};
ram[30476] = {9'd64,-10'd337};
ram[30477] = {9'd67,-10'd334};
ram[30478] = {9'd70,-10'd330};
ram[30479] = {9'd73,-10'd327};
ram[30480] = {9'd76,-10'd324};
ram[30481] = {9'd80,-10'd321};
ram[30482] = {9'd83,-10'd318};
ram[30483] = {9'd86,-10'd315};
ram[30484] = {9'd89,-10'd312};
ram[30485] = {9'd92,-10'd308};
ram[30486] = {9'd95,-10'd305};
ram[30487] = {9'd98,-10'd302};
ram[30488] = {-9'd99,-10'd299};
ram[30489] = {-9'd96,-10'd296};
ram[30490] = {-9'd92,-10'd293};
ram[30491] = {-9'd89,-10'd290};
ram[30492] = {-9'd86,-10'd286};
ram[30493] = {-9'd83,-10'd283};
ram[30494] = {-9'd80,-10'd280};
ram[30495] = {-9'd77,-10'd277};
ram[30496] = {-9'd74,-10'd274};
ram[30497] = {-9'd70,-10'd271};
ram[30498] = {-9'd67,-10'd268};
ram[30499] = {-9'd64,-10'd264};
ram[30500] = {-9'd61,-10'd261};
ram[30501] = {-9'd58,-10'd258};
ram[30502] = {-9'd55,-10'd255};
ram[30503] = {-9'd52,-10'd252};
ram[30504] = {-9'd48,-10'd249};
ram[30505] = {-9'd45,-10'd246};
ram[30506] = {-9'd42,-10'd242};
ram[30507] = {-9'd39,-10'd239};
ram[30508] = {-9'd36,-10'd236};
ram[30509] = {-9'd33,-10'd233};
ram[30510] = {-9'd30,-10'd230};
ram[30511] = {-9'd26,-10'd227};
ram[30512] = {-9'd23,-10'd224};
ram[30513] = {-9'd20,-10'd220};
ram[30514] = {-9'd17,-10'd217};
ram[30515] = {-9'd14,-10'd214};
ram[30516] = {-9'd11,-10'd211};
ram[30517] = {-9'd8,-10'd208};
ram[30518] = {-9'd4,-10'd205};
ram[30519] = {-9'd1,-10'd202};
ram[30520] = {9'd2,-10'd198};
ram[30521] = {9'd5,-10'd195};
ram[30522] = {9'd8,-10'd192};
ram[30523] = {9'd11,-10'd189};
ram[30524] = {9'd14,-10'd186};
ram[30525] = {9'd18,-10'd183};
ram[30526] = {9'd21,-10'd180};
ram[30527] = {9'd24,-10'd176};
ram[30528] = {9'd27,-10'd173};
ram[30529] = {9'd30,-10'd170};
ram[30530] = {9'd33,-10'd167};
ram[30531] = {9'd36,-10'd164};
ram[30532] = {9'd40,-10'd161};
ram[30533] = {9'd43,-10'd158};
ram[30534] = {9'd46,-10'd154};
ram[30535] = {9'd49,-10'd151};
ram[30536] = {9'd52,-10'd148};
ram[30537] = {9'd55,-10'd145};
ram[30538] = {9'd58,-10'd142};
ram[30539] = {9'd62,-10'd139};
ram[30540] = {9'd65,-10'd136};
ram[30541] = {9'd68,-10'd132};
ram[30542] = {9'd71,-10'd129};
ram[30543] = {9'd74,-10'd126};
ram[30544] = {9'd77,-10'd123};
ram[30545] = {9'd80,-10'd120};
ram[30546] = {9'd84,-10'd117};
ram[30547] = {9'd87,-10'd114};
ram[30548] = {9'd90,-10'd110};
ram[30549] = {9'd93,-10'd107};
ram[30550] = {9'd96,-10'd104};
ram[30551] = {9'd99,-10'd101};
ram[30552] = {-9'd98,-10'd98};
ram[30553] = {-9'd95,-10'd95};
ram[30554] = {-9'd92,-10'd92};
ram[30555] = {-9'd88,-10'd88};
ram[30556] = {-9'd85,-10'd85};
ram[30557] = {-9'd82,-10'd82};
ram[30558] = {-9'd79,-10'd79};
ram[30559] = {-9'd76,-10'd76};
ram[30560] = {-9'd73,-10'd73};
ram[30561] = {-9'd70,-10'd70};
ram[30562] = {-9'd66,-10'd66};
ram[30563] = {-9'd63,-10'd63};
ram[30564] = {-9'd60,-10'd60};
ram[30565] = {-9'd57,-10'd57};
ram[30566] = {-9'd54,-10'd54};
ram[30567] = {-9'd51,-10'd51};
ram[30568] = {-9'd48,-10'd48};
ram[30569] = {-9'd44,-10'd44};
ram[30570] = {-9'd41,-10'd41};
ram[30571] = {-9'd38,-10'd38};
ram[30572] = {-9'd35,-10'd35};
ram[30573] = {-9'd32,-10'd32};
ram[30574] = {-9'd29,-10'd29};
ram[30575] = {-9'd26,-10'd26};
ram[30576] = {-9'd22,-10'd22};
ram[30577] = {-9'd19,-10'd19};
ram[30578] = {-9'd16,-10'd16};
ram[30579] = {-9'd13,-10'd13};
ram[30580] = {-9'd10,-10'd10};
ram[30581] = {-9'd7,-10'd7};
ram[30582] = {-9'd4,-10'd4};
ram[30583] = {9'd0,10'd0};
ram[30584] = {9'd3,10'd3};
ram[30585] = {9'd6,10'd6};
ram[30586] = {9'd9,10'd9};
ram[30587] = {9'd12,10'd12};
ram[30588] = {9'd15,10'd15};
ram[30589] = {9'd18,10'd18};
ram[30590] = {9'd21,10'd21};
ram[30591] = {9'd25,10'd25};
ram[30592] = {9'd25,10'd25};
ram[30593] = {9'd28,10'd28};
ram[30594] = {9'd31,10'd31};
ram[30595] = {9'd34,10'd34};
ram[30596] = {9'd37,10'd37};
ram[30597] = {9'd40,10'd40};
ram[30598] = {9'd43,10'd43};
ram[30599] = {9'd47,10'd47};
ram[30600] = {9'd50,10'd50};
ram[30601] = {9'd53,10'd53};
ram[30602] = {9'd56,10'd56};
ram[30603] = {9'd59,10'd59};
ram[30604] = {9'd62,10'd62};
ram[30605] = {9'd65,10'd65};
ram[30606] = {9'd69,10'd69};
ram[30607] = {9'd72,10'd72};
ram[30608] = {9'd75,10'd75};
ram[30609] = {9'd78,10'd78};
ram[30610] = {9'd81,10'd81};
ram[30611] = {9'd84,10'd84};
ram[30612] = {9'd87,10'd87};
ram[30613] = {9'd91,10'd91};
ram[30614] = {9'd94,10'd94};
ram[30615] = {9'd97,10'd97};
ram[30616] = {-9'd100,10'd100};
ram[30617] = {-9'd97,10'd103};
ram[30618] = {-9'd94,10'd106};
ram[30619] = {-9'd91,10'd109};
ram[30620] = {-9'd88,10'd113};
ram[30621] = {-9'd85,10'd116};
ram[30622] = {-9'd81,10'd119};
ram[30623] = {-9'd78,10'd122};
ram[30624] = {-9'd75,10'd125};
ram[30625] = {-9'd72,10'd128};
ram[30626] = {-9'd69,10'd131};
ram[30627] = {-9'd66,10'd135};
ram[30628] = {-9'd63,10'd138};
ram[30629] = {-9'd59,10'd141};
ram[30630] = {-9'd56,10'd144};
ram[30631] = {-9'd53,10'd147};
ram[30632] = {-9'd50,10'd150};
ram[30633] = {-9'd47,10'd153};
ram[30634] = {-9'd44,10'd157};
ram[30635] = {-9'd41,10'd160};
ram[30636] = {-9'd37,10'd163};
ram[30637] = {-9'd34,10'd166};
ram[30638] = {-9'd31,10'd169};
ram[30639] = {-9'd28,10'd172};
ram[30640] = {-9'd25,10'd175};
ram[30641] = {-9'd22,10'd179};
ram[30642] = {-9'd19,10'd182};
ram[30643] = {-9'd15,10'd185};
ram[30644] = {-9'd12,10'd188};
ram[30645] = {-9'd9,10'd191};
ram[30646] = {-9'd6,10'd194};
ram[30647] = {-9'd3,10'd197};
ram[30648] = {9'd0,10'd201};
ram[30649] = {9'd3,10'd204};
ram[30650] = {9'd7,10'd207};
ram[30651] = {9'd10,10'd210};
ram[30652] = {9'd13,10'd213};
ram[30653] = {9'd16,10'd216};
ram[30654] = {9'd19,10'd219};
ram[30655] = {9'd22,10'd223};
ram[30656] = {9'd25,10'd226};
ram[30657] = {9'd29,10'd229};
ram[30658] = {9'd32,10'd232};
ram[30659] = {9'd35,10'd235};
ram[30660] = {9'd38,10'd238};
ram[30661] = {9'd41,10'd241};
ram[30662] = {9'd44,10'd245};
ram[30663] = {9'd47,10'd248};
ram[30664] = {9'd51,10'd251};
ram[30665] = {9'd54,10'd254};
ram[30666] = {9'd57,10'd257};
ram[30667] = {9'd60,10'd260};
ram[30668] = {9'd63,10'd263};
ram[30669] = {9'd66,10'd267};
ram[30670] = {9'd69,10'd270};
ram[30671] = {9'd73,10'd273};
ram[30672] = {9'd76,10'd276};
ram[30673] = {9'd79,10'd279};
ram[30674] = {9'd82,10'd282};
ram[30675] = {9'd85,10'd285};
ram[30676] = {9'd88,10'd289};
ram[30677] = {9'd91,10'd292};
ram[30678] = {9'd95,10'd295};
ram[30679] = {9'd98,10'd298};
ram[30680] = {-9'd99,10'd301};
ram[30681] = {-9'd96,10'd304};
ram[30682] = {-9'd93,10'd307};
ram[30683] = {-9'd90,10'd311};
ram[30684] = {-9'd87,10'd314};
ram[30685] = {-9'd84,10'd317};
ram[30686] = {-9'd81,10'd320};
ram[30687] = {-9'd77,10'd323};
ram[30688] = {-9'd74,10'd326};
ram[30689] = {-9'd71,10'd329};
ram[30690] = {-9'd68,10'd333};
ram[30691] = {-9'd65,10'd336};
ram[30692] = {-9'd62,10'd339};
ram[30693] = {-9'd59,10'd342};
ram[30694] = {-9'd55,10'd345};
ram[30695] = {-9'd52,10'd348};
ram[30696] = {-9'd49,10'd351};
ram[30697] = {-9'd46,10'd354};
ram[30698] = {-9'd43,10'd358};
ram[30699] = {-9'd40,10'd361};
ram[30700] = {-9'd37,10'd364};
ram[30701] = {-9'd33,10'd367};
ram[30702] = {-9'd30,10'd370};
ram[30703] = {-9'd27,10'd373};
ram[30704] = {-9'd24,10'd376};
ram[30705] = {-9'd21,10'd380};
ram[30706] = {-9'd18,10'd383};
ram[30707] = {-9'd15,10'd386};
ram[30708] = {-9'd11,10'd389};
ram[30709] = {-9'd8,10'd392};
ram[30710] = {-9'd5,10'd395};
ram[30711] = {-9'd2,10'd398};
ram[30712] = {9'd1,-10'd399};
ram[30713] = {9'd4,-10'd396};
ram[30714] = {9'd7,-10'd393};
ram[30715] = {9'd10,-10'd390};
ram[30716] = {9'd14,-10'd387};
ram[30717] = {9'd17,-10'd384};
ram[30718] = {9'd20,-10'd381};
ram[30719] = {9'd23,-10'd377};
ram[30720] = {9'd23,-10'd377};
ram[30721] = {9'd26,-10'd374};
ram[30722] = {9'd29,-10'd371};
ram[30723] = {9'd32,-10'd368};
ram[30724] = {9'd36,-10'd365};
ram[30725] = {9'd39,-10'd362};
ram[30726] = {9'd42,-10'd359};
ram[30727] = {9'd45,-10'd355};
ram[30728] = {9'd48,-10'd352};
ram[30729] = {9'd51,-10'd349};
ram[30730] = {9'd54,-10'd346};
ram[30731] = {9'd58,-10'd343};
ram[30732] = {9'd61,-10'd340};
ram[30733] = {9'd64,-10'd337};
ram[30734] = {9'd67,-10'd334};
ram[30735] = {9'd70,-10'd330};
ram[30736] = {9'd73,-10'd327};
ram[30737] = {9'd76,-10'd324};
ram[30738] = {9'd80,-10'd321};
ram[30739] = {9'd83,-10'd318};
ram[30740] = {9'd86,-10'd315};
ram[30741] = {9'd89,-10'd312};
ram[30742] = {9'd92,-10'd308};
ram[30743] = {9'd95,-10'd305};
ram[30744] = {9'd98,-10'd302};
ram[30745] = {-9'd99,-10'd299};
ram[30746] = {-9'd96,-10'd296};
ram[30747] = {-9'd92,-10'd293};
ram[30748] = {-9'd89,-10'd290};
ram[30749] = {-9'd86,-10'd286};
ram[30750] = {-9'd83,-10'd283};
ram[30751] = {-9'd80,-10'd280};
ram[30752] = {-9'd77,-10'd277};
ram[30753] = {-9'd74,-10'd274};
ram[30754] = {-9'd70,-10'd271};
ram[30755] = {-9'd67,-10'd268};
ram[30756] = {-9'd64,-10'd264};
ram[30757] = {-9'd61,-10'd261};
ram[30758] = {-9'd58,-10'd258};
ram[30759] = {-9'd55,-10'd255};
ram[30760] = {-9'd52,-10'd252};
ram[30761] = {-9'd48,-10'd249};
ram[30762] = {-9'd45,-10'd246};
ram[30763] = {-9'd42,-10'd242};
ram[30764] = {-9'd39,-10'd239};
ram[30765] = {-9'd36,-10'd236};
ram[30766] = {-9'd33,-10'd233};
ram[30767] = {-9'd30,-10'd230};
ram[30768] = {-9'd26,-10'd227};
ram[30769] = {-9'd23,-10'd224};
ram[30770] = {-9'd20,-10'd220};
ram[30771] = {-9'd17,-10'd217};
ram[30772] = {-9'd14,-10'd214};
ram[30773] = {-9'd11,-10'd211};
ram[30774] = {-9'd8,-10'd208};
ram[30775] = {-9'd4,-10'd205};
ram[30776] = {-9'd1,-10'd202};
ram[30777] = {9'd2,-10'd198};
ram[30778] = {9'd5,-10'd195};
ram[30779] = {9'd8,-10'd192};
ram[30780] = {9'd11,-10'd189};
ram[30781] = {9'd14,-10'd186};
ram[30782] = {9'd18,-10'd183};
ram[30783] = {9'd21,-10'd180};
ram[30784] = {9'd24,-10'd176};
ram[30785] = {9'd27,-10'd173};
ram[30786] = {9'd30,-10'd170};
ram[30787] = {9'd33,-10'd167};
ram[30788] = {9'd36,-10'd164};
ram[30789] = {9'd40,-10'd161};
ram[30790] = {9'd43,-10'd158};
ram[30791] = {9'd46,-10'd154};
ram[30792] = {9'd49,-10'd151};
ram[30793] = {9'd52,-10'd148};
ram[30794] = {9'd55,-10'd145};
ram[30795] = {9'd58,-10'd142};
ram[30796] = {9'd62,-10'd139};
ram[30797] = {9'd65,-10'd136};
ram[30798] = {9'd68,-10'd132};
ram[30799] = {9'd71,-10'd129};
ram[30800] = {9'd74,-10'd126};
ram[30801] = {9'd77,-10'd123};
ram[30802] = {9'd80,-10'd120};
ram[30803] = {9'd84,-10'd117};
ram[30804] = {9'd87,-10'd114};
ram[30805] = {9'd90,-10'd110};
ram[30806] = {9'd93,-10'd107};
ram[30807] = {9'd96,-10'd104};
ram[30808] = {9'd99,-10'd101};
ram[30809] = {-9'd98,-10'd98};
ram[30810] = {-9'd95,-10'd95};
ram[30811] = {-9'd92,-10'd92};
ram[30812] = {-9'd88,-10'd88};
ram[30813] = {-9'd85,-10'd85};
ram[30814] = {-9'd82,-10'd82};
ram[30815] = {-9'd79,-10'd79};
ram[30816] = {-9'd76,-10'd76};
ram[30817] = {-9'd73,-10'd73};
ram[30818] = {-9'd70,-10'd70};
ram[30819] = {-9'd66,-10'd66};
ram[30820] = {-9'd63,-10'd63};
ram[30821] = {-9'd60,-10'd60};
ram[30822] = {-9'd57,-10'd57};
ram[30823] = {-9'd54,-10'd54};
ram[30824] = {-9'd51,-10'd51};
ram[30825] = {-9'd48,-10'd48};
ram[30826] = {-9'd44,-10'd44};
ram[30827] = {-9'd41,-10'd41};
ram[30828] = {-9'd38,-10'd38};
ram[30829] = {-9'd35,-10'd35};
ram[30830] = {-9'd32,-10'd32};
ram[30831] = {-9'd29,-10'd29};
ram[30832] = {-9'd26,-10'd26};
ram[30833] = {-9'd22,-10'd22};
ram[30834] = {-9'd19,-10'd19};
ram[30835] = {-9'd16,-10'd16};
ram[30836] = {-9'd13,-10'd13};
ram[30837] = {-9'd10,-10'd10};
ram[30838] = {-9'd7,-10'd7};
ram[30839] = {-9'd4,-10'd4};
ram[30840] = {9'd0,10'd0};
ram[30841] = {9'd3,10'd3};
ram[30842] = {9'd6,10'd6};
ram[30843] = {9'd9,10'd9};
ram[30844] = {9'd12,10'd12};
ram[30845] = {9'd15,10'd15};
ram[30846] = {9'd18,10'd18};
ram[30847] = {9'd21,10'd21};
ram[30848] = {9'd21,10'd21};
ram[30849] = {9'd25,10'd25};
ram[30850] = {9'd28,10'd28};
ram[30851] = {9'd31,10'd31};
ram[30852] = {9'd34,10'd34};
ram[30853] = {9'd37,10'd37};
ram[30854] = {9'd40,10'd40};
ram[30855] = {9'd43,10'd43};
ram[30856] = {9'd47,10'd47};
ram[30857] = {9'd50,10'd50};
ram[30858] = {9'd53,10'd53};
ram[30859] = {9'd56,10'd56};
ram[30860] = {9'd59,10'd59};
ram[30861] = {9'd62,10'd62};
ram[30862] = {9'd65,10'd65};
ram[30863] = {9'd69,10'd69};
ram[30864] = {9'd72,10'd72};
ram[30865] = {9'd75,10'd75};
ram[30866] = {9'd78,10'd78};
ram[30867] = {9'd81,10'd81};
ram[30868] = {9'd84,10'd84};
ram[30869] = {9'd87,10'd87};
ram[30870] = {9'd91,10'd91};
ram[30871] = {9'd94,10'd94};
ram[30872] = {9'd97,10'd97};
ram[30873] = {-9'd100,10'd100};
ram[30874] = {-9'd97,10'd103};
ram[30875] = {-9'd94,10'd106};
ram[30876] = {-9'd91,10'd109};
ram[30877] = {-9'd88,10'd113};
ram[30878] = {-9'd85,10'd116};
ram[30879] = {-9'd81,10'd119};
ram[30880] = {-9'd78,10'd122};
ram[30881] = {-9'd75,10'd125};
ram[30882] = {-9'd72,10'd128};
ram[30883] = {-9'd69,10'd131};
ram[30884] = {-9'd66,10'd135};
ram[30885] = {-9'd63,10'd138};
ram[30886] = {-9'd59,10'd141};
ram[30887] = {-9'd56,10'd144};
ram[30888] = {-9'd53,10'd147};
ram[30889] = {-9'd50,10'd150};
ram[30890] = {-9'd47,10'd153};
ram[30891] = {-9'd44,10'd157};
ram[30892] = {-9'd41,10'd160};
ram[30893] = {-9'd37,10'd163};
ram[30894] = {-9'd34,10'd166};
ram[30895] = {-9'd31,10'd169};
ram[30896] = {-9'd28,10'd172};
ram[30897] = {-9'd25,10'd175};
ram[30898] = {-9'd22,10'd179};
ram[30899] = {-9'd19,10'd182};
ram[30900] = {-9'd15,10'd185};
ram[30901] = {-9'd12,10'd188};
ram[30902] = {-9'd9,10'd191};
ram[30903] = {-9'd6,10'd194};
ram[30904] = {-9'd3,10'd197};
ram[30905] = {9'd0,10'd201};
ram[30906] = {9'd3,10'd204};
ram[30907] = {9'd7,10'd207};
ram[30908] = {9'd10,10'd210};
ram[30909] = {9'd13,10'd213};
ram[30910] = {9'd16,10'd216};
ram[30911] = {9'd19,10'd219};
ram[30912] = {9'd22,10'd223};
ram[30913] = {9'd25,10'd226};
ram[30914] = {9'd29,10'd229};
ram[30915] = {9'd32,10'd232};
ram[30916] = {9'd35,10'd235};
ram[30917] = {9'd38,10'd238};
ram[30918] = {9'd41,10'd241};
ram[30919] = {9'd44,10'd245};
ram[30920] = {9'd47,10'd248};
ram[30921] = {9'd51,10'd251};
ram[30922] = {9'd54,10'd254};
ram[30923] = {9'd57,10'd257};
ram[30924] = {9'd60,10'd260};
ram[30925] = {9'd63,10'd263};
ram[30926] = {9'd66,10'd267};
ram[30927] = {9'd69,10'd270};
ram[30928] = {9'd73,10'd273};
ram[30929] = {9'd76,10'd276};
ram[30930] = {9'd79,10'd279};
ram[30931] = {9'd82,10'd282};
ram[30932] = {9'd85,10'd285};
ram[30933] = {9'd88,10'd289};
ram[30934] = {9'd91,10'd292};
ram[30935] = {9'd95,10'd295};
ram[30936] = {9'd98,10'd298};
ram[30937] = {-9'd99,10'd301};
ram[30938] = {-9'd96,10'd304};
ram[30939] = {-9'd93,10'd307};
ram[30940] = {-9'd90,10'd311};
ram[30941] = {-9'd87,10'd314};
ram[30942] = {-9'd84,10'd317};
ram[30943] = {-9'd81,10'd320};
ram[30944] = {-9'd77,10'd323};
ram[30945] = {-9'd74,10'd326};
ram[30946] = {-9'd71,10'd329};
ram[30947] = {-9'd68,10'd333};
ram[30948] = {-9'd65,10'd336};
ram[30949] = {-9'd62,10'd339};
ram[30950] = {-9'd59,10'd342};
ram[30951] = {-9'd55,10'd345};
ram[30952] = {-9'd52,10'd348};
ram[30953] = {-9'd49,10'd351};
ram[30954] = {-9'd46,10'd354};
ram[30955] = {-9'd43,10'd358};
ram[30956] = {-9'd40,10'd361};
ram[30957] = {-9'd37,10'd364};
ram[30958] = {-9'd33,10'd367};
ram[30959] = {-9'd30,10'd370};
ram[30960] = {-9'd27,10'd373};
ram[30961] = {-9'd24,10'd376};
ram[30962] = {-9'd21,10'd380};
ram[30963] = {-9'd18,10'd383};
ram[30964] = {-9'd15,10'd386};
ram[30965] = {-9'd11,10'd389};
ram[30966] = {-9'd8,10'd392};
ram[30967] = {-9'd5,10'd395};
ram[30968] = {-9'd2,10'd398};
ram[30969] = {9'd1,-10'd399};
ram[30970] = {9'd4,-10'd396};
ram[30971] = {9'd7,-10'd393};
ram[30972] = {9'd10,-10'd390};
ram[30973] = {9'd14,-10'd387};
ram[30974] = {9'd17,-10'd384};
ram[30975] = {9'd20,-10'd381};
ram[30976] = {9'd20,-10'd381};
ram[30977] = {9'd23,-10'd377};
ram[30978] = {9'd26,-10'd374};
ram[30979] = {9'd29,-10'd371};
ram[30980] = {9'd32,-10'd368};
ram[30981] = {9'd36,-10'd365};
ram[30982] = {9'd39,-10'd362};
ram[30983] = {9'd42,-10'd359};
ram[30984] = {9'd45,-10'd355};
ram[30985] = {9'd48,-10'd352};
ram[30986] = {9'd51,-10'd349};
ram[30987] = {9'd54,-10'd346};
ram[30988] = {9'd58,-10'd343};
ram[30989] = {9'd61,-10'd340};
ram[30990] = {9'd64,-10'd337};
ram[30991] = {9'd67,-10'd334};
ram[30992] = {9'd70,-10'd330};
ram[30993] = {9'd73,-10'd327};
ram[30994] = {9'd76,-10'd324};
ram[30995] = {9'd80,-10'd321};
ram[30996] = {9'd83,-10'd318};
ram[30997] = {9'd86,-10'd315};
ram[30998] = {9'd89,-10'd312};
ram[30999] = {9'd92,-10'd308};
ram[31000] = {9'd95,-10'd305};
ram[31001] = {9'd98,-10'd302};
ram[31002] = {-9'd99,-10'd299};
ram[31003] = {-9'd96,-10'd296};
ram[31004] = {-9'd92,-10'd293};
ram[31005] = {-9'd89,-10'd290};
ram[31006] = {-9'd86,-10'd286};
ram[31007] = {-9'd83,-10'd283};
ram[31008] = {-9'd80,-10'd280};
ram[31009] = {-9'd77,-10'd277};
ram[31010] = {-9'd74,-10'd274};
ram[31011] = {-9'd70,-10'd271};
ram[31012] = {-9'd67,-10'd268};
ram[31013] = {-9'd64,-10'd264};
ram[31014] = {-9'd61,-10'd261};
ram[31015] = {-9'd58,-10'd258};
ram[31016] = {-9'd55,-10'd255};
ram[31017] = {-9'd52,-10'd252};
ram[31018] = {-9'd48,-10'd249};
ram[31019] = {-9'd45,-10'd246};
ram[31020] = {-9'd42,-10'd242};
ram[31021] = {-9'd39,-10'd239};
ram[31022] = {-9'd36,-10'd236};
ram[31023] = {-9'd33,-10'd233};
ram[31024] = {-9'd30,-10'd230};
ram[31025] = {-9'd26,-10'd227};
ram[31026] = {-9'd23,-10'd224};
ram[31027] = {-9'd20,-10'd220};
ram[31028] = {-9'd17,-10'd217};
ram[31029] = {-9'd14,-10'd214};
ram[31030] = {-9'd11,-10'd211};
ram[31031] = {-9'd8,-10'd208};
ram[31032] = {-9'd4,-10'd205};
ram[31033] = {-9'd1,-10'd202};
ram[31034] = {9'd2,-10'd198};
ram[31035] = {9'd5,-10'd195};
ram[31036] = {9'd8,-10'd192};
ram[31037] = {9'd11,-10'd189};
ram[31038] = {9'd14,-10'd186};
ram[31039] = {9'd18,-10'd183};
ram[31040] = {9'd21,-10'd180};
ram[31041] = {9'd24,-10'd176};
ram[31042] = {9'd27,-10'd173};
ram[31043] = {9'd30,-10'd170};
ram[31044] = {9'd33,-10'd167};
ram[31045] = {9'd36,-10'd164};
ram[31046] = {9'd40,-10'd161};
ram[31047] = {9'd43,-10'd158};
ram[31048] = {9'd46,-10'd154};
ram[31049] = {9'd49,-10'd151};
ram[31050] = {9'd52,-10'd148};
ram[31051] = {9'd55,-10'd145};
ram[31052] = {9'd58,-10'd142};
ram[31053] = {9'd62,-10'd139};
ram[31054] = {9'd65,-10'd136};
ram[31055] = {9'd68,-10'd132};
ram[31056] = {9'd71,-10'd129};
ram[31057] = {9'd74,-10'd126};
ram[31058] = {9'd77,-10'd123};
ram[31059] = {9'd80,-10'd120};
ram[31060] = {9'd84,-10'd117};
ram[31061] = {9'd87,-10'd114};
ram[31062] = {9'd90,-10'd110};
ram[31063] = {9'd93,-10'd107};
ram[31064] = {9'd96,-10'd104};
ram[31065] = {9'd99,-10'd101};
ram[31066] = {-9'd98,-10'd98};
ram[31067] = {-9'd95,-10'd95};
ram[31068] = {-9'd92,-10'd92};
ram[31069] = {-9'd88,-10'd88};
ram[31070] = {-9'd85,-10'd85};
ram[31071] = {-9'd82,-10'd82};
ram[31072] = {-9'd79,-10'd79};
ram[31073] = {-9'd76,-10'd76};
ram[31074] = {-9'd73,-10'd73};
ram[31075] = {-9'd70,-10'd70};
ram[31076] = {-9'd66,-10'd66};
ram[31077] = {-9'd63,-10'd63};
ram[31078] = {-9'd60,-10'd60};
ram[31079] = {-9'd57,-10'd57};
ram[31080] = {-9'd54,-10'd54};
ram[31081] = {-9'd51,-10'd51};
ram[31082] = {-9'd48,-10'd48};
ram[31083] = {-9'd44,-10'd44};
ram[31084] = {-9'd41,-10'd41};
ram[31085] = {-9'd38,-10'd38};
ram[31086] = {-9'd35,-10'd35};
ram[31087] = {-9'd32,-10'd32};
ram[31088] = {-9'd29,-10'd29};
ram[31089] = {-9'd26,-10'd26};
ram[31090] = {-9'd22,-10'd22};
ram[31091] = {-9'd19,-10'd19};
ram[31092] = {-9'd16,-10'd16};
ram[31093] = {-9'd13,-10'd13};
ram[31094] = {-9'd10,-10'd10};
ram[31095] = {-9'd7,-10'd7};
ram[31096] = {-9'd4,-10'd4};
ram[31097] = {9'd0,10'd0};
ram[31098] = {9'd3,10'd3};
ram[31099] = {9'd6,10'd6};
ram[31100] = {9'd9,10'd9};
ram[31101] = {9'd12,10'd12};
ram[31102] = {9'd15,10'd15};
ram[31103] = {9'd18,10'd18};
ram[31104] = {9'd18,10'd18};
ram[31105] = {9'd21,10'd21};
ram[31106] = {9'd25,10'd25};
ram[31107] = {9'd28,10'd28};
ram[31108] = {9'd31,10'd31};
ram[31109] = {9'd34,10'd34};
ram[31110] = {9'd37,10'd37};
ram[31111] = {9'd40,10'd40};
ram[31112] = {9'd43,10'd43};
ram[31113] = {9'd47,10'd47};
ram[31114] = {9'd50,10'd50};
ram[31115] = {9'd53,10'd53};
ram[31116] = {9'd56,10'd56};
ram[31117] = {9'd59,10'd59};
ram[31118] = {9'd62,10'd62};
ram[31119] = {9'd65,10'd65};
ram[31120] = {9'd69,10'd69};
ram[31121] = {9'd72,10'd72};
ram[31122] = {9'd75,10'd75};
ram[31123] = {9'd78,10'd78};
ram[31124] = {9'd81,10'd81};
ram[31125] = {9'd84,10'd84};
ram[31126] = {9'd87,10'd87};
ram[31127] = {9'd91,10'd91};
ram[31128] = {9'd94,10'd94};
ram[31129] = {9'd97,10'd97};
ram[31130] = {-9'd100,10'd100};
ram[31131] = {-9'd97,10'd103};
ram[31132] = {-9'd94,10'd106};
ram[31133] = {-9'd91,10'd109};
ram[31134] = {-9'd88,10'd113};
ram[31135] = {-9'd85,10'd116};
ram[31136] = {-9'd81,10'd119};
ram[31137] = {-9'd78,10'd122};
ram[31138] = {-9'd75,10'd125};
ram[31139] = {-9'd72,10'd128};
ram[31140] = {-9'd69,10'd131};
ram[31141] = {-9'd66,10'd135};
ram[31142] = {-9'd63,10'd138};
ram[31143] = {-9'd59,10'd141};
ram[31144] = {-9'd56,10'd144};
ram[31145] = {-9'd53,10'd147};
ram[31146] = {-9'd50,10'd150};
ram[31147] = {-9'd47,10'd153};
ram[31148] = {-9'd44,10'd157};
ram[31149] = {-9'd41,10'd160};
ram[31150] = {-9'd37,10'd163};
ram[31151] = {-9'd34,10'd166};
ram[31152] = {-9'd31,10'd169};
ram[31153] = {-9'd28,10'd172};
ram[31154] = {-9'd25,10'd175};
ram[31155] = {-9'd22,10'd179};
ram[31156] = {-9'd19,10'd182};
ram[31157] = {-9'd15,10'd185};
ram[31158] = {-9'd12,10'd188};
ram[31159] = {-9'd9,10'd191};
ram[31160] = {-9'd6,10'd194};
ram[31161] = {-9'd3,10'd197};
ram[31162] = {9'd0,10'd201};
ram[31163] = {9'd3,10'd204};
ram[31164] = {9'd7,10'd207};
ram[31165] = {9'd10,10'd210};
ram[31166] = {9'd13,10'd213};
ram[31167] = {9'd16,10'd216};
ram[31168] = {9'd19,10'd219};
ram[31169] = {9'd22,10'd223};
ram[31170] = {9'd25,10'd226};
ram[31171] = {9'd29,10'd229};
ram[31172] = {9'd32,10'd232};
ram[31173] = {9'd35,10'd235};
ram[31174] = {9'd38,10'd238};
ram[31175] = {9'd41,10'd241};
ram[31176] = {9'd44,10'd245};
ram[31177] = {9'd47,10'd248};
ram[31178] = {9'd51,10'd251};
ram[31179] = {9'd54,10'd254};
ram[31180] = {9'd57,10'd257};
ram[31181] = {9'd60,10'd260};
ram[31182] = {9'd63,10'd263};
ram[31183] = {9'd66,10'd267};
ram[31184] = {9'd69,10'd270};
ram[31185] = {9'd73,10'd273};
ram[31186] = {9'd76,10'd276};
ram[31187] = {9'd79,10'd279};
ram[31188] = {9'd82,10'd282};
ram[31189] = {9'd85,10'd285};
ram[31190] = {9'd88,10'd289};
ram[31191] = {9'd91,10'd292};
ram[31192] = {9'd95,10'd295};
ram[31193] = {9'd98,10'd298};
ram[31194] = {-9'd99,10'd301};
ram[31195] = {-9'd96,10'd304};
ram[31196] = {-9'd93,10'd307};
ram[31197] = {-9'd90,10'd311};
ram[31198] = {-9'd87,10'd314};
ram[31199] = {-9'd84,10'd317};
ram[31200] = {-9'd81,10'd320};
ram[31201] = {-9'd77,10'd323};
ram[31202] = {-9'd74,10'd326};
ram[31203] = {-9'd71,10'd329};
ram[31204] = {-9'd68,10'd333};
ram[31205] = {-9'd65,10'd336};
ram[31206] = {-9'd62,10'd339};
ram[31207] = {-9'd59,10'd342};
ram[31208] = {-9'd55,10'd345};
ram[31209] = {-9'd52,10'd348};
ram[31210] = {-9'd49,10'd351};
ram[31211] = {-9'd46,10'd354};
ram[31212] = {-9'd43,10'd358};
ram[31213] = {-9'd40,10'd361};
ram[31214] = {-9'd37,10'd364};
ram[31215] = {-9'd33,10'd367};
ram[31216] = {-9'd30,10'd370};
ram[31217] = {-9'd27,10'd373};
ram[31218] = {-9'd24,10'd376};
ram[31219] = {-9'd21,10'd380};
ram[31220] = {-9'd18,10'd383};
ram[31221] = {-9'd15,10'd386};
ram[31222] = {-9'd11,10'd389};
ram[31223] = {-9'd8,10'd392};
ram[31224] = {-9'd5,10'd395};
ram[31225] = {-9'd2,10'd398};
ram[31226] = {9'd1,-10'd399};
ram[31227] = {9'd4,-10'd396};
ram[31228] = {9'd7,-10'd393};
ram[31229] = {9'd10,-10'd390};
ram[31230] = {9'd14,-10'd387};
ram[31231] = {9'd17,-10'd384};
ram[31232] = {9'd17,-10'd384};
ram[31233] = {9'd20,-10'd381};
ram[31234] = {9'd23,-10'd377};
ram[31235] = {9'd26,-10'd374};
ram[31236] = {9'd29,-10'd371};
ram[31237] = {9'd32,-10'd368};
ram[31238] = {9'd36,-10'd365};
ram[31239] = {9'd39,-10'd362};
ram[31240] = {9'd42,-10'd359};
ram[31241] = {9'd45,-10'd355};
ram[31242] = {9'd48,-10'd352};
ram[31243] = {9'd51,-10'd349};
ram[31244] = {9'd54,-10'd346};
ram[31245] = {9'd58,-10'd343};
ram[31246] = {9'd61,-10'd340};
ram[31247] = {9'd64,-10'd337};
ram[31248] = {9'd67,-10'd334};
ram[31249] = {9'd70,-10'd330};
ram[31250] = {9'd73,-10'd327};
ram[31251] = {9'd76,-10'd324};
ram[31252] = {9'd80,-10'd321};
ram[31253] = {9'd83,-10'd318};
ram[31254] = {9'd86,-10'd315};
ram[31255] = {9'd89,-10'd312};
ram[31256] = {9'd92,-10'd308};
ram[31257] = {9'd95,-10'd305};
ram[31258] = {9'd98,-10'd302};
ram[31259] = {-9'd99,-10'd299};
ram[31260] = {-9'd96,-10'd296};
ram[31261] = {-9'd92,-10'd293};
ram[31262] = {-9'd89,-10'd290};
ram[31263] = {-9'd86,-10'd286};
ram[31264] = {-9'd83,-10'd283};
ram[31265] = {-9'd80,-10'd280};
ram[31266] = {-9'd77,-10'd277};
ram[31267] = {-9'd74,-10'd274};
ram[31268] = {-9'd70,-10'd271};
ram[31269] = {-9'd67,-10'd268};
ram[31270] = {-9'd64,-10'd264};
ram[31271] = {-9'd61,-10'd261};
ram[31272] = {-9'd58,-10'd258};
ram[31273] = {-9'd55,-10'd255};
ram[31274] = {-9'd52,-10'd252};
ram[31275] = {-9'd48,-10'd249};
ram[31276] = {-9'd45,-10'd246};
ram[31277] = {-9'd42,-10'd242};
ram[31278] = {-9'd39,-10'd239};
ram[31279] = {-9'd36,-10'd236};
ram[31280] = {-9'd33,-10'd233};
ram[31281] = {-9'd30,-10'd230};
ram[31282] = {-9'd26,-10'd227};
ram[31283] = {-9'd23,-10'd224};
ram[31284] = {-9'd20,-10'd220};
ram[31285] = {-9'd17,-10'd217};
ram[31286] = {-9'd14,-10'd214};
ram[31287] = {-9'd11,-10'd211};
ram[31288] = {-9'd8,-10'd208};
ram[31289] = {-9'd4,-10'd205};
ram[31290] = {-9'd1,-10'd202};
ram[31291] = {9'd2,-10'd198};
ram[31292] = {9'd5,-10'd195};
ram[31293] = {9'd8,-10'd192};
ram[31294] = {9'd11,-10'd189};
ram[31295] = {9'd14,-10'd186};
ram[31296] = {9'd18,-10'd183};
ram[31297] = {9'd21,-10'd180};
ram[31298] = {9'd24,-10'd176};
ram[31299] = {9'd27,-10'd173};
ram[31300] = {9'd30,-10'd170};
ram[31301] = {9'd33,-10'd167};
ram[31302] = {9'd36,-10'd164};
ram[31303] = {9'd40,-10'd161};
ram[31304] = {9'd43,-10'd158};
ram[31305] = {9'd46,-10'd154};
ram[31306] = {9'd49,-10'd151};
ram[31307] = {9'd52,-10'd148};
ram[31308] = {9'd55,-10'd145};
ram[31309] = {9'd58,-10'd142};
ram[31310] = {9'd62,-10'd139};
ram[31311] = {9'd65,-10'd136};
ram[31312] = {9'd68,-10'd132};
ram[31313] = {9'd71,-10'd129};
ram[31314] = {9'd74,-10'd126};
ram[31315] = {9'd77,-10'd123};
ram[31316] = {9'd80,-10'd120};
ram[31317] = {9'd84,-10'd117};
ram[31318] = {9'd87,-10'd114};
ram[31319] = {9'd90,-10'd110};
ram[31320] = {9'd93,-10'd107};
ram[31321] = {9'd96,-10'd104};
ram[31322] = {9'd99,-10'd101};
ram[31323] = {-9'd98,-10'd98};
ram[31324] = {-9'd95,-10'd95};
ram[31325] = {-9'd92,-10'd92};
ram[31326] = {-9'd88,-10'd88};
ram[31327] = {-9'd85,-10'd85};
ram[31328] = {-9'd82,-10'd82};
ram[31329] = {-9'd79,-10'd79};
ram[31330] = {-9'd76,-10'd76};
ram[31331] = {-9'd73,-10'd73};
ram[31332] = {-9'd70,-10'd70};
ram[31333] = {-9'd66,-10'd66};
ram[31334] = {-9'd63,-10'd63};
ram[31335] = {-9'd60,-10'd60};
ram[31336] = {-9'd57,-10'd57};
ram[31337] = {-9'd54,-10'd54};
ram[31338] = {-9'd51,-10'd51};
ram[31339] = {-9'd48,-10'd48};
ram[31340] = {-9'd44,-10'd44};
ram[31341] = {-9'd41,-10'd41};
ram[31342] = {-9'd38,-10'd38};
ram[31343] = {-9'd35,-10'd35};
ram[31344] = {-9'd32,-10'd32};
ram[31345] = {-9'd29,-10'd29};
ram[31346] = {-9'd26,-10'd26};
ram[31347] = {-9'd22,-10'd22};
ram[31348] = {-9'd19,-10'd19};
ram[31349] = {-9'd16,-10'd16};
ram[31350] = {-9'd13,-10'd13};
ram[31351] = {-9'd10,-10'd10};
ram[31352] = {-9'd7,-10'd7};
ram[31353] = {-9'd4,-10'd4};
ram[31354] = {9'd0,10'd0};
ram[31355] = {9'd3,10'd3};
ram[31356] = {9'd6,10'd6};
ram[31357] = {9'd9,10'd9};
ram[31358] = {9'd12,10'd12};
ram[31359] = {9'd15,10'd15};
ram[31360] = {9'd15,10'd15};
ram[31361] = {9'd18,10'd18};
ram[31362] = {9'd21,10'd21};
ram[31363] = {9'd25,10'd25};
ram[31364] = {9'd28,10'd28};
ram[31365] = {9'd31,10'd31};
ram[31366] = {9'd34,10'd34};
ram[31367] = {9'd37,10'd37};
ram[31368] = {9'd40,10'd40};
ram[31369] = {9'd43,10'd43};
ram[31370] = {9'd47,10'd47};
ram[31371] = {9'd50,10'd50};
ram[31372] = {9'd53,10'd53};
ram[31373] = {9'd56,10'd56};
ram[31374] = {9'd59,10'd59};
ram[31375] = {9'd62,10'd62};
ram[31376] = {9'd65,10'd65};
ram[31377] = {9'd69,10'd69};
ram[31378] = {9'd72,10'd72};
ram[31379] = {9'd75,10'd75};
ram[31380] = {9'd78,10'd78};
ram[31381] = {9'd81,10'd81};
ram[31382] = {9'd84,10'd84};
ram[31383] = {9'd87,10'd87};
ram[31384] = {9'd91,10'd91};
ram[31385] = {9'd94,10'd94};
ram[31386] = {9'd97,10'd97};
ram[31387] = {-9'd100,10'd100};
ram[31388] = {-9'd97,10'd103};
ram[31389] = {-9'd94,10'd106};
ram[31390] = {-9'd91,10'd109};
ram[31391] = {-9'd88,10'd113};
ram[31392] = {-9'd85,10'd116};
ram[31393] = {-9'd81,10'd119};
ram[31394] = {-9'd78,10'd122};
ram[31395] = {-9'd75,10'd125};
ram[31396] = {-9'd72,10'd128};
ram[31397] = {-9'd69,10'd131};
ram[31398] = {-9'd66,10'd135};
ram[31399] = {-9'd63,10'd138};
ram[31400] = {-9'd59,10'd141};
ram[31401] = {-9'd56,10'd144};
ram[31402] = {-9'd53,10'd147};
ram[31403] = {-9'd50,10'd150};
ram[31404] = {-9'd47,10'd153};
ram[31405] = {-9'd44,10'd157};
ram[31406] = {-9'd41,10'd160};
ram[31407] = {-9'd37,10'd163};
ram[31408] = {-9'd34,10'd166};
ram[31409] = {-9'd31,10'd169};
ram[31410] = {-9'd28,10'd172};
ram[31411] = {-9'd25,10'd175};
ram[31412] = {-9'd22,10'd179};
ram[31413] = {-9'd19,10'd182};
ram[31414] = {-9'd15,10'd185};
ram[31415] = {-9'd12,10'd188};
ram[31416] = {-9'd9,10'd191};
ram[31417] = {-9'd6,10'd194};
ram[31418] = {-9'd3,10'd197};
ram[31419] = {9'd0,10'd201};
ram[31420] = {9'd3,10'd204};
ram[31421] = {9'd7,10'd207};
ram[31422] = {9'd10,10'd210};
ram[31423] = {9'd13,10'd213};
ram[31424] = {9'd16,10'd216};
ram[31425] = {9'd19,10'd219};
ram[31426] = {9'd22,10'd223};
ram[31427] = {9'd25,10'd226};
ram[31428] = {9'd29,10'd229};
ram[31429] = {9'd32,10'd232};
ram[31430] = {9'd35,10'd235};
ram[31431] = {9'd38,10'd238};
ram[31432] = {9'd41,10'd241};
ram[31433] = {9'd44,10'd245};
ram[31434] = {9'd47,10'd248};
ram[31435] = {9'd51,10'd251};
ram[31436] = {9'd54,10'd254};
ram[31437] = {9'd57,10'd257};
ram[31438] = {9'd60,10'd260};
ram[31439] = {9'd63,10'd263};
ram[31440] = {9'd66,10'd267};
ram[31441] = {9'd69,10'd270};
ram[31442] = {9'd73,10'd273};
ram[31443] = {9'd76,10'd276};
ram[31444] = {9'd79,10'd279};
ram[31445] = {9'd82,10'd282};
ram[31446] = {9'd85,10'd285};
ram[31447] = {9'd88,10'd289};
ram[31448] = {9'd91,10'd292};
ram[31449] = {9'd95,10'd295};
ram[31450] = {9'd98,10'd298};
ram[31451] = {-9'd99,10'd301};
ram[31452] = {-9'd96,10'd304};
ram[31453] = {-9'd93,10'd307};
ram[31454] = {-9'd90,10'd311};
ram[31455] = {-9'd87,10'd314};
ram[31456] = {-9'd84,10'd317};
ram[31457] = {-9'd81,10'd320};
ram[31458] = {-9'd77,10'd323};
ram[31459] = {-9'd74,10'd326};
ram[31460] = {-9'd71,10'd329};
ram[31461] = {-9'd68,10'd333};
ram[31462] = {-9'd65,10'd336};
ram[31463] = {-9'd62,10'd339};
ram[31464] = {-9'd59,10'd342};
ram[31465] = {-9'd55,10'd345};
ram[31466] = {-9'd52,10'd348};
ram[31467] = {-9'd49,10'd351};
ram[31468] = {-9'd46,10'd354};
ram[31469] = {-9'd43,10'd358};
ram[31470] = {-9'd40,10'd361};
ram[31471] = {-9'd37,10'd364};
ram[31472] = {-9'd33,10'd367};
ram[31473] = {-9'd30,10'd370};
ram[31474] = {-9'd27,10'd373};
ram[31475] = {-9'd24,10'd376};
ram[31476] = {-9'd21,10'd380};
ram[31477] = {-9'd18,10'd383};
ram[31478] = {-9'd15,10'd386};
ram[31479] = {-9'd11,10'd389};
ram[31480] = {-9'd8,10'd392};
ram[31481] = {-9'd5,10'd395};
ram[31482] = {-9'd2,10'd398};
ram[31483] = {9'd1,-10'd399};
ram[31484] = {9'd4,-10'd396};
ram[31485] = {9'd7,-10'd393};
ram[31486] = {9'd10,-10'd390};
ram[31487] = {9'd14,-10'd387};
ram[31488] = {9'd14,-10'd387};
ram[31489] = {9'd17,-10'd384};
ram[31490] = {9'd20,-10'd381};
ram[31491] = {9'd23,-10'd377};
ram[31492] = {9'd26,-10'd374};
ram[31493] = {9'd29,-10'd371};
ram[31494] = {9'd32,-10'd368};
ram[31495] = {9'd36,-10'd365};
ram[31496] = {9'd39,-10'd362};
ram[31497] = {9'd42,-10'd359};
ram[31498] = {9'd45,-10'd355};
ram[31499] = {9'd48,-10'd352};
ram[31500] = {9'd51,-10'd349};
ram[31501] = {9'd54,-10'd346};
ram[31502] = {9'd58,-10'd343};
ram[31503] = {9'd61,-10'd340};
ram[31504] = {9'd64,-10'd337};
ram[31505] = {9'd67,-10'd334};
ram[31506] = {9'd70,-10'd330};
ram[31507] = {9'd73,-10'd327};
ram[31508] = {9'd76,-10'd324};
ram[31509] = {9'd80,-10'd321};
ram[31510] = {9'd83,-10'd318};
ram[31511] = {9'd86,-10'd315};
ram[31512] = {9'd89,-10'd312};
ram[31513] = {9'd92,-10'd308};
ram[31514] = {9'd95,-10'd305};
ram[31515] = {9'd98,-10'd302};
ram[31516] = {-9'd99,-10'd299};
ram[31517] = {-9'd96,-10'd296};
ram[31518] = {-9'd92,-10'd293};
ram[31519] = {-9'd89,-10'd290};
ram[31520] = {-9'd86,-10'd286};
ram[31521] = {-9'd83,-10'd283};
ram[31522] = {-9'd80,-10'd280};
ram[31523] = {-9'd77,-10'd277};
ram[31524] = {-9'd74,-10'd274};
ram[31525] = {-9'd70,-10'd271};
ram[31526] = {-9'd67,-10'd268};
ram[31527] = {-9'd64,-10'd264};
ram[31528] = {-9'd61,-10'd261};
ram[31529] = {-9'd58,-10'd258};
ram[31530] = {-9'd55,-10'd255};
ram[31531] = {-9'd52,-10'd252};
ram[31532] = {-9'd48,-10'd249};
ram[31533] = {-9'd45,-10'd246};
ram[31534] = {-9'd42,-10'd242};
ram[31535] = {-9'd39,-10'd239};
ram[31536] = {-9'd36,-10'd236};
ram[31537] = {-9'd33,-10'd233};
ram[31538] = {-9'd30,-10'd230};
ram[31539] = {-9'd26,-10'd227};
ram[31540] = {-9'd23,-10'd224};
ram[31541] = {-9'd20,-10'd220};
ram[31542] = {-9'd17,-10'd217};
ram[31543] = {-9'd14,-10'd214};
ram[31544] = {-9'd11,-10'd211};
ram[31545] = {-9'd8,-10'd208};
ram[31546] = {-9'd4,-10'd205};
ram[31547] = {-9'd1,-10'd202};
ram[31548] = {9'd2,-10'd198};
ram[31549] = {9'd5,-10'd195};
ram[31550] = {9'd8,-10'd192};
ram[31551] = {9'd11,-10'd189};
ram[31552] = {9'd14,-10'd186};
ram[31553] = {9'd18,-10'd183};
ram[31554] = {9'd21,-10'd180};
ram[31555] = {9'd24,-10'd176};
ram[31556] = {9'd27,-10'd173};
ram[31557] = {9'd30,-10'd170};
ram[31558] = {9'd33,-10'd167};
ram[31559] = {9'd36,-10'd164};
ram[31560] = {9'd40,-10'd161};
ram[31561] = {9'd43,-10'd158};
ram[31562] = {9'd46,-10'd154};
ram[31563] = {9'd49,-10'd151};
ram[31564] = {9'd52,-10'd148};
ram[31565] = {9'd55,-10'd145};
ram[31566] = {9'd58,-10'd142};
ram[31567] = {9'd62,-10'd139};
ram[31568] = {9'd65,-10'd136};
ram[31569] = {9'd68,-10'd132};
ram[31570] = {9'd71,-10'd129};
ram[31571] = {9'd74,-10'd126};
ram[31572] = {9'd77,-10'd123};
ram[31573] = {9'd80,-10'd120};
ram[31574] = {9'd84,-10'd117};
ram[31575] = {9'd87,-10'd114};
ram[31576] = {9'd90,-10'd110};
ram[31577] = {9'd93,-10'd107};
ram[31578] = {9'd96,-10'd104};
ram[31579] = {9'd99,-10'd101};
ram[31580] = {-9'd98,-10'd98};
ram[31581] = {-9'd95,-10'd95};
ram[31582] = {-9'd92,-10'd92};
ram[31583] = {-9'd88,-10'd88};
ram[31584] = {-9'd85,-10'd85};
ram[31585] = {-9'd82,-10'd82};
ram[31586] = {-9'd79,-10'd79};
ram[31587] = {-9'd76,-10'd76};
ram[31588] = {-9'd73,-10'd73};
ram[31589] = {-9'd70,-10'd70};
ram[31590] = {-9'd66,-10'd66};
ram[31591] = {-9'd63,-10'd63};
ram[31592] = {-9'd60,-10'd60};
ram[31593] = {-9'd57,-10'd57};
ram[31594] = {-9'd54,-10'd54};
ram[31595] = {-9'd51,-10'd51};
ram[31596] = {-9'd48,-10'd48};
ram[31597] = {-9'd44,-10'd44};
ram[31598] = {-9'd41,-10'd41};
ram[31599] = {-9'd38,-10'd38};
ram[31600] = {-9'd35,-10'd35};
ram[31601] = {-9'd32,-10'd32};
ram[31602] = {-9'd29,-10'd29};
ram[31603] = {-9'd26,-10'd26};
ram[31604] = {-9'd22,-10'd22};
ram[31605] = {-9'd19,-10'd19};
ram[31606] = {-9'd16,-10'd16};
ram[31607] = {-9'd13,-10'd13};
ram[31608] = {-9'd10,-10'd10};
ram[31609] = {-9'd7,-10'd7};
ram[31610] = {-9'd4,-10'd4};
ram[31611] = {9'd0,10'd0};
ram[31612] = {9'd3,10'd3};
ram[31613] = {9'd6,10'd6};
ram[31614] = {9'd9,10'd9};
ram[31615] = {9'd12,10'd12};
ram[31616] = {9'd12,10'd12};
ram[31617] = {9'd15,10'd15};
ram[31618] = {9'd18,10'd18};
ram[31619] = {9'd21,10'd21};
ram[31620] = {9'd25,10'd25};
ram[31621] = {9'd28,10'd28};
ram[31622] = {9'd31,10'd31};
ram[31623] = {9'd34,10'd34};
ram[31624] = {9'd37,10'd37};
ram[31625] = {9'd40,10'd40};
ram[31626] = {9'd43,10'd43};
ram[31627] = {9'd47,10'd47};
ram[31628] = {9'd50,10'd50};
ram[31629] = {9'd53,10'd53};
ram[31630] = {9'd56,10'd56};
ram[31631] = {9'd59,10'd59};
ram[31632] = {9'd62,10'd62};
ram[31633] = {9'd65,10'd65};
ram[31634] = {9'd69,10'd69};
ram[31635] = {9'd72,10'd72};
ram[31636] = {9'd75,10'd75};
ram[31637] = {9'd78,10'd78};
ram[31638] = {9'd81,10'd81};
ram[31639] = {9'd84,10'd84};
ram[31640] = {9'd87,10'd87};
ram[31641] = {9'd91,10'd91};
ram[31642] = {9'd94,10'd94};
ram[31643] = {9'd97,10'd97};
ram[31644] = {-9'd100,10'd100};
ram[31645] = {-9'd97,10'd103};
ram[31646] = {-9'd94,10'd106};
ram[31647] = {-9'd91,10'd109};
ram[31648] = {-9'd88,10'd113};
ram[31649] = {-9'd85,10'd116};
ram[31650] = {-9'd81,10'd119};
ram[31651] = {-9'd78,10'd122};
ram[31652] = {-9'd75,10'd125};
ram[31653] = {-9'd72,10'd128};
ram[31654] = {-9'd69,10'd131};
ram[31655] = {-9'd66,10'd135};
ram[31656] = {-9'd63,10'd138};
ram[31657] = {-9'd59,10'd141};
ram[31658] = {-9'd56,10'd144};
ram[31659] = {-9'd53,10'd147};
ram[31660] = {-9'd50,10'd150};
ram[31661] = {-9'd47,10'd153};
ram[31662] = {-9'd44,10'd157};
ram[31663] = {-9'd41,10'd160};
ram[31664] = {-9'd37,10'd163};
ram[31665] = {-9'd34,10'd166};
ram[31666] = {-9'd31,10'd169};
ram[31667] = {-9'd28,10'd172};
ram[31668] = {-9'd25,10'd175};
ram[31669] = {-9'd22,10'd179};
ram[31670] = {-9'd19,10'd182};
ram[31671] = {-9'd15,10'd185};
ram[31672] = {-9'd12,10'd188};
ram[31673] = {-9'd9,10'd191};
ram[31674] = {-9'd6,10'd194};
ram[31675] = {-9'd3,10'd197};
ram[31676] = {9'd0,10'd201};
ram[31677] = {9'd3,10'd204};
ram[31678] = {9'd7,10'd207};
ram[31679] = {9'd10,10'd210};
ram[31680] = {9'd13,10'd213};
ram[31681] = {9'd16,10'd216};
ram[31682] = {9'd19,10'd219};
ram[31683] = {9'd22,10'd223};
ram[31684] = {9'd25,10'd226};
ram[31685] = {9'd29,10'd229};
ram[31686] = {9'd32,10'd232};
ram[31687] = {9'd35,10'd235};
ram[31688] = {9'd38,10'd238};
ram[31689] = {9'd41,10'd241};
ram[31690] = {9'd44,10'd245};
ram[31691] = {9'd47,10'd248};
ram[31692] = {9'd51,10'd251};
ram[31693] = {9'd54,10'd254};
ram[31694] = {9'd57,10'd257};
ram[31695] = {9'd60,10'd260};
ram[31696] = {9'd63,10'd263};
ram[31697] = {9'd66,10'd267};
ram[31698] = {9'd69,10'd270};
ram[31699] = {9'd73,10'd273};
ram[31700] = {9'd76,10'd276};
ram[31701] = {9'd79,10'd279};
ram[31702] = {9'd82,10'd282};
ram[31703] = {9'd85,10'd285};
ram[31704] = {9'd88,10'd289};
ram[31705] = {9'd91,10'd292};
ram[31706] = {9'd95,10'd295};
ram[31707] = {9'd98,10'd298};
ram[31708] = {-9'd99,10'd301};
ram[31709] = {-9'd96,10'd304};
ram[31710] = {-9'd93,10'd307};
ram[31711] = {-9'd90,10'd311};
ram[31712] = {-9'd87,10'd314};
ram[31713] = {-9'd84,10'd317};
ram[31714] = {-9'd81,10'd320};
ram[31715] = {-9'd77,10'd323};
ram[31716] = {-9'd74,10'd326};
ram[31717] = {-9'd71,10'd329};
ram[31718] = {-9'd68,10'd333};
ram[31719] = {-9'd65,10'd336};
ram[31720] = {-9'd62,10'd339};
ram[31721] = {-9'd59,10'd342};
ram[31722] = {-9'd55,10'd345};
ram[31723] = {-9'd52,10'd348};
ram[31724] = {-9'd49,10'd351};
ram[31725] = {-9'd46,10'd354};
ram[31726] = {-9'd43,10'd358};
ram[31727] = {-9'd40,10'd361};
ram[31728] = {-9'd37,10'd364};
ram[31729] = {-9'd33,10'd367};
ram[31730] = {-9'd30,10'd370};
ram[31731] = {-9'd27,10'd373};
ram[31732] = {-9'd24,10'd376};
ram[31733] = {-9'd21,10'd380};
ram[31734] = {-9'd18,10'd383};
ram[31735] = {-9'd15,10'd386};
ram[31736] = {-9'd11,10'd389};
ram[31737] = {-9'd8,10'd392};
ram[31738] = {-9'd5,10'd395};
ram[31739] = {-9'd2,10'd398};
ram[31740] = {9'd1,-10'd399};
ram[31741] = {9'd4,-10'd396};
ram[31742] = {9'd7,-10'd393};
ram[31743] = {9'd10,-10'd390};
ram[31744] = {9'd10,-10'd390};
ram[31745] = {9'd14,-10'd387};
ram[31746] = {9'd17,-10'd384};
ram[31747] = {9'd20,-10'd381};
ram[31748] = {9'd23,-10'd377};
ram[31749] = {9'd26,-10'd374};
ram[31750] = {9'd29,-10'd371};
ram[31751] = {9'd32,-10'd368};
ram[31752] = {9'd36,-10'd365};
ram[31753] = {9'd39,-10'd362};
ram[31754] = {9'd42,-10'd359};
ram[31755] = {9'd45,-10'd355};
ram[31756] = {9'd48,-10'd352};
ram[31757] = {9'd51,-10'd349};
ram[31758] = {9'd54,-10'd346};
ram[31759] = {9'd58,-10'd343};
ram[31760] = {9'd61,-10'd340};
ram[31761] = {9'd64,-10'd337};
ram[31762] = {9'd67,-10'd334};
ram[31763] = {9'd70,-10'd330};
ram[31764] = {9'd73,-10'd327};
ram[31765] = {9'd76,-10'd324};
ram[31766] = {9'd80,-10'd321};
ram[31767] = {9'd83,-10'd318};
ram[31768] = {9'd86,-10'd315};
ram[31769] = {9'd89,-10'd312};
ram[31770] = {9'd92,-10'd308};
ram[31771] = {9'd95,-10'd305};
ram[31772] = {9'd98,-10'd302};
ram[31773] = {-9'd99,-10'd299};
ram[31774] = {-9'd96,-10'd296};
ram[31775] = {-9'd92,-10'd293};
ram[31776] = {-9'd89,-10'd290};
ram[31777] = {-9'd86,-10'd286};
ram[31778] = {-9'd83,-10'd283};
ram[31779] = {-9'd80,-10'd280};
ram[31780] = {-9'd77,-10'd277};
ram[31781] = {-9'd74,-10'd274};
ram[31782] = {-9'd70,-10'd271};
ram[31783] = {-9'd67,-10'd268};
ram[31784] = {-9'd64,-10'd264};
ram[31785] = {-9'd61,-10'd261};
ram[31786] = {-9'd58,-10'd258};
ram[31787] = {-9'd55,-10'd255};
ram[31788] = {-9'd52,-10'd252};
ram[31789] = {-9'd48,-10'd249};
ram[31790] = {-9'd45,-10'd246};
ram[31791] = {-9'd42,-10'd242};
ram[31792] = {-9'd39,-10'd239};
ram[31793] = {-9'd36,-10'd236};
ram[31794] = {-9'd33,-10'd233};
ram[31795] = {-9'd30,-10'd230};
ram[31796] = {-9'd26,-10'd227};
ram[31797] = {-9'd23,-10'd224};
ram[31798] = {-9'd20,-10'd220};
ram[31799] = {-9'd17,-10'd217};
ram[31800] = {-9'd14,-10'd214};
ram[31801] = {-9'd11,-10'd211};
ram[31802] = {-9'd8,-10'd208};
ram[31803] = {-9'd4,-10'd205};
ram[31804] = {-9'd1,-10'd202};
ram[31805] = {9'd2,-10'd198};
ram[31806] = {9'd5,-10'd195};
ram[31807] = {9'd8,-10'd192};
ram[31808] = {9'd11,-10'd189};
ram[31809] = {9'd14,-10'd186};
ram[31810] = {9'd18,-10'd183};
ram[31811] = {9'd21,-10'd180};
ram[31812] = {9'd24,-10'd176};
ram[31813] = {9'd27,-10'd173};
ram[31814] = {9'd30,-10'd170};
ram[31815] = {9'd33,-10'd167};
ram[31816] = {9'd36,-10'd164};
ram[31817] = {9'd40,-10'd161};
ram[31818] = {9'd43,-10'd158};
ram[31819] = {9'd46,-10'd154};
ram[31820] = {9'd49,-10'd151};
ram[31821] = {9'd52,-10'd148};
ram[31822] = {9'd55,-10'd145};
ram[31823] = {9'd58,-10'd142};
ram[31824] = {9'd62,-10'd139};
ram[31825] = {9'd65,-10'd136};
ram[31826] = {9'd68,-10'd132};
ram[31827] = {9'd71,-10'd129};
ram[31828] = {9'd74,-10'd126};
ram[31829] = {9'd77,-10'd123};
ram[31830] = {9'd80,-10'd120};
ram[31831] = {9'd84,-10'd117};
ram[31832] = {9'd87,-10'd114};
ram[31833] = {9'd90,-10'd110};
ram[31834] = {9'd93,-10'd107};
ram[31835] = {9'd96,-10'd104};
ram[31836] = {9'd99,-10'd101};
ram[31837] = {-9'd98,-10'd98};
ram[31838] = {-9'd95,-10'd95};
ram[31839] = {-9'd92,-10'd92};
ram[31840] = {-9'd88,-10'd88};
ram[31841] = {-9'd85,-10'd85};
ram[31842] = {-9'd82,-10'd82};
ram[31843] = {-9'd79,-10'd79};
ram[31844] = {-9'd76,-10'd76};
ram[31845] = {-9'd73,-10'd73};
ram[31846] = {-9'd70,-10'd70};
ram[31847] = {-9'd66,-10'd66};
ram[31848] = {-9'd63,-10'd63};
ram[31849] = {-9'd60,-10'd60};
ram[31850] = {-9'd57,-10'd57};
ram[31851] = {-9'd54,-10'd54};
ram[31852] = {-9'd51,-10'd51};
ram[31853] = {-9'd48,-10'd48};
ram[31854] = {-9'd44,-10'd44};
ram[31855] = {-9'd41,-10'd41};
ram[31856] = {-9'd38,-10'd38};
ram[31857] = {-9'd35,-10'd35};
ram[31858] = {-9'd32,-10'd32};
ram[31859] = {-9'd29,-10'd29};
ram[31860] = {-9'd26,-10'd26};
ram[31861] = {-9'd22,-10'd22};
ram[31862] = {-9'd19,-10'd19};
ram[31863] = {-9'd16,-10'd16};
ram[31864] = {-9'd13,-10'd13};
ram[31865] = {-9'd10,-10'd10};
ram[31866] = {-9'd7,-10'd7};
ram[31867] = {-9'd4,-10'd4};
ram[31868] = {9'd0,10'd0};
ram[31869] = {9'd3,10'd3};
ram[31870] = {9'd6,10'd6};
ram[31871] = {9'd9,10'd9};
ram[31872] = {9'd9,10'd9};
ram[31873] = {9'd12,10'd12};
ram[31874] = {9'd15,10'd15};
ram[31875] = {9'd18,10'd18};
ram[31876] = {9'd21,10'd21};
ram[31877] = {9'd25,10'd25};
ram[31878] = {9'd28,10'd28};
ram[31879] = {9'd31,10'd31};
ram[31880] = {9'd34,10'd34};
ram[31881] = {9'd37,10'd37};
ram[31882] = {9'd40,10'd40};
ram[31883] = {9'd43,10'd43};
ram[31884] = {9'd47,10'd47};
ram[31885] = {9'd50,10'd50};
ram[31886] = {9'd53,10'd53};
ram[31887] = {9'd56,10'd56};
ram[31888] = {9'd59,10'd59};
ram[31889] = {9'd62,10'd62};
ram[31890] = {9'd65,10'd65};
ram[31891] = {9'd69,10'd69};
ram[31892] = {9'd72,10'd72};
ram[31893] = {9'd75,10'd75};
ram[31894] = {9'd78,10'd78};
ram[31895] = {9'd81,10'd81};
ram[31896] = {9'd84,10'd84};
ram[31897] = {9'd87,10'd87};
ram[31898] = {9'd91,10'd91};
ram[31899] = {9'd94,10'd94};
ram[31900] = {9'd97,10'd97};
ram[31901] = {-9'd100,10'd100};
ram[31902] = {-9'd97,10'd103};
ram[31903] = {-9'd94,10'd106};
ram[31904] = {-9'd91,10'd109};
ram[31905] = {-9'd88,10'd113};
ram[31906] = {-9'd85,10'd116};
ram[31907] = {-9'd81,10'd119};
ram[31908] = {-9'd78,10'd122};
ram[31909] = {-9'd75,10'd125};
ram[31910] = {-9'd72,10'd128};
ram[31911] = {-9'd69,10'd131};
ram[31912] = {-9'd66,10'd135};
ram[31913] = {-9'd63,10'd138};
ram[31914] = {-9'd59,10'd141};
ram[31915] = {-9'd56,10'd144};
ram[31916] = {-9'd53,10'd147};
ram[31917] = {-9'd50,10'd150};
ram[31918] = {-9'd47,10'd153};
ram[31919] = {-9'd44,10'd157};
ram[31920] = {-9'd41,10'd160};
ram[31921] = {-9'd37,10'd163};
ram[31922] = {-9'd34,10'd166};
ram[31923] = {-9'd31,10'd169};
ram[31924] = {-9'd28,10'd172};
ram[31925] = {-9'd25,10'd175};
ram[31926] = {-9'd22,10'd179};
ram[31927] = {-9'd19,10'd182};
ram[31928] = {-9'd15,10'd185};
ram[31929] = {-9'd12,10'd188};
ram[31930] = {-9'd9,10'd191};
ram[31931] = {-9'd6,10'd194};
ram[31932] = {-9'd3,10'd197};
ram[31933] = {9'd0,10'd201};
ram[31934] = {9'd3,10'd204};
ram[31935] = {9'd7,10'd207};
ram[31936] = {9'd10,10'd210};
ram[31937] = {9'd13,10'd213};
ram[31938] = {9'd16,10'd216};
ram[31939] = {9'd19,10'd219};
ram[31940] = {9'd22,10'd223};
ram[31941] = {9'd25,10'd226};
ram[31942] = {9'd29,10'd229};
ram[31943] = {9'd32,10'd232};
ram[31944] = {9'd35,10'd235};
ram[31945] = {9'd38,10'd238};
ram[31946] = {9'd41,10'd241};
ram[31947] = {9'd44,10'd245};
ram[31948] = {9'd47,10'd248};
ram[31949] = {9'd51,10'd251};
ram[31950] = {9'd54,10'd254};
ram[31951] = {9'd57,10'd257};
ram[31952] = {9'd60,10'd260};
ram[31953] = {9'd63,10'd263};
ram[31954] = {9'd66,10'd267};
ram[31955] = {9'd69,10'd270};
ram[31956] = {9'd73,10'd273};
ram[31957] = {9'd76,10'd276};
ram[31958] = {9'd79,10'd279};
ram[31959] = {9'd82,10'd282};
ram[31960] = {9'd85,10'd285};
ram[31961] = {9'd88,10'd289};
ram[31962] = {9'd91,10'd292};
ram[31963] = {9'd95,10'd295};
ram[31964] = {9'd98,10'd298};
ram[31965] = {-9'd99,10'd301};
ram[31966] = {-9'd96,10'd304};
ram[31967] = {-9'd93,10'd307};
ram[31968] = {-9'd90,10'd311};
ram[31969] = {-9'd87,10'd314};
ram[31970] = {-9'd84,10'd317};
ram[31971] = {-9'd81,10'd320};
ram[31972] = {-9'd77,10'd323};
ram[31973] = {-9'd74,10'd326};
ram[31974] = {-9'd71,10'd329};
ram[31975] = {-9'd68,10'd333};
ram[31976] = {-9'd65,10'd336};
ram[31977] = {-9'd62,10'd339};
ram[31978] = {-9'd59,10'd342};
ram[31979] = {-9'd55,10'd345};
ram[31980] = {-9'd52,10'd348};
ram[31981] = {-9'd49,10'd351};
ram[31982] = {-9'd46,10'd354};
ram[31983] = {-9'd43,10'd358};
ram[31984] = {-9'd40,10'd361};
ram[31985] = {-9'd37,10'd364};
ram[31986] = {-9'd33,10'd367};
ram[31987] = {-9'd30,10'd370};
ram[31988] = {-9'd27,10'd373};
ram[31989] = {-9'd24,10'd376};
ram[31990] = {-9'd21,10'd380};
ram[31991] = {-9'd18,10'd383};
ram[31992] = {-9'd15,10'd386};
ram[31993] = {-9'd11,10'd389};
ram[31994] = {-9'd8,10'd392};
ram[31995] = {-9'd5,10'd395};
ram[31996] = {-9'd2,10'd398};
ram[31997] = {9'd1,-10'd399};
ram[31998] = {9'd4,-10'd396};
ram[31999] = {9'd7,-10'd393};
ram[32000] = {9'd7,-10'd393};
ram[32001] = {9'd10,-10'd390};
ram[32002] = {9'd14,-10'd387};
ram[32003] = {9'd17,-10'd384};
ram[32004] = {9'd20,-10'd381};
ram[32005] = {9'd23,-10'd377};
ram[32006] = {9'd26,-10'd374};
ram[32007] = {9'd29,-10'd371};
ram[32008] = {9'd32,-10'd368};
ram[32009] = {9'd36,-10'd365};
ram[32010] = {9'd39,-10'd362};
ram[32011] = {9'd42,-10'd359};
ram[32012] = {9'd45,-10'd355};
ram[32013] = {9'd48,-10'd352};
ram[32014] = {9'd51,-10'd349};
ram[32015] = {9'd54,-10'd346};
ram[32016] = {9'd58,-10'd343};
ram[32017] = {9'd61,-10'd340};
ram[32018] = {9'd64,-10'd337};
ram[32019] = {9'd67,-10'd334};
ram[32020] = {9'd70,-10'd330};
ram[32021] = {9'd73,-10'd327};
ram[32022] = {9'd76,-10'd324};
ram[32023] = {9'd80,-10'd321};
ram[32024] = {9'd83,-10'd318};
ram[32025] = {9'd86,-10'd315};
ram[32026] = {9'd89,-10'd312};
ram[32027] = {9'd92,-10'd308};
ram[32028] = {9'd95,-10'd305};
ram[32029] = {9'd98,-10'd302};
ram[32030] = {-9'd99,-10'd299};
ram[32031] = {-9'd96,-10'd296};
ram[32032] = {-9'd92,-10'd293};
ram[32033] = {-9'd89,-10'd290};
ram[32034] = {-9'd86,-10'd286};
ram[32035] = {-9'd83,-10'd283};
ram[32036] = {-9'd80,-10'd280};
ram[32037] = {-9'd77,-10'd277};
ram[32038] = {-9'd74,-10'd274};
ram[32039] = {-9'd70,-10'd271};
ram[32040] = {-9'd67,-10'd268};
ram[32041] = {-9'd64,-10'd264};
ram[32042] = {-9'd61,-10'd261};
ram[32043] = {-9'd58,-10'd258};
ram[32044] = {-9'd55,-10'd255};
ram[32045] = {-9'd52,-10'd252};
ram[32046] = {-9'd48,-10'd249};
ram[32047] = {-9'd45,-10'd246};
ram[32048] = {-9'd42,-10'd242};
ram[32049] = {-9'd39,-10'd239};
ram[32050] = {-9'd36,-10'd236};
ram[32051] = {-9'd33,-10'd233};
ram[32052] = {-9'd30,-10'd230};
ram[32053] = {-9'd26,-10'd227};
ram[32054] = {-9'd23,-10'd224};
ram[32055] = {-9'd20,-10'd220};
ram[32056] = {-9'd17,-10'd217};
ram[32057] = {-9'd14,-10'd214};
ram[32058] = {-9'd11,-10'd211};
ram[32059] = {-9'd8,-10'd208};
ram[32060] = {-9'd4,-10'd205};
ram[32061] = {-9'd1,-10'd202};
ram[32062] = {9'd2,-10'd198};
ram[32063] = {9'd5,-10'd195};
ram[32064] = {9'd8,-10'd192};
ram[32065] = {9'd11,-10'd189};
ram[32066] = {9'd14,-10'd186};
ram[32067] = {9'd18,-10'd183};
ram[32068] = {9'd21,-10'd180};
ram[32069] = {9'd24,-10'd176};
ram[32070] = {9'd27,-10'd173};
ram[32071] = {9'd30,-10'd170};
ram[32072] = {9'd33,-10'd167};
ram[32073] = {9'd36,-10'd164};
ram[32074] = {9'd40,-10'd161};
ram[32075] = {9'd43,-10'd158};
ram[32076] = {9'd46,-10'd154};
ram[32077] = {9'd49,-10'd151};
ram[32078] = {9'd52,-10'd148};
ram[32079] = {9'd55,-10'd145};
ram[32080] = {9'd58,-10'd142};
ram[32081] = {9'd62,-10'd139};
ram[32082] = {9'd65,-10'd136};
ram[32083] = {9'd68,-10'd132};
ram[32084] = {9'd71,-10'd129};
ram[32085] = {9'd74,-10'd126};
ram[32086] = {9'd77,-10'd123};
ram[32087] = {9'd80,-10'd120};
ram[32088] = {9'd84,-10'd117};
ram[32089] = {9'd87,-10'd114};
ram[32090] = {9'd90,-10'd110};
ram[32091] = {9'd93,-10'd107};
ram[32092] = {9'd96,-10'd104};
ram[32093] = {9'd99,-10'd101};
ram[32094] = {-9'd98,-10'd98};
ram[32095] = {-9'd95,-10'd95};
ram[32096] = {-9'd92,-10'd92};
ram[32097] = {-9'd88,-10'd88};
ram[32098] = {-9'd85,-10'd85};
ram[32099] = {-9'd82,-10'd82};
ram[32100] = {-9'd79,-10'd79};
ram[32101] = {-9'd76,-10'd76};
ram[32102] = {-9'd73,-10'd73};
ram[32103] = {-9'd70,-10'd70};
ram[32104] = {-9'd66,-10'd66};
ram[32105] = {-9'd63,-10'd63};
ram[32106] = {-9'd60,-10'd60};
ram[32107] = {-9'd57,-10'd57};
ram[32108] = {-9'd54,-10'd54};
ram[32109] = {-9'd51,-10'd51};
ram[32110] = {-9'd48,-10'd48};
ram[32111] = {-9'd44,-10'd44};
ram[32112] = {-9'd41,-10'd41};
ram[32113] = {-9'd38,-10'd38};
ram[32114] = {-9'd35,-10'd35};
ram[32115] = {-9'd32,-10'd32};
ram[32116] = {-9'd29,-10'd29};
ram[32117] = {-9'd26,-10'd26};
ram[32118] = {-9'd22,-10'd22};
ram[32119] = {-9'd19,-10'd19};
ram[32120] = {-9'd16,-10'd16};
ram[32121] = {-9'd13,-10'd13};
ram[32122] = {-9'd10,-10'd10};
ram[32123] = {-9'd7,-10'd7};
ram[32124] = {-9'd4,-10'd4};
ram[32125] = {9'd0,10'd0};
ram[32126] = {9'd3,10'd3};
ram[32127] = {9'd6,10'd6};
ram[32128] = {9'd6,10'd6};
ram[32129] = {9'd9,10'd9};
ram[32130] = {9'd12,10'd12};
ram[32131] = {9'd15,10'd15};
ram[32132] = {9'd18,10'd18};
ram[32133] = {9'd21,10'd21};
ram[32134] = {9'd25,10'd25};
ram[32135] = {9'd28,10'd28};
ram[32136] = {9'd31,10'd31};
ram[32137] = {9'd34,10'd34};
ram[32138] = {9'd37,10'd37};
ram[32139] = {9'd40,10'd40};
ram[32140] = {9'd43,10'd43};
ram[32141] = {9'd47,10'd47};
ram[32142] = {9'd50,10'd50};
ram[32143] = {9'd53,10'd53};
ram[32144] = {9'd56,10'd56};
ram[32145] = {9'd59,10'd59};
ram[32146] = {9'd62,10'd62};
ram[32147] = {9'd65,10'd65};
ram[32148] = {9'd69,10'd69};
ram[32149] = {9'd72,10'd72};
ram[32150] = {9'd75,10'd75};
ram[32151] = {9'd78,10'd78};
ram[32152] = {9'd81,10'd81};
ram[32153] = {9'd84,10'd84};
ram[32154] = {9'd87,10'd87};
ram[32155] = {9'd91,10'd91};
ram[32156] = {9'd94,10'd94};
ram[32157] = {9'd97,10'd97};
ram[32158] = {-9'd100,10'd100};
ram[32159] = {-9'd97,10'd103};
ram[32160] = {-9'd94,10'd106};
ram[32161] = {-9'd91,10'd109};
ram[32162] = {-9'd88,10'd113};
ram[32163] = {-9'd85,10'd116};
ram[32164] = {-9'd81,10'd119};
ram[32165] = {-9'd78,10'd122};
ram[32166] = {-9'd75,10'd125};
ram[32167] = {-9'd72,10'd128};
ram[32168] = {-9'd69,10'd131};
ram[32169] = {-9'd66,10'd135};
ram[32170] = {-9'd63,10'd138};
ram[32171] = {-9'd59,10'd141};
ram[32172] = {-9'd56,10'd144};
ram[32173] = {-9'd53,10'd147};
ram[32174] = {-9'd50,10'd150};
ram[32175] = {-9'd47,10'd153};
ram[32176] = {-9'd44,10'd157};
ram[32177] = {-9'd41,10'd160};
ram[32178] = {-9'd37,10'd163};
ram[32179] = {-9'd34,10'd166};
ram[32180] = {-9'd31,10'd169};
ram[32181] = {-9'd28,10'd172};
ram[32182] = {-9'd25,10'd175};
ram[32183] = {-9'd22,10'd179};
ram[32184] = {-9'd19,10'd182};
ram[32185] = {-9'd15,10'd185};
ram[32186] = {-9'd12,10'd188};
ram[32187] = {-9'd9,10'd191};
ram[32188] = {-9'd6,10'd194};
ram[32189] = {-9'd3,10'd197};
ram[32190] = {9'd0,10'd201};
ram[32191] = {9'd3,10'd204};
ram[32192] = {9'd7,10'd207};
ram[32193] = {9'd10,10'd210};
ram[32194] = {9'd13,10'd213};
ram[32195] = {9'd16,10'd216};
ram[32196] = {9'd19,10'd219};
ram[32197] = {9'd22,10'd223};
ram[32198] = {9'd25,10'd226};
ram[32199] = {9'd29,10'd229};
ram[32200] = {9'd32,10'd232};
ram[32201] = {9'd35,10'd235};
ram[32202] = {9'd38,10'd238};
ram[32203] = {9'd41,10'd241};
ram[32204] = {9'd44,10'd245};
ram[32205] = {9'd47,10'd248};
ram[32206] = {9'd51,10'd251};
ram[32207] = {9'd54,10'd254};
ram[32208] = {9'd57,10'd257};
ram[32209] = {9'd60,10'd260};
ram[32210] = {9'd63,10'd263};
ram[32211] = {9'd66,10'd267};
ram[32212] = {9'd69,10'd270};
ram[32213] = {9'd73,10'd273};
ram[32214] = {9'd76,10'd276};
ram[32215] = {9'd79,10'd279};
ram[32216] = {9'd82,10'd282};
ram[32217] = {9'd85,10'd285};
ram[32218] = {9'd88,10'd289};
ram[32219] = {9'd91,10'd292};
ram[32220] = {9'd95,10'd295};
ram[32221] = {9'd98,10'd298};
ram[32222] = {-9'd99,10'd301};
ram[32223] = {-9'd96,10'd304};
ram[32224] = {-9'd93,10'd307};
ram[32225] = {-9'd90,10'd311};
ram[32226] = {-9'd87,10'd314};
ram[32227] = {-9'd84,10'd317};
ram[32228] = {-9'd81,10'd320};
ram[32229] = {-9'd77,10'd323};
ram[32230] = {-9'd74,10'd326};
ram[32231] = {-9'd71,10'd329};
ram[32232] = {-9'd68,10'd333};
ram[32233] = {-9'd65,10'd336};
ram[32234] = {-9'd62,10'd339};
ram[32235] = {-9'd59,10'd342};
ram[32236] = {-9'd55,10'd345};
ram[32237] = {-9'd52,10'd348};
ram[32238] = {-9'd49,10'd351};
ram[32239] = {-9'd46,10'd354};
ram[32240] = {-9'd43,10'd358};
ram[32241] = {-9'd40,10'd361};
ram[32242] = {-9'd37,10'd364};
ram[32243] = {-9'd33,10'd367};
ram[32244] = {-9'd30,10'd370};
ram[32245] = {-9'd27,10'd373};
ram[32246] = {-9'd24,10'd376};
ram[32247] = {-9'd21,10'd380};
ram[32248] = {-9'd18,10'd383};
ram[32249] = {-9'd15,10'd386};
ram[32250] = {-9'd11,10'd389};
ram[32251] = {-9'd8,10'd392};
ram[32252] = {-9'd5,10'd395};
ram[32253] = {-9'd2,10'd398};
ram[32254] = {9'd1,-10'd399};
ram[32255] = {9'd4,-10'd396};
ram[32256] = {9'd4,-10'd396};
ram[32257] = {9'd7,-10'd393};
ram[32258] = {9'd10,-10'd390};
ram[32259] = {9'd14,-10'd387};
ram[32260] = {9'd17,-10'd384};
ram[32261] = {9'd20,-10'd381};
ram[32262] = {9'd23,-10'd377};
ram[32263] = {9'd26,-10'd374};
ram[32264] = {9'd29,-10'd371};
ram[32265] = {9'd32,-10'd368};
ram[32266] = {9'd36,-10'd365};
ram[32267] = {9'd39,-10'd362};
ram[32268] = {9'd42,-10'd359};
ram[32269] = {9'd45,-10'd355};
ram[32270] = {9'd48,-10'd352};
ram[32271] = {9'd51,-10'd349};
ram[32272] = {9'd54,-10'd346};
ram[32273] = {9'd58,-10'd343};
ram[32274] = {9'd61,-10'd340};
ram[32275] = {9'd64,-10'd337};
ram[32276] = {9'd67,-10'd334};
ram[32277] = {9'd70,-10'd330};
ram[32278] = {9'd73,-10'd327};
ram[32279] = {9'd76,-10'd324};
ram[32280] = {9'd80,-10'd321};
ram[32281] = {9'd83,-10'd318};
ram[32282] = {9'd86,-10'd315};
ram[32283] = {9'd89,-10'd312};
ram[32284] = {9'd92,-10'd308};
ram[32285] = {9'd95,-10'd305};
ram[32286] = {9'd98,-10'd302};
ram[32287] = {-9'd99,-10'd299};
ram[32288] = {-9'd96,-10'd296};
ram[32289] = {-9'd92,-10'd293};
ram[32290] = {-9'd89,-10'd290};
ram[32291] = {-9'd86,-10'd286};
ram[32292] = {-9'd83,-10'd283};
ram[32293] = {-9'd80,-10'd280};
ram[32294] = {-9'd77,-10'd277};
ram[32295] = {-9'd74,-10'd274};
ram[32296] = {-9'd70,-10'd271};
ram[32297] = {-9'd67,-10'd268};
ram[32298] = {-9'd64,-10'd264};
ram[32299] = {-9'd61,-10'd261};
ram[32300] = {-9'd58,-10'd258};
ram[32301] = {-9'd55,-10'd255};
ram[32302] = {-9'd52,-10'd252};
ram[32303] = {-9'd48,-10'd249};
ram[32304] = {-9'd45,-10'd246};
ram[32305] = {-9'd42,-10'd242};
ram[32306] = {-9'd39,-10'd239};
ram[32307] = {-9'd36,-10'd236};
ram[32308] = {-9'd33,-10'd233};
ram[32309] = {-9'd30,-10'd230};
ram[32310] = {-9'd26,-10'd227};
ram[32311] = {-9'd23,-10'd224};
ram[32312] = {-9'd20,-10'd220};
ram[32313] = {-9'd17,-10'd217};
ram[32314] = {-9'd14,-10'd214};
ram[32315] = {-9'd11,-10'd211};
ram[32316] = {-9'd8,-10'd208};
ram[32317] = {-9'd4,-10'd205};
ram[32318] = {-9'd1,-10'd202};
ram[32319] = {9'd2,-10'd198};
ram[32320] = {9'd5,-10'd195};
ram[32321] = {9'd8,-10'd192};
ram[32322] = {9'd11,-10'd189};
ram[32323] = {9'd14,-10'd186};
ram[32324] = {9'd18,-10'd183};
ram[32325] = {9'd21,-10'd180};
ram[32326] = {9'd24,-10'd176};
ram[32327] = {9'd27,-10'd173};
ram[32328] = {9'd30,-10'd170};
ram[32329] = {9'd33,-10'd167};
ram[32330] = {9'd36,-10'd164};
ram[32331] = {9'd40,-10'd161};
ram[32332] = {9'd43,-10'd158};
ram[32333] = {9'd46,-10'd154};
ram[32334] = {9'd49,-10'd151};
ram[32335] = {9'd52,-10'd148};
ram[32336] = {9'd55,-10'd145};
ram[32337] = {9'd58,-10'd142};
ram[32338] = {9'd62,-10'd139};
ram[32339] = {9'd65,-10'd136};
ram[32340] = {9'd68,-10'd132};
ram[32341] = {9'd71,-10'd129};
ram[32342] = {9'd74,-10'd126};
ram[32343] = {9'd77,-10'd123};
ram[32344] = {9'd80,-10'd120};
ram[32345] = {9'd84,-10'd117};
ram[32346] = {9'd87,-10'd114};
ram[32347] = {9'd90,-10'd110};
ram[32348] = {9'd93,-10'd107};
ram[32349] = {9'd96,-10'd104};
ram[32350] = {9'd99,-10'd101};
ram[32351] = {-9'd98,-10'd98};
ram[32352] = {-9'd95,-10'd95};
ram[32353] = {-9'd92,-10'd92};
ram[32354] = {-9'd88,-10'd88};
ram[32355] = {-9'd85,-10'd85};
ram[32356] = {-9'd82,-10'd82};
ram[32357] = {-9'd79,-10'd79};
ram[32358] = {-9'd76,-10'd76};
ram[32359] = {-9'd73,-10'd73};
ram[32360] = {-9'd70,-10'd70};
ram[32361] = {-9'd66,-10'd66};
ram[32362] = {-9'd63,-10'd63};
ram[32363] = {-9'd60,-10'd60};
ram[32364] = {-9'd57,-10'd57};
ram[32365] = {-9'd54,-10'd54};
ram[32366] = {-9'd51,-10'd51};
ram[32367] = {-9'd48,-10'd48};
ram[32368] = {-9'd44,-10'd44};
ram[32369] = {-9'd41,-10'd41};
ram[32370] = {-9'd38,-10'd38};
ram[32371] = {-9'd35,-10'd35};
ram[32372] = {-9'd32,-10'd32};
ram[32373] = {-9'd29,-10'd29};
ram[32374] = {-9'd26,-10'd26};
ram[32375] = {-9'd22,-10'd22};
ram[32376] = {-9'd19,-10'd19};
ram[32377] = {-9'd16,-10'd16};
ram[32378] = {-9'd13,-10'd13};
ram[32379] = {-9'd10,-10'd10};
ram[32380] = {-9'd7,-10'd7};
ram[32381] = {-9'd4,-10'd4};
ram[32382] = {9'd0,10'd0};
ram[32383] = {9'd3,10'd3};
ram[32384] = {9'd3,10'd3};
ram[32385] = {9'd6,10'd6};
ram[32386] = {9'd9,10'd9};
ram[32387] = {9'd12,10'd12};
ram[32388] = {9'd15,10'd15};
ram[32389] = {9'd18,10'd18};
ram[32390] = {9'd21,10'd21};
ram[32391] = {9'd25,10'd25};
ram[32392] = {9'd28,10'd28};
ram[32393] = {9'd31,10'd31};
ram[32394] = {9'd34,10'd34};
ram[32395] = {9'd37,10'd37};
ram[32396] = {9'd40,10'd40};
ram[32397] = {9'd43,10'd43};
ram[32398] = {9'd47,10'd47};
ram[32399] = {9'd50,10'd50};
ram[32400] = {9'd53,10'd53};
ram[32401] = {9'd56,10'd56};
ram[32402] = {9'd59,10'd59};
ram[32403] = {9'd62,10'd62};
ram[32404] = {9'd65,10'd65};
ram[32405] = {9'd69,10'd69};
ram[32406] = {9'd72,10'd72};
ram[32407] = {9'd75,10'd75};
ram[32408] = {9'd78,10'd78};
ram[32409] = {9'd81,10'd81};
ram[32410] = {9'd84,10'd84};
ram[32411] = {9'd87,10'd87};
ram[32412] = {9'd91,10'd91};
ram[32413] = {9'd94,10'd94};
ram[32414] = {9'd97,10'd97};
ram[32415] = {-9'd100,10'd100};
ram[32416] = {-9'd97,10'd103};
ram[32417] = {-9'd94,10'd106};
ram[32418] = {-9'd91,10'd109};
ram[32419] = {-9'd88,10'd113};
ram[32420] = {-9'd85,10'd116};
ram[32421] = {-9'd81,10'd119};
ram[32422] = {-9'd78,10'd122};
ram[32423] = {-9'd75,10'd125};
ram[32424] = {-9'd72,10'd128};
ram[32425] = {-9'd69,10'd131};
ram[32426] = {-9'd66,10'd135};
ram[32427] = {-9'd63,10'd138};
ram[32428] = {-9'd59,10'd141};
ram[32429] = {-9'd56,10'd144};
ram[32430] = {-9'd53,10'd147};
ram[32431] = {-9'd50,10'd150};
ram[32432] = {-9'd47,10'd153};
ram[32433] = {-9'd44,10'd157};
ram[32434] = {-9'd41,10'd160};
ram[32435] = {-9'd37,10'd163};
ram[32436] = {-9'd34,10'd166};
ram[32437] = {-9'd31,10'd169};
ram[32438] = {-9'd28,10'd172};
ram[32439] = {-9'd25,10'd175};
ram[32440] = {-9'd22,10'd179};
ram[32441] = {-9'd19,10'd182};
ram[32442] = {-9'd15,10'd185};
ram[32443] = {-9'd12,10'd188};
ram[32444] = {-9'd9,10'd191};
ram[32445] = {-9'd6,10'd194};
ram[32446] = {-9'd3,10'd197};
ram[32447] = {9'd0,10'd201};
ram[32448] = {9'd3,10'd204};
ram[32449] = {9'd7,10'd207};
ram[32450] = {9'd10,10'd210};
ram[32451] = {9'd13,10'd213};
ram[32452] = {9'd16,10'd216};
ram[32453] = {9'd19,10'd219};
ram[32454] = {9'd22,10'd223};
ram[32455] = {9'd25,10'd226};
ram[32456] = {9'd29,10'd229};
ram[32457] = {9'd32,10'd232};
ram[32458] = {9'd35,10'd235};
ram[32459] = {9'd38,10'd238};
ram[32460] = {9'd41,10'd241};
ram[32461] = {9'd44,10'd245};
ram[32462] = {9'd47,10'd248};
ram[32463] = {9'd51,10'd251};
ram[32464] = {9'd54,10'd254};
ram[32465] = {9'd57,10'd257};
ram[32466] = {9'd60,10'd260};
ram[32467] = {9'd63,10'd263};
ram[32468] = {9'd66,10'd267};
ram[32469] = {9'd69,10'd270};
ram[32470] = {9'd73,10'd273};
ram[32471] = {9'd76,10'd276};
ram[32472] = {9'd79,10'd279};
ram[32473] = {9'd82,10'd282};
ram[32474] = {9'd85,10'd285};
ram[32475] = {9'd88,10'd289};
ram[32476] = {9'd91,10'd292};
ram[32477] = {9'd95,10'd295};
ram[32478] = {9'd98,10'd298};
ram[32479] = {-9'd99,10'd301};
ram[32480] = {-9'd96,10'd304};
ram[32481] = {-9'd93,10'd307};
ram[32482] = {-9'd90,10'd311};
ram[32483] = {-9'd87,10'd314};
ram[32484] = {-9'd84,10'd317};
ram[32485] = {-9'd81,10'd320};
ram[32486] = {-9'd77,10'd323};
ram[32487] = {-9'd74,10'd326};
ram[32488] = {-9'd71,10'd329};
ram[32489] = {-9'd68,10'd333};
ram[32490] = {-9'd65,10'd336};
ram[32491] = {-9'd62,10'd339};
ram[32492] = {-9'd59,10'd342};
ram[32493] = {-9'd55,10'd345};
ram[32494] = {-9'd52,10'd348};
ram[32495] = {-9'd49,10'd351};
ram[32496] = {-9'd46,10'd354};
ram[32497] = {-9'd43,10'd358};
ram[32498] = {-9'd40,10'd361};
ram[32499] = {-9'd37,10'd364};
ram[32500] = {-9'd33,10'd367};
ram[32501] = {-9'd30,10'd370};
ram[32502] = {-9'd27,10'd373};
ram[32503] = {-9'd24,10'd376};
ram[32504] = {-9'd21,10'd380};
ram[32505] = {-9'd18,10'd383};
ram[32506] = {-9'd15,10'd386};
ram[32507] = {-9'd11,10'd389};
ram[32508] = {-9'd8,10'd392};
ram[32509] = {-9'd5,10'd395};
ram[32510] = {-9'd2,10'd398};
ram[32511] = {9'd1,-10'd399};
ram[32512] = {9'd1,-10'd399};
ram[32513] = {9'd4,-10'd396};
ram[32514] = {9'd7,-10'd393};
ram[32515] = {9'd10,-10'd390};
ram[32516] = {9'd14,-10'd387};
ram[32517] = {9'd17,-10'd384};
ram[32518] = {9'd20,-10'd381};
ram[32519] = {9'd23,-10'd377};
ram[32520] = {9'd26,-10'd374};
ram[32521] = {9'd29,-10'd371};
ram[32522] = {9'd32,-10'd368};
ram[32523] = {9'd36,-10'd365};
ram[32524] = {9'd39,-10'd362};
ram[32525] = {9'd42,-10'd359};
ram[32526] = {9'd45,-10'd355};
ram[32527] = {9'd48,-10'd352};
ram[32528] = {9'd51,-10'd349};
ram[32529] = {9'd54,-10'd346};
ram[32530] = {9'd58,-10'd343};
ram[32531] = {9'd61,-10'd340};
ram[32532] = {9'd64,-10'd337};
ram[32533] = {9'd67,-10'd334};
ram[32534] = {9'd70,-10'd330};
ram[32535] = {9'd73,-10'd327};
ram[32536] = {9'd76,-10'd324};
ram[32537] = {9'd80,-10'd321};
ram[32538] = {9'd83,-10'd318};
ram[32539] = {9'd86,-10'd315};
ram[32540] = {9'd89,-10'd312};
ram[32541] = {9'd92,-10'd308};
ram[32542] = {9'd95,-10'd305};
ram[32543] = {9'd98,-10'd302};
ram[32544] = {-9'd99,-10'd299};
ram[32545] = {-9'd96,-10'd296};
ram[32546] = {-9'd92,-10'd293};
ram[32547] = {-9'd89,-10'd290};
ram[32548] = {-9'd86,-10'd286};
ram[32549] = {-9'd83,-10'd283};
ram[32550] = {-9'd80,-10'd280};
ram[32551] = {-9'd77,-10'd277};
ram[32552] = {-9'd74,-10'd274};
ram[32553] = {-9'd70,-10'd271};
ram[32554] = {-9'd67,-10'd268};
ram[32555] = {-9'd64,-10'd264};
ram[32556] = {-9'd61,-10'd261};
ram[32557] = {-9'd58,-10'd258};
ram[32558] = {-9'd55,-10'd255};
ram[32559] = {-9'd52,-10'd252};
ram[32560] = {-9'd48,-10'd249};
ram[32561] = {-9'd45,-10'd246};
ram[32562] = {-9'd42,-10'd242};
ram[32563] = {-9'd39,-10'd239};
ram[32564] = {-9'd36,-10'd236};
ram[32565] = {-9'd33,-10'd233};
ram[32566] = {-9'd30,-10'd230};
ram[32567] = {-9'd26,-10'd227};
ram[32568] = {-9'd23,-10'd224};
ram[32569] = {-9'd20,-10'd220};
ram[32570] = {-9'd17,-10'd217};
ram[32571] = {-9'd14,-10'd214};
ram[32572] = {-9'd11,-10'd211};
ram[32573] = {-9'd8,-10'd208};
ram[32574] = {-9'd4,-10'd205};
ram[32575] = {-9'd1,-10'd202};
ram[32576] = {9'd2,-10'd198};
ram[32577] = {9'd5,-10'd195};
ram[32578] = {9'd8,-10'd192};
ram[32579] = {9'd11,-10'd189};
ram[32580] = {9'd14,-10'd186};
ram[32581] = {9'd18,-10'd183};
ram[32582] = {9'd21,-10'd180};
ram[32583] = {9'd24,-10'd176};
ram[32584] = {9'd27,-10'd173};
ram[32585] = {9'd30,-10'd170};
ram[32586] = {9'd33,-10'd167};
ram[32587] = {9'd36,-10'd164};
ram[32588] = {9'd40,-10'd161};
ram[32589] = {9'd43,-10'd158};
ram[32590] = {9'd46,-10'd154};
ram[32591] = {9'd49,-10'd151};
ram[32592] = {9'd52,-10'd148};
ram[32593] = {9'd55,-10'd145};
ram[32594] = {9'd58,-10'd142};
ram[32595] = {9'd62,-10'd139};
ram[32596] = {9'd65,-10'd136};
ram[32597] = {9'd68,-10'd132};
ram[32598] = {9'd71,-10'd129};
ram[32599] = {9'd74,-10'd126};
ram[32600] = {9'd77,-10'd123};
ram[32601] = {9'd80,-10'd120};
ram[32602] = {9'd84,-10'd117};
ram[32603] = {9'd87,-10'd114};
ram[32604] = {9'd90,-10'd110};
ram[32605] = {9'd93,-10'd107};
ram[32606] = {9'd96,-10'd104};
ram[32607] = {9'd99,-10'd101};
ram[32608] = {-9'd98,-10'd98};
ram[32609] = {-9'd95,-10'd95};
ram[32610] = {-9'd92,-10'd92};
ram[32611] = {-9'd88,-10'd88};
ram[32612] = {-9'd85,-10'd85};
ram[32613] = {-9'd82,-10'd82};
ram[32614] = {-9'd79,-10'd79};
ram[32615] = {-9'd76,-10'd76};
ram[32616] = {-9'd73,-10'd73};
ram[32617] = {-9'd70,-10'd70};
ram[32618] = {-9'd66,-10'd66};
ram[32619] = {-9'd63,-10'd63};
ram[32620] = {-9'd60,-10'd60};
ram[32621] = {-9'd57,-10'd57};
ram[32622] = {-9'd54,-10'd54};
ram[32623] = {-9'd51,-10'd51};
ram[32624] = {-9'd48,-10'd48};
ram[32625] = {-9'd44,-10'd44};
ram[32626] = {-9'd41,-10'd41};
ram[32627] = {-9'd38,-10'd38};
ram[32628] = {-9'd35,-10'd35};
ram[32629] = {-9'd32,-10'd32};
ram[32630] = {-9'd29,-10'd29};
ram[32631] = {-9'd26,-10'd26};
ram[32632] = {-9'd22,-10'd22};
ram[32633] = {-9'd19,-10'd19};
ram[32634] = {-9'd16,-10'd16};
ram[32635] = {-9'd13,-10'd13};
ram[32636] = {-9'd10,-10'd10};
ram[32637] = {-9'd7,-10'd7};
ram[32638] = {-9'd4,-10'd4};
ram[32639] = {9'd0,10'd0};
ram[32640] = {9'd0,10'd0};
ram[32641] = {9'd3,10'd3};
ram[32642] = {9'd6,10'd6};
ram[32643] = {9'd9,10'd9};
ram[32644] = {9'd12,10'd12};
ram[32645] = {9'd15,10'd15};
ram[32646] = {9'd18,10'd18};
ram[32647] = {9'd21,10'd21};
ram[32648] = {9'd25,10'd25};
ram[32649] = {9'd28,10'd28};
ram[32650] = {9'd31,10'd31};
ram[32651] = {9'd34,10'd34};
ram[32652] = {9'd37,10'd37};
ram[32653] = {9'd40,10'd40};
ram[32654] = {9'd43,10'd43};
ram[32655] = {9'd47,10'd47};
ram[32656] = {9'd50,10'd50};
ram[32657] = {9'd53,10'd53};
ram[32658] = {9'd56,10'd56};
ram[32659] = {9'd59,10'd59};
ram[32660] = {9'd62,10'd62};
ram[32661] = {9'd65,10'd65};
ram[32662] = {9'd69,10'd69};
ram[32663] = {9'd72,10'd72};
ram[32664] = {9'd75,10'd75};
ram[32665] = {9'd78,10'd78};
ram[32666] = {9'd81,10'd81};
ram[32667] = {9'd84,10'd84};
ram[32668] = {9'd87,10'd87};
ram[32669] = {9'd91,10'd91};
ram[32670] = {9'd94,10'd94};
ram[32671] = {9'd97,10'd97};
ram[32672] = {-9'd100,10'd100};
ram[32673] = {-9'd97,10'd103};
ram[32674] = {-9'd94,10'd106};
ram[32675] = {-9'd91,10'd109};
ram[32676] = {-9'd88,10'd113};
ram[32677] = {-9'd85,10'd116};
ram[32678] = {-9'd81,10'd119};
ram[32679] = {-9'd78,10'd122};
ram[32680] = {-9'd75,10'd125};
ram[32681] = {-9'd72,10'd128};
ram[32682] = {-9'd69,10'd131};
ram[32683] = {-9'd66,10'd135};
ram[32684] = {-9'd63,10'd138};
ram[32685] = {-9'd59,10'd141};
ram[32686] = {-9'd56,10'd144};
ram[32687] = {-9'd53,10'd147};
ram[32688] = {-9'd50,10'd150};
ram[32689] = {-9'd47,10'd153};
ram[32690] = {-9'd44,10'd157};
ram[32691] = {-9'd41,10'd160};
ram[32692] = {-9'd37,10'd163};
ram[32693] = {-9'd34,10'd166};
ram[32694] = {-9'd31,10'd169};
ram[32695] = {-9'd28,10'd172};
ram[32696] = {-9'd25,10'd175};
ram[32697] = {-9'd22,10'd179};
ram[32698] = {-9'd19,10'd182};
ram[32699] = {-9'd15,10'd185};
ram[32700] = {-9'd12,10'd188};
ram[32701] = {-9'd9,10'd191};
ram[32702] = {-9'd6,10'd194};
ram[32703] = {-9'd3,10'd197};
ram[32704] = {9'd0,10'd201};
ram[32705] = {9'd3,10'd204};
ram[32706] = {9'd7,10'd207};
ram[32707] = {9'd10,10'd210};
ram[32708] = {9'd13,10'd213};
ram[32709] = {9'd16,10'd216};
ram[32710] = {9'd19,10'd219};
ram[32711] = {9'd22,10'd223};
ram[32712] = {9'd25,10'd226};
ram[32713] = {9'd29,10'd229};
ram[32714] = {9'd32,10'd232};
ram[32715] = {9'd35,10'd235};
ram[32716] = {9'd38,10'd238};
ram[32717] = {9'd41,10'd241};
ram[32718] = {9'd44,10'd245};
ram[32719] = {9'd47,10'd248};
ram[32720] = {9'd51,10'd251};
ram[32721] = {9'd54,10'd254};
ram[32722] = {9'd57,10'd257};
ram[32723] = {9'd60,10'd260};
ram[32724] = {9'd63,10'd263};
ram[32725] = {9'd66,10'd267};
ram[32726] = {9'd69,10'd270};
ram[32727] = {9'd73,10'd273};
ram[32728] = {9'd76,10'd276};
ram[32729] = {9'd79,10'd279};
ram[32730] = {9'd82,10'd282};
ram[32731] = {9'd85,10'd285};
ram[32732] = {9'd88,10'd289};
ram[32733] = {9'd91,10'd292};
ram[32734] = {9'd95,10'd295};
ram[32735] = {9'd98,10'd298};
ram[32736] = {-9'd99,10'd301};
ram[32737] = {-9'd96,10'd304};
ram[32738] = {-9'd93,10'd307};
ram[32739] = {-9'd90,10'd311};
ram[32740] = {-9'd87,10'd314};
ram[32741] = {-9'd84,10'd317};
ram[32742] = {-9'd81,10'd320};
ram[32743] = {-9'd77,10'd323};
ram[32744] = {-9'd74,10'd326};
ram[32745] = {-9'd71,10'd329};
ram[32746] = {-9'd68,10'd333};
ram[32747] = {-9'd65,10'd336};
ram[32748] = {-9'd62,10'd339};
ram[32749] = {-9'd59,10'd342};
ram[32750] = {-9'd55,10'd345};
ram[32751] = {-9'd52,10'd348};
ram[32752] = {-9'd49,10'd351};
ram[32753] = {-9'd46,10'd354};
ram[32754] = {-9'd43,10'd358};
ram[32755] = {-9'd40,10'd361};
ram[32756] = {-9'd37,10'd364};
ram[32757] = {-9'd33,10'd367};
ram[32758] = {-9'd30,10'd370};
ram[32759] = {-9'd27,10'd373};
ram[32760] = {-9'd24,10'd376};
ram[32761] = {-9'd21,10'd380};
ram[32762] = {-9'd18,10'd383};
ram[32763] = {-9'd15,10'd386};
ram[32764] = {-9'd11,10'd389};
ram[32765] = {-9'd8,10'd392};
ram[32766] = {-9'd5,10'd395};
ram[32767] = {-9'd2,10'd398};
ram[32768] = {-9'd2,10'd398};
ram[32769] = {9'd1,-10'd399};
ram[32770] = {9'd4,-10'd396};
ram[32771] = {9'd7,-10'd393};
ram[32772] = {9'd10,-10'd390};
ram[32773] = {9'd14,-10'd387};
ram[32774] = {9'd17,-10'd384};
ram[32775] = {9'd20,-10'd381};
ram[32776] = {9'd23,-10'd377};
ram[32777] = {9'd26,-10'd374};
ram[32778] = {9'd29,-10'd371};
ram[32779] = {9'd32,-10'd368};
ram[32780] = {9'd36,-10'd365};
ram[32781] = {9'd39,-10'd362};
ram[32782] = {9'd42,-10'd359};
ram[32783] = {9'd45,-10'd355};
ram[32784] = {9'd48,-10'd352};
ram[32785] = {9'd51,-10'd349};
ram[32786] = {9'd54,-10'd346};
ram[32787] = {9'd58,-10'd343};
ram[32788] = {9'd61,-10'd340};
ram[32789] = {9'd64,-10'd337};
ram[32790] = {9'd67,-10'd334};
ram[32791] = {9'd70,-10'd330};
ram[32792] = {9'd73,-10'd327};
ram[32793] = {9'd76,-10'd324};
ram[32794] = {9'd80,-10'd321};
ram[32795] = {9'd83,-10'd318};
ram[32796] = {9'd86,-10'd315};
ram[32797] = {9'd89,-10'd312};
ram[32798] = {9'd92,-10'd308};
ram[32799] = {9'd95,-10'd305};
ram[32800] = {9'd98,-10'd302};
ram[32801] = {-9'd99,-10'd299};
ram[32802] = {-9'd96,-10'd296};
ram[32803] = {-9'd92,-10'd293};
ram[32804] = {-9'd89,-10'd290};
ram[32805] = {-9'd86,-10'd286};
ram[32806] = {-9'd83,-10'd283};
ram[32807] = {-9'd80,-10'd280};
ram[32808] = {-9'd77,-10'd277};
ram[32809] = {-9'd74,-10'd274};
ram[32810] = {-9'd70,-10'd271};
ram[32811] = {-9'd67,-10'd268};
ram[32812] = {-9'd64,-10'd264};
ram[32813] = {-9'd61,-10'd261};
ram[32814] = {-9'd58,-10'd258};
ram[32815] = {-9'd55,-10'd255};
ram[32816] = {-9'd52,-10'd252};
ram[32817] = {-9'd48,-10'd249};
ram[32818] = {-9'd45,-10'd246};
ram[32819] = {-9'd42,-10'd242};
ram[32820] = {-9'd39,-10'd239};
ram[32821] = {-9'd36,-10'd236};
ram[32822] = {-9'd33,-10'd233};
ram[32823] = {-9'd30,-10'd230};
ram[32824] = {-9'd26,-10'd227};
ram[32825] = {-9'd23,-10'd224};
ram[32826] = {-9'd20,-10'd220};
ram[32827] = {-9'd17,-10'd217};
ram[32828] = {-9'd14,-10'd214};
ram[32829] = {-9'd11,-10'd211};
ram[32830] = {-9'd8,-10'd208};
ram[32831] = {-9'd4,-10'd205};
ram[32832] = {-9'd1,-10'd202};
ram[32833] = {9'd2,-10'd198};
ram[32834] = {9'd5,-10'd195};
ram[32835] = {9'd8,-10'd192};
ram[32836] = {9'd11,-10'd189};
ram[32837] = {9'd14,-10'd186};
ram[32838] = {9'd18,-10'd183};
ram[32839] = {9'd21,-10'd180};
ram[32840] = {9'd24,-10'd176};
ram[32841] = {9'd27,-10'd173};
ram[32842] = {9'd30,-10'd170};
ram[32843] = {9'd33,-10'd167};
ram[32844] = {9'd36,-10'd164};
ram[32845] = {9'd40,-10'd161};
ram[32846] = {9'd43,-10'd158};
ram[32847] = {9'd46,-10'd154};
ram[32848] = {9'd49,-10'd151};
ram[32849] = {9'd52,-10'd148};
ram[32850] = {9'd55,-10'd145};
ram[32851] = {9'd58,-10'd142};
ram[32852] = {9'd62,-10'd139};
ram[32853] = {9'd65,-10'd136};
ram[32854] = {9'd68,-10'd132};
ram[32855] = {9'd71,-10'd129};
ram[32856] = {9'd74,-10'd126};
ram[32857] = {9'd77,-10'd123};
ram[32858] = {9'd80,-10'd120};
ram[32859] = {9'd84,-10'd117};
ram[32860] = {9'd87,-10'd114};
ram[32861] = {9'd90,-10'd110};
ram[32862] = {9'd93,-10'd107};
ram[32863] = {9'd96,-10'd104};
ram[32864] = {9'd99,-10'd101};
ram[32865] = {-9'd98,-10'd98};
ram[32866] = {-9'd95,-10'd95};
ram[32867] = {-9'd92,-10'd92};
ram[32868] = {-9'd88,-10'd88};
ram[32869] = {-9'd85,-10'd85};
ram[32870] = {-9'd82,-10'd82};
ram[32871] = {-9'd79,-10'd79};
ram[32872] = {-9'd76,-10'd76};
ram[32873] = {-9'd73,-10'd73};
ram[32874] = {-9'd70,-10'd70};
ram[32875] = {-9'd66,-10'd66};
ram[32876] = {-9'd63,-10'd63};
ram[32877] = {-9'd60,-10'd60};
ram[32878] = {-9'd57,-10'd57};
ram[32879] = {-9'd54,-10'd54};
ram[32880] = {-9'd51,-10'd51};
ram[32881] = {-9'd48,-10'd48};
ram[32882] = {-9'd44,-10'd44};
ram[32883] = {-9'd41,-10'd41};
ram[32884] = {-9'd38,-10'd38};
ram[32885] = {-9'd35,-10'd35};
ram[32886] = {-9'd32,-10'd32};
ram[32887] = {-9'd29,-10'd29};
ram[32888] = {-9'd26,-10'd26};
ram[32889] = {-9'd22,-10'd22};
ram[32890] = {-9'd19,-10'd19};
ram[32891] = {-9'd16,-10'd16};
ram[32892] = {-9'd13,-10'd13};
ram[32893] = {-9'd10,-10'd10};
ram[32894] = {-9'd7,-10'd7};
ram[32895] = {-9'd4,-10'd4};
ram[32896] = {-9'd4,-10'd4};
ram[32897] = {9'd0,10'd0};
ram[32898] = {9'd3,10'd3};
ram[32899] = {9'd6,10'd6};
ram[32900] = {9'd9,10'd9};
ram[32901] = {9'd12,10'd12};
ram[32902] = {9'd15,10'd15};
ram[32903] = {9'd18,10'd18};
ram[32904] = {9'd21,10'd21};
ram[32905] = {9'd25,10'd25};
ram[32906] = {9'd28,10'd28};
ram[32907] = {9'd31,10'd31};
ram[32908] = {9'd34,10'd34};
ram[32909] = {9'd37,10'd37};
ram[32910] = {9'd40,10'd40};
ram[32911] = {9'd43,10'd43};
ram[32912] = {9'd47,10'd47};
ram[32913] = {9'd50,10'd50};
ram[32914] = {9'd53,10'd53};
ram[32915] = {9'd56,10'd56};
ram[32916] = {9'd59,10'd59};
ram[32917] = {9'd62,10'd62};
ram[32918] = {9'd65,10'd65};
ram[32919] = {9'd69,10'd69};
ram[32920] = {9'd72,10'd72};
ram[32921] = {9'd75,10'd75};
ram[32922] = {9'd78,10'd78};
ram[32923] = {9'd81,10'd81};
ram[32924] = {9'd84,10'd84};
ram[32925] = {9'd87,10'd87};
ram[32926] = {9'd91,10'd91};
ram[32927] = {9'd94,10'd94};
ram[32928] = {9'd97,10'd97};
ram[32929] = {-9'd100,10'd100};
ram[32930] = {-9'd97,10'd103};
ram[32931] = {-9'd94,10'd106};
ram[32932] = {-9'd91,10'd109};
ram[32933] = {-9'd88,10'd113};
ram[32934] = {-9'd85,10'd116};
ram[32935] = {-9'd81,10'd119};
ram[32936] = {-9'd78,10'd122};
ram[32937] = {-9'd75,10'd125};
ram[32938] = {-9'd72,10'd128};
ram[32939] = {-9'd69,10'd131};
ram[32940] = {-9'd66,10'd135};
ram[32941] = {-9'd63,10'd138};
ram[32942] = {-9'd59,10'd141};
ram[32943] = {-9'd56,10'd144};
ram[32944] = {-9'd53,10'd147};
ram[32945] = {-9'd50,10'd150};
ram[32946] = {-9'd47,10'd153};
ram[32947] = {-9'd44,10'd157};
ram[32948] = {-9'd41,10'd160};
ram[32949] = {-9'd37,10'd163};
ram[32950] = {-9'd34,10'd166};
ram[32951] = {-9'd31,10'd169};
ram[32952] = {-9'd28,10'd172};
ram[32953] = {-9'd25,10'd175};
ram[32954] = {-9'd22,10'd179};
ram[32955] = {-9'd19,10'd182};
ram[32956] = {-9'd15,10'd185};
ram[32957] = {-9'd12,10'd188};
ram[32958] = {-9'd9,10'd191};
ram[32959] = {-9'd6,10'd194};
ram[32960] = {-9'd3,10'd197};
ram[32961] = {9'd0,10'd201};
ram[32962] = {9'd3,10'd204};
ram[32963] = {9'd7,10'd207};
ram[32964] = {9'd10,10'd210};
ram[32965] = {9'd13,10'd213};
ram[32966] = {9'd16,10'd216};
ram[32967] = {9'd19,10'd219};
ram[32968] = {9'd22,10'd223};
ram[32969] = {9'd25,10'd226};
ram[32970] = {9'd29,10'd229};
ram[32971] = {9'd32,10'd232};
ram[32972] = {9'd35,10'd235};
ram[32973] = {9'd38,10'd238};
ram[32974] = {9'd41,10'd241};
ram[32975] = {9'd44,10'd245};
ram[32976] = {9'd47,10'd248};
ram[32977] = {9'd51,10'd251};
ram[32978] = {9'd54,10'd254};
ram[32979] = {9'd57,10'd257};
ram[32980] = {9'd60,10'd260};
ram[32981] = {9'd63,10'd263};
ram[32982] = {9'd66,10'd267};
ram[32983] = {9'd69,10'd270};
ram[32984] = {9'd73,10'd273};
ram[32985] = {9'd76,10'd276};
ram[32986] = {9'd79,10'd279};
ram[32987] = {9'd82,10'd282};
ram[32988] = {9'd85,10'd285};
ram[32989] = {9'd88,10'd289};
ram[32990] = {9'd91,10'd292};
ram[32991] = {9'd95,10'd295};
ram[32992] = {9'd98,10'd298};
ram[32993] = {-9'd99,10'd301};
ram[32994] = {-9'd96,10'd304};
ram[32995] = {-9'd93,10'd307};
ram[32996] = {-9'd90,10'd311};
ram[32997] = {-9'd87,10'd314};
ram[32998] = {-9'd84,10'd317};
ram[32999] = {-9'd81,10'd320};
ram[33000] = {-9'd77,10'd323};
ram[33001] = {-9'd74,10'd326};
ram[33002] = {-9'd71,10'd329};
ram[33003] = {-9'd68,10'd333};
ram[33004] = {-9'd65,10'd336};
ram[33005] = {-9'd62,10'd339};
ram[33006] = {-9'd59,10'd342};
ram[33007] = {-9'd55,10'd345};
ram[33008] = {-9'd52,10'd348};
ram[33009] = {-9'd49,10'd351};
ram[33010] = {-9'd46,10'd354};
ram[33011] = {-9'd43,10'd358};
ram[33012] = {-9'd40,10'd361};
ram[33013] = {-9'd37,10'd364};
ram[33014] = {-9'd33,10'd367};
ram[33015] = {-9'd30,10'd370};
ram[33016] = {-9'd27,10'd373};
ram[33017] = {-9'd24,10'd376};
ram[33018] = {-9'd21,10'd380};
ram[33019] = {-9'd18,10'd383};
ram[33020] = {-9'd15,10'd386};
ram[33021] = {-9'd11,10'd389};
ram[33022] = {-9'd8,10'd392};
ram[33023] = {-9'd5,10'd395};
ram[33024] = {-9'd5,10'd395};
ram[33025] = {-9'd2,10'd398};
ram[33026] = {9'd1,-10'd399};
ram[33027] = {9'd4,-10'd396};
ram[33028] = {9'd7,-10'd393};
ram[33029] = {9'd10,-10'd390};
ram[33030] = {9'd14,-10'd387};
ram[33031] = {9'd17,-10'd384};
ram[33032] = {9'd20,-10'd381};
ram[33033] = {9'd23,-10'd377};
ram[33034] = {9'd26,-10'd374};
ram[33035] = {9'd29,-10'd371};
ram[33036] = {9'd32,-10'd368};
ram[33037] = {9'd36,-10'd365};
ram[33038] = {9'd39,-10'd362};
ram[33039] = {9'd42,-10'd359};
ram[33040] = {9'd45,-10'd355};
ram[33041] = {9'd48,-10'd352};
ram[33042] = {9'd51,-10'd349};
ram[33043] = {9'd54,-10'd346};
ram[33044] = {9'd58,-10'd343};
ram[33045] = {9'd61,-10'd340};
ram[33046] = {9'd64,-10'd337};
ram[33047] = {9'd67,-10'd334};
ram[33048] = {9'd70,-10'd330};
ram[33049] = {9'd73,-10'd327};
ram[33050] = {9'd76,-10'd324};
ram[33051] = {9'd80,-10'd321};
ram[33052] = {9'd83,-10'd318};
ram[33053] = {9'd86,-10'd315};
ram[33054] = {9'd89,-10'd312};
ram[33055] = {9'd92,-10'd308};
ram[33056] = {9'd95,-10'd305};
ram[33057] = {9'd98,-10'd302};
ram[33058] = {-9'd99,-10'd299};
ram[33059] = {-9'd96,-10'd296};
ram[33060] = {-9'd92,-10'd293};
ram[33061] = {-9'd89,-10'd290};
ram[33062] = {-9'd86,-10'd286};
ram[33063] = {-9'd83,-10'd283};
ram[33064] = {-9'd80,-10'd280};
ram[33065] = {-9'd77,-10'd277};
ram[33066] = {-9'd74,-10'd274};
ram[33067] = {-9'd70,-10'd271};
ram[33068] = {-9'd67,-10'd268};
ram[33069] = {-9'd64,-10'd264};
ram[33070] = {-9'd61,-10'd261};
ram[33071] = {-9'd58,-10'd258};
ram[33072] = {-9'd55,-10'd255};
ram[33073] = {-9'd52,-10'd252};
ram[33074] = {-9'd48,-10'd249};
ram[33075] = {-9'd45,-10'd246};
ram[33076] = {-9'd42,-10'd242};
ram[33077] = {-9'd39,-10'd239};
ram[33078] = {-9'd36,-10'd236};
ram[33079] = {-9'd33,-10'd233};
ram[33080] = {-9'd30,-10'd230};
ram[33081] = {-9'd26,-10'd227};
ram[33082] = {-9'd23,-10'd224};
ram[33083] = {-9'd20,-10'd220};
ram[33084] = {-9'd17,-10'd217};
ram[33085] = {-9'd14,-10'd214};
ram[33086] = {-9'd11,-10'd211};
ram[33087] = {-9'd8,-10'd208};
ram[33088] = {-9'd4,-10'd205};
ram[33089] = {-9'd1,-10'd202};
ram[33090] = {9'd2,-10'd198};
ram[33091] = {9'd5,-10'd195};
ram[33092] = {9'd8,-10'd192};
ram[33093] = {9'd11,-10'd189};
ram[33094] = {9'd14,-10'd186};
ram[33095] = {9'd18,-10'd183};
ram[33096] = {9'd21,-10'd180};
ram[33097] = {9'd24,-10'd176};
ram[33098] = {9'd27,-10'd173};
ram[33099] = {9'd30,-10'd170};
ram[33100] = {9'd33,-10'd167};
ram[33101] = {9'd36,-10'd164};
ram[33102] = {9'd40,-10'd161};
ram[33103] = {9'd43,-10'd158};
ram[33104] = {9'd46,-10'd154};
ram[33105] = {9'd49,-10'd151};
ram[33106] = {9'd52,-10'd148};
ram[33107] = {9'd55,-10'd145};
ram[33108] = {9'd58,-10'd142};
ram[33109] = {9'd62,-10'd139};
ram[33110] = {9'd65,-10'd136};
ram[33111] = {9'd68,-10'd132};
ram[33112] = {9'd71,-10'd129};
ram[33113] = {9'd74,-10'd126};
ram[33114] = {9'd77,-10'd123};
ram[33115] = {9'd80,-10'd120};
ram[33116] = {9'd84,-10'd117};
ram[33117] = {9'd87,-10'd114};
ram[33118] = {9'd90,-10'd110};
ram[33119] = {9'd93,-10'd107};
ram[33120] = {9'd96,-10'd104};
ram[33121] = {9'd99,-10'd101};
ram[33122] = {-9'd98,-10'd98};
ram[33123] = {-9'd95,-10'd95};
ram[33124] = {-9'd92,-10'd92};
ram[33125] = {-9'd88,-10'd88};
ram[33126] = {-9'd85,-10'd85};
ram[33127] = {-9'd82,-10'd82};
ram[33128] = {-9'd79,-10'd79};
ram[33129] = {-9'd76,-10'd76};
ram[33130] = {-9'd73,-10'd73};
ram[33131] = {-9'd70,-10'd70};
ram[33132] = {-9'd66,-10'd66};
ram[33133] = {-9'd63,-10'd63};
ram[33134] = {-9'd60,-10'd60};
ram[33135] = {-9'd57,-10'd57};
ram[33136] = {-9'd54,-10'd54};
ram[33137] = {-9'd51,-10'd51};
ram[33138] = {-9'd48,-10'd48};
ram[33139] = {-9'd44,-10'd44};
ram[33140] = {-9'd41,-10'd41};
ram[33141] = {-9'd38,-10'd38};
ram[33142] = {-9'd35,-10'd35};
ram[33143] = {-9'd32,-10'd32};
ram[33144] = {-9'd29,-10'd29};
ram[33145] = {-9'd26,-10'd26};
ram[33146] = {-9'd22,-10'd22};
ram[33147] = {-9'd19,-10'd19};
ram[33148] = {-9'd16,-10'd16};
ram[33149] = {-9'd13,-10'd13};
ram[33150] = {-9'd10,-10'd10};
ram[33151] = {-9'd7,-10'd7};
ram[33152] = {-9'd7,-10'd7};
ram[33153] = {-9'd4,-10'd4};
ram[33154] = {9'd0,10'd0};
ram[33155] = {9'd3,10'd3};
ram[33156] = {9'd6,10'd6};
ram[33157] = {9'd9,10'd9};
ram[33158] = {9'd12,10'd12};
ram[33159] = {9'd15,10'd15};
ram[33160] = {9'd18,10'd18};
ram[33161] = {9'd21,10'd21};
ram[33162] = {9'd25,10'd25};
ram[33163] = {9'd28,10'd28};
ram[33164] = {9'd31,10'd31};
ram[33165] = {9'd34,10'd34};
ram[33166] = {9'd37,10'd37};
ram[33167] = {9'd40,10'd40};
ram[33168] = {9'd43,10'd43};
ram[33169] = {9'd47,10'd47};
ram[33170] = {9'd50,10'd50};
ram[33171] = {9'd53,10'd53};
ram[33172] = {9'd56,10'd56};
ram[33173] = {9'd59,10'd59};
ram[33174] = {9'd62,10'd62};
ram[33175] = {9'd65,10'd65};
ram[33176] = {9'd69,10'd69};
ram[33177] = {9'd72,10'd72};
ram[33178] = {9'd75,10'd75};
ram[33179] = {9'd78,10'd78};
ram[33180] = {9'd81,10'd81};
ram[33181] = {9'd84,10'd84};
ram[33182] = {9'd87,10'd87};
ram[33183] = {9'd91,10'd91};
ram[33184] = {9'd94,10'd94};
ram[33185] = {9'd97,10'd97};
ram[33186] = {-9'd100,10'd100};
ram[33187] = {-9'd97,10'd103};
ram[33188] = {-9'd94,10'd106};
ram[33189] = {-9'd91,10'd109};
ram[33190] = {-9'd88,10'd113};
ram[33191] = {-9'd85,10'd116};
ram[33192] = {-9'd81,10'd119};
ram[33193] = {-9'd78,10'd122};
ram[33194] = {-9'd75,10'd125};
ram[33195] = {-9'd72,10'd128};
ram[33196] = {-9'd69,10'd131};
ram[33197] = {-9'd66,10'd135};
ram[33198] = {-9'd63,10'd138};
ram[33199] = {-9'd59,10'd141};
ram[33200] = {-9'd56,10'd144};
ram[33201] = {-9'd53,10'd147};
ram[33202] = {-9'd50,10'd150};
ram[33203] = {-9'd47,10'd153};
ram[33204] = {-9'd44,10'd157};
ram[33205] = {-9'd41,10'd160};
ram[33206] = {-9'd37,10'd163};
ram[33207] = {-9'd34,10'd166};
ram[33208] = {-9'd31,10'd169};
ram[33209] = {-9'd28,10'd172};
ram[33210] = {-9'd25,10'd175};
ram[33211] = {-9'd22,10'd179};
ram[33212] = {-9'd19,10'd182};
ram[33213] = {-9'd15,10'd185};
ram[33214] = {-9'd12,10'd188};
ram[33215] = {-9'd9,10'd191};
ram[33216] = {-9'd6,10'd194};
ram[33217] = {-9'd3,10'd197};
ram[33218] = {9'd0,10'd201};
ram[33219] = {9'd3,10'd204};
ram[33220] = {9'd7,10'd207};
ram[33221] = {9'd10,10'd210};
ram[33222] = {9'd13,10'd213};
ram[33223] = {9'd16,10'd216};
ram[33224] = {9'd19,10'd219};
ram[33225] = {9'd22,10'd223};
ram[33226] = {9'd25,10'd226};
ram[33227] = {9'd29,10'd229};
ram[33228] = {9'd32,10'd232};
ram[33229] = {9'd35,10'd235};
ram[33230] = {9'd38,10'd238};
ram[33231] = {9'd41,10'd241};
ram[33232] = {9'd44,10'd245};
ram[33233] = {9'd47,10'd248};
ram[33234] = {9'd51,10'd251};
ram[33235] = {9'd54,10'd254};
ram[33236] = {9'd57,10'd257};
ram[33237] = {9'd60,10'd260};
ram[33238] = {9'd63,10'd263};
ram[33239] = {9'd66,10'd267};
ram[33240] = {9'd69,10'd270};
ram[33241] = {9'd73,10'd273};
ram[33242] = {9'd76,10'd276};
ram[33243] = {9'd79,10'd279};
ram[33244] = {9'd82,10'd282};
ram[33245] = {9'd85,10'd285};
ram[33246] = {9'd88,10'd289};
ram[33247] = {9'd91,10'd292};
ram[33248] = {9'd95,10'd295};
ram[33249] = {9'd98,10'd298};
ram[33250] = {-9'd99,10'd301};
ram[33251] = {-9'd96,10'd304};
ram[33252] = {-9'd93,10'd307};
ram[33253] = {-9'd90,10'd311};
ram[33254] = {-9'd87,10'd314};
ram[33255] = {-9'd84,10'd317};
ram[33256] = {-9'd81,10'd320};
ram[33257] = {-9'd77,10'd323};
ram[33258] = {-9'd74,10'd326};
ram[33259] = {-9'd71,10'd329};
ram[33260] = {-9'd68,10'd333};
ram[33261] = {-9'd65,10'd336};
ram[33262] = {-9'd62,10'd339};
ram[33263] = {-9'd59,10'd342};
ram[33264] = {-9'd55,10'd345};
ram[33265] = {-9'd52,10'd348};
ram[33266] = {-9'd49,10'd351};
ram[33267] = {-9'd46,10'd354};
ram[33268] = {-9'd43,10'd358};
ram[33269] = {-9'd40,10'd361};
ram[33270] = {-9'd37,10'd364};
ram[33271] = {-9'd33,10'd367};
ram[33272] = {-9'd30,10'd370};
ram[33273] = {-9'd27,10'd373};
ram[33274] = {-9'd24,10'd376};
ram[33275] = {-9'd21,10'd380};
ram[33276] = {-9'd18,10'd383};
ram[33277] = {-9'd15,10'd386};
ram[33278] = {-9'd11,10'd389};
ram[33279] = {-9'd8,10'd392};
ram[33280] = {-9'd8,10'd392};
ram[33281] = {-9'd5,10'd395};
ram[33282] = {-9'd2,10'd398};
ram[33283] = {9'd1,-10'd399};
ram[33284] = {9'd4,-10'd396};
ram[33285] = {9'd7,-10'd393};
ram[33286] = {9'd10,-10'd390};
ram[33287] = {9'd14,-10'd387};
ram[33288] = {9'd17,-10'd384};
ram[33289] = {9'd20,-10'd381};
ram[33290] = {9'd23,-10'd377};
ram[33291] = {9'd26,-10'd374};
ram[33292] = {9'd29,-10'd371};
ram[33293] = {9'd32,-10'd368};
ram[33294] = {9'd36,-10'd365};
ram[33295] = {9'd39,-10'd362};
ram[33296] = {9'd42,-10'd359};
ram[33297] = {9'd45,-10'd355};
ram[33298] = {9'd48,-10'd352};
ram[33299] = {9'd51,-10'd349};
ram[33300] = {9'd54,-10'd346};
ram[33301] = {9'd58,-10'd343};
ram[33302] = {9'd61,-10'd340};
ram[33303] = {9'd64,-10'd337};
ram[33304] = {9'd67,-10'd334};
ram[33305] = {9'd70,-10'd330};
ram[33306] = {9'd73,-10'd327};
ram[33307] = {9'd76,-10'd324};
ram[33308] = {9'd80,-10'd321};
ram[33309] = {9'd83,-10'd318};
ram[33310] = {9'd86,-10'd315};
ram[33311] = {9'd89,-10'd312};
ram[33312] = {9'd92,-10'd308};
ram[33313] = {9'd95,-10'd305};
ram[33314] = {9'd98,-10'd302};
ram[33315] = {-9'd99,-10'd299};
ram[33316] = {-9'd96,-10'd296};
ram[33317] = {-9'd92,-10'd293};
ram[33318] = {-9'd89,-10'd290};
ram[33319] = {-9'd86,-10'd286};
ram[33320] = {-9'd83,-10'd283};
ram[33321] = {-9'd80,-10'd280};
ram[33322] = {-9'd77,-10'd277};
ram[33323] = {-9'd74,-10'd274};
ram[33324] = {-9'd70,-10'd271};
ram[33325] = {-9'd67,-10'd268};
ram[33326] = {-9'd64,-10'd264};
ram[33327] = {-9'd61,-10'd261};
ram[33328] = {-9'd58,-10'd258};
ram[33329] = {-9'd55,-10'd255};
ram[33330] = {-9'd52,-10'd252};
ram[33331] = {-9'd48,-10'd249};
ram[33332] = {-9'd45,-10'd246};
ram[33333] = {-9'd42,-10'd242};
ram[33334] = {-9'd39,-10'd239};
ram[33335] = {-9'd36,-10'd236};
ram[33336] = {-9'd33,-10'd233};
ram[33337] = {-9'd30,-10'd230};
ram[33338] = {-9'd26,-10'd227};
ram[33339] = {-9'd23,-10'd224};
ram[33340] = {-9'd20,-10'd220};
ram[33341] = {-9'd17,-10'd217};
ram[33342] = {-9'd14,-10'd214};
ram[33343] = {-9'd11,-10'd211};
ram[33344] = {-9'd8,-10'd208};
ram[33345] = {-9'd4,-10'd205};
ram[33346] = {-9'd1,-10'd202};
ram[33347] = {9'd2,-10'd198};
ram[33348] = {9'd5,-10'd195};
ram[33349] = {9'd8,-10'd192};
ram[33350] = {9'd11,-10'd189};
ram[33351] = {9'd14,-10'd186};
ram[33352] = {9'd18,-10'd183};
ram[33353] = {9'd21,-10'd180};
ram[33354] = {9'd24,-10'd176};
ram[33355] = {9'd27,-10'd173};
ram[33356] = {9'd30,-10'd170};
ram[33357] = {9'd33,-10'd167};
ram[33358] = {9'd36,-10'd164};
ram[33359] = {9'd40,-10'd161};
ram[33360] = {9'd43,-10'd158};
ram[33361] = {9'd46,-10'd154};
ram[33362] = {9'd49,-10'd151};
ram[33363] = {9'd52,-10'd148};
ram[33364] = {9'd55,-10'd145};
ram[33365] = {9'd58,-10'd142};
ram[33366] = {9'd62,-10'd139};
ram[33367] = {9'd65,-10'd136};
ram[33368] = {9'd68,-10'd132};
ram[33369] = {9'd71,-10'd129};
ram[33370] = {9'd74,-10'd126};
ram[33371] = {9'd77,-10'd123};
ram[33372] = {9'd80,-10'd120};
ram[33373] = {9'd84,-10'd117};
ram[33374] = {9'd87,-10'd114};
ram[33375] = {9'd90,-10'd110};
ram[33376] = {9'd93,-10'd107};
ram[33377] = {9'd96,-10'd104};
ram[33378] = {9'd99,-10'd101};
ram[33379] = {-9'd98,-10'd98};
ram[33380] = {-9'd95,-10'd95};
ram[33381] = {-9'd92,-10'd92};
ram[33382] = {-9'd88,-10'd88};
ram[33383] = {-9'd85,-10'd85};
ram[33384] = {-9'd82,-10'd82};
ram[33385] = {-9'd79,-10'd79};
ram[33386] = {-9'd76,-10'd76};
ram[33387] = {-9'd73,-10'd73};
ram[33388] = {-9'd70,-10'd70};
ram[33389] = {-9'd66,-10'd66};
ram[33390] = {-9'd63,-10'd63};
ram[33391] = {-9'd60,-10'd60};
ram[33392] = {-9'd57,-10'd57};
ram[33393] = {-9'd54,-10'd54};
ram[33394] = {-9'd51,-10'd51};
ram[33395] = {-9'd48,-10'd48};
ram[33396] = {-9'd44,-10'd44};
ram[33397] = {-9'd41,-10'd41};
ram[33398] = {-9'd38,-10'd38};
ram[33399] = {-9'd35,-10'd35};
ram[33400] = {-9'd32,-10'd32};
ram[33401] = {-9'd29,-10'd29};
ram[33402] = {-9'd26,-10'd26};
ram[33403] = {-9'd22,-10'd22};
ram[33404] = {-9'd19,-10'd19};
ram[33405] = {-9'd16,-10'd16};
ram[33406] = {-9'd13,-10'd13};
ram[33407] = {-9'd10,-10'd10};
ram[33408] = {-9'd10,-10'd10};
ram[33409] = {-9'd7,-10'd7};
ram[33410] = {-9'd4,-10'd4};
ram[33411] = {9'd0,10'd0};
ram[33412] = {9'd3,10'd3};
ram[33413] = {9'd6,10'd6};
ram[33414] = {9'd9,10'd9};
ram[33415] = {9'd12,10'd12};
ram[33416] = {9'd15,10'd15};
ram[33417] = {9'd18,10'd18};
ram[33418] = {9'd21,10'd21};
ram[33419] = {9'd25,10'd25};
ram[33420] = {9'd28,10'd28};
ram[33421] = {9'd31,10'd31};
ram[33422] = {9'd34,10'd34};
ram[33423] = {9'd37,10'd37};
ram[33424] = {9'd40,10'd40};
ram[33425] = {9'd43,10'd43};
ram[33426] = {9'd47,10'd47};
ram[33427] = {9'd50,10'd50};
ram[33428] = {9'd53,10'd53};
ram[33429] = {9'd56,10'd56};
ram[33430] = {9'd59,10'd59};
ram[33431] = {9'd62,10'd62};
ram[33432] = {9'd65,10'd65};
ram[33433] = {9'd69,10'd69};
ram[33434] = {9'd72,10'd72};
ram[33435] = {9'd75,10'd75};
ram[33436] = {9'd78,10'd78};
ram[33437] = {9'd81,10'd81};
ram[33438] = {9'd84,10'd84};
ram[33439] = {9'd87,10'd87};
ram[33440] = {9'd91,10'd91};
ram[33441] = {9'd94,10'd94};
ram[33442] = {9'd97,10'd97};
ram[33443] = {-9'd100,10'd100};
ram[33444] = {-9'd97,10'd103};
ram[33445] = {-9'd94,10'd106};
ram[33446] = {-9'd91,10'd109};
ram[33447] = {-9'd88,10'd113};
ram[33448] = {-9'd85,10'd116};
ram[33449] = {-9'd81,10'd119};
ram[33450] = {-9'd78,10'd122};
ram[33451] = {-9'd75,10'd125};
ram[33452] = {-9'd72,10'd128};
ram[33453] = {-9'd69,10'd131};
ram[33454] = {-9'd66,10'd135};
ram[33455] = {-9'd63,10'd138};
ram[33456] = {-9'd59,10'd141};
ram[33457] = {-9'd56,10'd144};
ram[33458] = {-9'd53,10'd147};
ram[33459] = {-9'd50,10'd150};
ram[33460] = {-9'd47,10'd153};
ram[33461] = {-9'd44,10'd157};
ram[33462] = {-9'd41,10'd160};
ram[33463] = {-9'd37,10'd163};
ram[33464] = {-9'd34,10'd166};
ram[33465] = {-9'd31,10'd169};
ram[33466] = {-9'd28,10'd172};
ram[33467] = {-9'd25,10'd175};
ram[33468] = {-9'd22,10'd179};
ram[33469] = {-9'd19,10'd182};
ram[33470] = {-9'd15,10'd185};
ram[33471] = {-9'd12,10'd188};
ram[33472] = {-9'd9,10'd191};
ram[33473] = {-9'd6,10'd194};
ram[33474] = {-9'd3,10'd197};
ram[33475] = {9'd0,10'd201};
ram[33476] = {9'd3,10'd204};
ram[33477] = {9'd7,10'd207};
ram[33478] = {9'd10,10'd210};
ram[33479] = {9'd13,10'd213};
ram[33480] = {9'd16,10'd216};
ram[33481] = {9'd19,10'd219};
ram[33482] = {9'd22,10'd223};
ram[33483] = {9'd25,10'd226};
ram[33484] = {9'd29,10'd229};
ram[33485] = {9'd32,10'd232};
ram[33486] = {9'd35,10'd235};
ram[33487] = {9'd38,10'd238};
ram[33488] = {9'd41,10'd241};
ram[33489] = {9'd44,10'd245};
ram[33490] = {9'd47,10'd248};
ram[33491] = {9'd51,10'd251};
ram[33492] = {9'd54,10'd254};
ram[33493] = {9'd57,10'd257};
ram[33494] = {9'd60,10'd260};
ram[33495] = {9'd63,10'd263};
ram[33496] = {9'd66,10'd267};
ram[33497] = {9'd69,10'd270};
ram[33498] = {9'd73,10'd273};
ram[33499] = {9'd76,10'd276};
ram[33500] = {9'd79,10'd279};
ram[33501] = {9'd82,10'd282};
ram[33502] = {9'd85,10'd285};
ram[33503] = {9'd88,10'd289};
ram[33504] = {9'd91,10'd292};
ram[33505] = {9'd95,10'd295};
ram[33506] = {9'd98,10'd298};
ram[33507] = {-9'd99,10'd301};
ram[33508] = {-9'd96,10'd304};
ram[33509] = {-9'd93,10'd307};
ram[33510] = {-9'd90,10'd311};
ram[33511] = {-9'd87,10'd314};
ram[33512] = {-9'd84,10'd317};
ram[33513] = {-9'd81,10'd320};
ram[33514] = {-9'd77,10'd323};
ram[33515] = {-9'd74,10'd326};
ram[33516] = {-9'd71,10'd329};
ram[33517] = {-9'd68,10'd333};
ram[33518] = {-9'd65,10'd336};
ram[33519] = {-9'd62,10'd339};
ram[33520] = {-9'd59,10'd342};
ram[33521] = {-9'd55,10'd345};
ram[33522] = {-9'd52,10'd348};
ram[33523] = {-9'd49,10'd351};
ram[33524] = {-9'd46,10'd354};
ram[33525] = {-9'd43,10'd358};
ram[33526] = {-9'd40,10'd361};
ram[33527] = {-9'd37,10'd364};
ram[33528] = {-9'd33,10'd367};
ram[33529] = {-9'd30,10'd370};
ram[33530] = {-9'd27,10'd373};
ram[33531] = {-9'd24,10'd376};
ram[33532] = {-9'd21,10'd380};
ram[33533] = {-9'd18,10'd383};
ram[33534] = {-9'd15,10'd386};
ram[33535] = {-9'd11,10'd389};
ram[33536] = {-9'd11,10'd389};
ram[33537] = {-9'd8,10'd392};
ram[33538] = {-9'd5,10'd395};
ram[33539] = {-9'd2,10'd398};
ram[33540] = {9'd1,-10'd399};
ram[33541] = {9'd4,-10'd396};
ram[33542] = {9'd7,-10'd393};
ram[33543] = {9'd10,-10'd390};
ram[33544] = {9'd14,-10'd387};
ram[33545] = {9'd17,-10'd384};
ram[33546] = {9'd20,-10'd381};
ram[33547] = {9'd23,-10'd377};
ram[33548] = {9'd26,-10'd374};
ram[33549] = {9'd29,-10'd371};
ram[33550] = {9'd32,-10'd368};
ram[33551] = {9'd36,-10'd365};
ram[33552] = {9'd39,-10'd362};
ram[33553] = {9'd42,-10'd359};
ram[33554] = {9'd45,-10'd355};
ram[33555] = {9'd48,-10'd352};
ram[33556] = {9'd51,-10'd349};
ram[33557] = {9'd54,-10'd346};
ram[33558] = {9'd58,-10'd343};
ram[33559] = {9'd61,-10'd340};
ram[33560] = {9'd64,-10'd337};
ram[33561] = {9'd67,-10'd334};
ram[33562] = {9'd70,-10'd330};
ram[33563] = {9'd73,-10'd327};
ram[33564] = {9'd76,-10'd324};
ram[33565] = {9'd80,-10'd321};
ram[33566] = {9'd83,-10'd318};
ram[33567] = {9'd86,-10'd315};
ram[33568] = {9'd89,-10'd312};
ram[33569] = {9'd92,-10'd308};
ram[33570] = {9'd95,-10'd305};
ram[33571] = {9'd98,-10'd302};
ram[33572] = {-9'd99,-10'd299};
ram[33573] = {-9'd96,-10'd296};
ram[33574] = {-9'd92,-10'd293};
ram[33575] = {-9'd89,-10'd290};
ram[33576] = {-9'd86,-10'd286};
ram[33577] = {-9'd83,-10'd283};
ram[33578] = {-9'd80,-10'd280};
ram[33579] = {-9'd77,-10'd277};
ram[33580] = {-9'd74,-10'd274};
ram[33581] = {-9'd70,-10'd271};
ram[33582] = {-9'd67,-10'd268};
ram[33583] = {-9'd64,-10'd264};
ram[33584] = {-9'd61,-10'd261};
ram[33585] = {-9'd58,-10'd258};
ram[33586] = {-9'd55,-10'd255};
ram[33587] = {-9'd52,-10'd252};
ram[33588] = {-9'd48,-10'd249};
ram[33589] = {-9'd45,-10'd246};
ram[33590] = {-9'd42,-10'd242};
ram[33591] = {-9'd39,-10'd239};
ram[33592] = {-9'd36,-10'd236};
ram[33593] = {-9'd33,-10'd233};
ram[33594] = {-9'd30,-10'd230};
ram[33595] = {-9'd26,-10'd227};
ram[33596] = {-9'd23,-10'd224};
ram[33597] = {-9'd20,-10'd220};
ram[33598] = {-9'd17,-10'd217};
ram[33599] = {-9'd14,-10'd214};
ram[33600] = {-9'd11,-10'd211};
ram[33601] = {-9'd8,-10'd208};
ram[33602] = {-9'd4,-10'd205};
ram[33603] = {-9'd1,-10'd202};
ram[33604] = {9'd2,-10'd198};
ram[33605] = {9'd5,-10'd195};
ram[33606] = {9'd8,-10'd192};
ram[33607] = {9'd11,-10'd189};
ram[33608] = {9'd14,-10'd186};
ram[33609] = {9'd18,-10'd183};
ram[33610] = {9'd21,-10'd180};
ram[33611] = {9'd24,-10'd176};
ram[33612] = {9'd27,-10'd173};
ram[33613] = {9'd30,-10'd170};
ram[33614] = {9'd33,-10'd167};
ram[33615] = {9'd36,-10'd164};
ram[33616] = {9'd40,-10'd161};
ram[33617] = {9'd43,-10'd158};
ram[33618] = {9'd46,-10'd154};
ram[33619] = {9'd49,-10'd151};
ram[33620] = {9'd52,-10'd148};
ram[33621] = {9'd55,-10'd145};
ram[33622] = {9'd58,-10'd142};
ram[33623] = {9'd62,-10'd139};
ram[33624] = {9'd65,-10'd136};
ram[33625] = {9'd68,-10'd132};
ram[33626] = {9'd71,-10'd129};
ram[33627] = {9'd74,-10'd126};
ram[33628] = {9'd77,-10'd123};
ram[33629] = {9'd80,-10'd120};
ram[33630] = {9'd84,-10'd117};
ram[33631] = {9'd87,-10'd114};
ram[33632] = {9'd90,-10'd110};
ram[33633] = {9'd93,-10'd107};
ram[33634] = {9'd96,-10'd104};
ram[33635] = {9'd99,-10'd101};
ram[33636] = {-9'd98,-10'd98};
ram[33637] = {-9'd95,-10'd95};
ram[33638] = {-9'd92,-10'd92};
ram[33639] = {-9'd88,-10'd88};
ram[33640] = {-9'd85,-10'd85};
ram[33641] = {-9'd82,-10'd82};
ram[33642] = {-9'd79,-10'd79};
ram[33643] = {-9'd76,-10'd76};
ram[33644] = {-9'd73,-10'd73};
ram[33645] = {-9'd70,-10'd70};
ram[33646] = {-9'd66,-10'd66};
ram[33647] = {-9'd63,-10'd63};
ram[33648] = {-9'd60,-10'd60};
ram[33649] = {-9'd57,-10'd57};
ram[33650] = {-9'd54,-10'd54};
ram[33651] = {-9'd51,-10'd51};
ram[33652] = {-9'd48,-10'd48};
ram[33653] = {-9'd44,-10'd44};
ram[33654] = {-9'd41,-10'd41};
ram[33655] = {-9'd38,-10'd38};
ram[33656] = {-9'd35,-10'd35};
ram[33657] = {-9'd32,-10'd32};
ram[33658] = {-9'd29,-10'd29};
ram[33659] = {-9'd26,-10'd26};
ram[33660] = {-9'd22,-10'd22};
ram[33661] = {-9'd19,-10'd19};
ram[33662] = {-9'd16,-10'd16};
ram[33663] = {-9'd13,-10'd13};
ram[33664] = {-9'd13,-10'd13};
ram[33665] = {-9'd10,-10'd10};
ram[33666] = {-9'd7,-10'd7};
ram[33667] = {-9'd4,-10'd4};
ram[33668] = {9'd0,10'd0};
ram[33669] = {9'd3,10'd3};
ram[33670] = {9'd6,10'd6};
ram[33671] = {9'd9,10'd9};
ram[33672] = {9'd12,10'd12};
ram[33673] = {9'd15,10'd15};
ram[33674] = {9'd18,10'd18};
ram[33675] = {9'd21,10'd21};
ram[33676] = {9'd25,10'd25};
ram[33677] = {9'd28,10'd28};
ram[33678] = {9'd31,10'd31};
ram[33679] = {9'd34,10'd34};
ram[33680] = {9'd37,10'd37};
ram[33681] = {9'd40,10'd40};
ram[33682] = {9'd43,10'd43};
ram[33683] = {9'd47,10'd47};
ram[33684] = {9'd50,10'd50};
ram[33685] = {9'd53,10'd53};
ram[33686] = {9'd56,10'd56};
ram[33687] = {9'd59,10'd59};
ram[33688] = {9'd62,10'd62};
ram[33689] = {9'd65,10'd65};
ram[33690] = {9'd69,10'd69};
ram[33691] = {9'd72,10'd72};
ram[33692] = {9'd75,10'd75};
ram[33693] = {9'd78,10'd78};
ram[33694] = {9'd81,10'd81};
ram[33695] = {9'd84,10'd84};
ram[33696] = {9'd87,10'd87};
ram[33697] = {9'd91,10'd91};
ram[33698] = {9'd94,10'd94};
ram[33699] = {9'd97,10'd97};
ram[33700] = {-9'd100,10'd100};
ram[33701] = {-9'd97,10'd103};
ram[33702] = {-9'd94,10'd106};
ram[33703] = {-9'd91,10'd109};
ram[33704] = {-9'd88,10'd113};
ram[33705] = {-9'd85,10'd116};
ram[33706] = {-9'd81,10'd119};
ram[33707] = {-9'd78,10'd122};
ram[33708] = {-9'd75,10'd125};
ram[33709] = {-9'd72,10'd128};
ram[33710] = {-9'd69,10'd131};
ram[33711] = {-9'd66,10'd135};
ram[33712] = {-9'd63,10'd138};
ram[33713] = {-9'd59,10'd141};
ram[33714] = {-9'd56,10'd144};
ram[33715] = {-9'd53,10'd147};
ram[33716] = {-9'd50,10'd150};
ram[33717] = {-9'd47,10'd153};
ram[33718] = {-9'd44,10'd157};
ram[33719] = {-9'd41,10'd160};
ram[33720] = {-9'd37,10'd163};
ram[33721] = {-9'd34,10'd166};
ram[33722] = {-9'd31,10'd169};
ram[33723] = {-9'd28,10'd172};
ram[33724] = {-9'd25,10'd175};
ram[33725] = {-9'd22,10'd179};
ram[33726] = {-9'd19,10'd182};
ram[33727] = {-9'd15,10'd185};
ram[33728] = {-9'd12,10'd188};
ram[33729] = {-9'd9,10'd191};
ram[33730] = {-9'd6,10'd194};
ram[33731] = {-9'd3,10'd197};
ram[33732] = {9'd0,10'd201};
ram[33733] = {9'd3,10'd204};
ram[33734] = {9'd7,10'd207};
ram[33735] = {9'd10,10'd210};
ram[33736] = {9'd13,10'd213};
ram[33737] = {9'd16,10'd216};
ram[33738] = {9'd19,10'd219};
ram[33739] = {9'd22,10'd223};
ram[33740] = {9'd25,10'd226};
ram[33741] = {9'd29,10'd229};
ram[33742] = {9'd32,10'd232};
ram[33743] = {9'd35,10'd235};
ram[33744] = {9'd38,10'd238};
ram[33745] = {9'd41,10'd241};
ram[33746] = {9'd44,10'd245};
ram[33747] = {9'd47,10'd248};
ram[33748] = {9'd51,10'd251};
ram[33749] = {9'd54,10'd254};
ram[33750] = {9'd57,10'd257};
ram[33751] = {9'd60,10'd260};
ram[33752] = {9'd63,10'd263};
ram[33753] = {9'd66,10'd267};
ram[33754] = {9'd69,10'd270};
ram[33755] = {9'd73,10'd273};
ram[33756] = {9'd76,10'd276};
ram[33757] = {9'd79,10'd279};
ram[33758] = {9'd82,10'd282};
ram[33759] = {9'd85,10'd285};
ram[33760] = {9'd88,10'd289};
ram[33761] = {9'd91,10'd292};
ram[33762] = {9'd95,10'd295};
ram[33763] = {9'd98,10'd298};
ram[33764] = {-9'd99,10'd301};
ram[33765] = {-9'd96,10'd304};
ram[33766] = {-9'd93,10'd307};
ram[33767] = {-9'd90,10'd311};
ram[33768] = {-9'd87,10'd314};
ram[33769] = {-9'd84,10'd317};
ram[33770] = {-9'd81,10'd320};
ram[33771] = {-9'd77,10'd323};
ram[33772] = {-9'd74,10'd326};
ram[33773] = {-9'd71,10'd329};
ram[33774] = {-9'd68,10'd333};
ram[33775] = {-9'd65,10'd336};
ram[33776] = {-9'd62,10'd339};
ram[33777] = {-9'd59,10'd342};
ram[33778] = {-9'd55,10'd345};
ram[33779] = {-9'd52,10'd348};
ram[33780] = {-9'd49,10'd351};
ram[33781] = {-9'd46,10'd354};
ram[33782] = {-9'd43,10'd358};
ram[33783] = {-9'd40,10'd361};
ram[33784] = {-9'd37,10'd364};
ram[33785] = {-9'd33,10'd367};
ram[33786] = {-9'd30,10'd370};
ram[33787] = {-9'd27,10'd373};
ram[33788] = {-9'd24,10'd376};
ram[33789] = {-9'd21,10'd380};
ram[33790] = {-9'd18,10'd383};
ram[33791] = {-9'd15,10'd386};
ram[33792] = {-9'd15,10'd386};
ram[33793] = {-9'd11,10'd389};
ram[33794] = {-9'd8,10'd392};
ram[33795] = {-9'd5,10'd395};
ram[33796] = {-9'd2,10'd398};
ram[33797] = {9'd1,-10'd399};
ram[33798] = {9'd4,-10'd396};
ram[33799] = {9'd7,-10'd393};
ram[33800] = {9'd10,-10'd390};
ram[33801] = {9'd14,-10'd387};
ram[33802] = {9'd17,-10'd384};
ram[33803] = {9'd20,-10'd381};
ram[33804] = {9'd23,-10'd377};
ram[33805] = {9'd26,-10'd374};
ram[33806] = {9'd29,-10'd371};
ram[33807] = {9'd32,-10'd368};
ram[33808] = {9'd36,-10'd365};
ram[33809] = {9'd39,-10'd362};
ram[33810] = {9'd42,-10'd359};
ram[33811] = {9'd45,-10'd355};
ram[33812] = {9'd48,-10'd352};
ram[33813] = {9'd51,-10'd349};
ram[33814] = {9'd54,-10'd346};
ram[33815] = {9'd58,-10'd343};
ram[33816] = {9'd61,-10'd340};
ram[33817] = {9'd64,-10'd337};
ram[33818] = {9'd67,-10'd334};
ram[33819] = {9'd70,-10'd330};
ram[33820] = {9'd73,-10'd327};
ram[33821] = {9'd76,-10'd324};
ram[33822] = {9'd80,-10'd321};
ram[33823] = {9'd83,-10'd318};
ram[33824] = {9'd86,-10'd315};
ram[33825] = {9'd89,-10'd312};
ram[33826] = {9'd92,-10'd308};
ram[33827] = {9'd95,-10'd305};
ram[33828] = {9'd98,-10'd302};
ram[33829] = {-9'd99,-10'd299};
ram[33830] = {-9'd96,-10'd296};
ram[33831] = {-9'd92,-10'd293};
ram[33832] = {-9'd89,-10'd290};
ram[33833] = {-9'd86,-10'd286};
ram[33834] = {-9'd83,-10'd283};
ram[33835] = {-9'd80,-10'd280};
ram[33836] = {-9'd77,-10'd277};
ram[33837] = {-9'd74,-10'd274};
ram[33838] = {-9'd70,-10'd271};
ram[33839] = {-9'd67,-10'd268};
ram[33840] = {-9'd64,-10'd264};
ram[33841] = {-9'd61,-10'd261};
ram[33842] = {-9'd58,-10'd258};
ram[33843] = {-9'd55,-10'd255};
ram[33844] = {-9'd52,-10'd252};
ram[33845] = {-9'd48,-10'd249};
ram[33846] = {-9'd45,-10'd246};
ram[33847] = {-9'd42,-10'd242};
ram[33848] = {-9'd39,-10'd239};
ram[33849] = {-9'd36,-10'd236};
ram[33850] = {-9'd33,-10'd233};
ram[33851] = {-9'd30,-10'd230};
ram[33852] = {-9'd26,-10'd227};
ram[33853] = {-9'd23,-10'd224};
ram[33854] = {-9'd20,-10'd220};
ram[33855] = {-9'd17,-10'd217};
ram[33856] = {-9'd14,-10'd214};
ram[33857] = {-9'd11,-10'd211};
ram[33858] = {-9'd8,-10'd208};
ram[33859] = {-9'd4,-10'd205};
ram[33860] = {-9'd1,-10'd202};
ram[33861] = {9'd2,-10'd198};
ram[33862] = {9'd5,-10'd195};
ram[33863] = {9'd8,-10'd192};
ram[33864] = {9'd11,-10'd189};
ram[33865] = {9'd14,-10'd186};
ram[33866] = {9'd18,-10'd183};
ram[33867] = {9'd21,-10'd180};
ram[33868] = {9'd24,-10'd176};
ram[33869] = {9'd27,-10'd173};
ram[33870] = {9'd30,-10'd170};
ram[33871] = {9'd33,-10'd167};
ram[33872] = {9'd36,-10'd164};
ram[33873] = {9'd40,-10'd161};
ram[33874] = {9'd43,-10'd158};
ram[33875] = {9'd46,-10'd154};
ram[33876] = {9'd49,-10'd151};
ram[33877] = {9'd52,-10'd148};
ram[33878] = {9'd55,-10'd145};
ram[33879] = {9'd58,-10'd142};
ram[33880] = {9'd62,-10'd139};
ram[33881] = {9'd65,-10'd136};
ram[33882] = {9'd68,-10'd132};
ram[33883] = {9'd71,-10'd129};
ram[33884] = {9'd74,-10'd126};
ram[33885] = {9'd77,-10'd123};
ram[33886] = {9'd80,-10'd120};
ram[33887] = {9'd84,-10'd117};
ram[33888] = {9'd87,-10'd114};
ram[33889] = {9'd90,-10'd110};
ram[33890] = {9'd93,-10'd107};
ram[33891] = {9'd96,-10'd104};
ram[33892] = {9'd99,-10'd101};
ram[33893] = {-9'd98,-10'd98};
ram[33894] = {-9'd95,-10'd95};
ram[33895] = {-9'd92,-10'd92};
ram[33896] = {-9'd88,-10'd88};
ram[33897] = {-9'd85,-10'd85};
ram[33898] = {-9'd82,-10'd82};
ram[33899] = {-9'd79,-10'd79};
ram[33900] = {-9'd76,-10'd76};
ram[33901] = {-9'd73,-10'd73};
ram[33902] = {-9'd70,-10'd70};
ram[33903] = {-9'd66,-10'd66};
ram[33904] = {-9'd63,-10'd63};
ram[33905] = {-9'd60,-10'd60};
ram[33906] = {-9'd57,-10'd57};
ram[33907] = {-9'd54,-10'd54};
ram[33908] = {-9'd51,-10'd51};
ram[33909] = {-9'd48,-10'd48};
ram[33910] = {-9'd44,-10'd44};
ram[33911] = {-9'd41,-10'd41};
ram[33912] = {-9'd38,-10'd38};
ram[33913] = {-9'd35,-10'd35};
ram[33914] = {-9'd32,-10'd32};
ram[33915] = {-9'd29,-10'd29};
ram[33916] = {-9'd26,-10'd26};
ram[33917] = {-9'd22,-10'd22};
ram[33918] = {-9'd19,-10'd19};
ram[33919] = {-9'd16,-10'd16};
ram[33920] = {-9'd16,-10'd16};
ram[33921] = {-9'd13,-10'd13};
ram[33922] = {-9'd10,-10'd10};
ram[33923] = {-9'd7,-10'd7};
ram[33924] = {-9'd4,-10'd4};
ram[33925] = {9'd0,10'd0};
ram[33926] = {9'd3,10'd3};
ram[33927] = {9'd6,10'd6};
ram[33928] = {9'd9,10'd9};
ram[33929] = {9'd12,10'd12};
ram[33930] = {9'd15,10'd15};
ram[33931] = {9'd18,10'd18};
ram[33932] = {9'd21,10'd21};
ram[33933] = {9'd25,10'd25};
ram[33934] = {9'd28,10'd28};
ram[33935] = {9'd31,10'd31};
ram[33936] = {9'd34,10'd34};
ram[33937] = {9'd37,10'd37};
ram[33938] = {9'd40,10'd40};
ram[33939] = {9'd43,10'd43};
ram[33940] = {9'd47,10'd47};
ram[33941] = {9'd50,10'd50};
ram[33942] = {9'd53,10'd53};
ram[33943] = {9'd56,10'd56};
ram[33944] = {9'd59,10'd59};
ram[33945] = {9'd62,10'd62};
ram[33946] = {9'd65,10'd65};
ram[33947] = {9'd69,10'd69};
ram[33948] = {9'd72,10'd72};
ram[33949] = {9'd75,10'd75};
ram[33950] = {9'd78,10'd78};
ram[33951] = {9'd81,10'd81};
ram[33952] = {9'd84,10'd84};
ram[33953] = {9'd87,10'd87};
ram[33954] = {9'd91,10'd91};
ram[33955] = {9'd94,10'd94};
ram[33956] = {9'd97,10'd97};
ram[33957] = {-9'd100,10'd100};
ram[33958] = {-9'd97,10'd103};
ram[33959] = {-9'd94,10'd106};
ram[33960] = {-9'd91,10'd109};
ram[33961] = {-9'd88,10'd113};
ram[33962] = {-9'd85,10'd116};
ram[33963] = {-9'd81,10'd119};
ram[33964] = {-9'd78,10'd122};
ram[33965] = {-9'd75,10'd125};
ram[33966] = {-9'd72,10'd128};
ram[33967] = {-9'd69,10'd131};
ram[33968] = {-9'd66,10'd135};
ram[33969] = {-9'd63,10'd138};
ram[33970] = {-9'd59,10'd141};
ram[33971] = {-9'd56,10'd144};
ram[33972] = {-9'd53,10'd147};
ram[33973] = {-9'd50,10'd150};
ram[33974] = {-9'd47,10'd153};
ram[33975] = {-9'd44,10'd157};
ram[33976] = {-9'd41,10'd160};
ram[33977] = {-9'd37,10'd163};
ram[33978] = {-9'd34,10'd166};
ram[33979] = {-9'd31,10'd169};
ram[33980] = {-9'd28,10'd172};
ram[33981] = {-9'd25,10'd175};
ram[33982] = {-9'd22,10'd179};
ram[33983] = {-9'd19,10'd182};
ram[33984] = {-9'd15,10'd185};
ram[33985] = {-9'd12,10'd188};
ram[33986] = {-9'd9,10'd191};
ram[33987] = {-9'd6,10'd194};
ram[33988] = {-9'd3,10'd197};
ram[33989] = {9'd0,10'd201};
ram[33990] = {9'd3,10'd204};
ram[33991] = {9'd7,10'd207};
ram[33992] = {9'd10,10'd210};
ram[33993] = {9'd13,10'd213};
ram[33994] = {9'd16,10'd216};
ram[33995] = {9'd19,10'd219};
ram[33996] = {9'd22,10'd223};
ram[33997] = {9'd25,10'd226};
ram[33998] = {9'd29,10'd229};
ram[33999] = {9'd32,10'd232};
ram[34000] = {9'd35,10'd235};
ram[34001] = {9'd38,10'd238};
ram[34002] = {9'd41,10'd241};
ram[34003] = {9'd44,10'd245};
ram[34004] = {9'd47,10'd248};
ram[34005] = {9'd51,10'd251};
ram[34006] = {9'd54,10'd254};
ram[34007] = {9'd57,10'd257};
ram[34008] = {9'd60,10'd260};
ram[34009] = {9'd63,10'd263};
ram[34010] = {9'd66,10'd267};
ram[34011] = {9'd69,10'd270};
ram[34012] = {9'd73,10'd273};
ram[34013] = {9'd76,10'd276};
ram[34014] = {9'd79,10'd279};
ram[34015] = {9'd82,10'd282};
ram[34016] = {9'd85,10'd285};
ram[34017] = {9'd88,10'd289};
ram[34018] = {9'd91,10'd292};
ram[34019] = {9'd95,10'd295};
ram[34020] = {9'd98,10'd298};
ram[34021] = {-9'd99,10'd301};
ram[34022] = {-9'd96,10'd304};
ram[34023] = {-9'd93,10'd307};
ram[34024] = {-9'd90,10'd311};
ram[34025] = {-9'd87,10'd314};
ram[34026] = {-9'd84,10'd317};
ram[34027] = {-9'd81,10'd320};
ram[34028] = {-9'd77,10'd323};
ram[34029] = {-9'd74,10'd326};
ram[34030] = {-9'd71,10'd329};
ram[34031] = {-9'd68,10'd333};
ram[34032] = {-9'd65,10'd336};
ram[34033] = {-9'd62,10'd339};
ram[34034] = {-9'd59,10'd342};
ram[34035] = {-9'd55,10'd345};
ram[34036] = {-9'd52,10'd348};
ram[34037] = {-9'd49,10'd351};
ram[34038] = {-9'd46,10'd354};
ram[34039] = {-9'd43,10'd358};
ram[34040] = {-9'd40,10'd361};
ram[34041] = {-9'd37,10'd364};
ram[34042] = {-9'd33,10'd367};
ram[34043] = {-9'd30,10'd370};
ram[34044] = {-9'd27,10'd373};
ram[34045] = {-9'd24,10'd376};
ram[34046] = {-9'd21,10'd380};
ram[34047] = {-9'd18,10'd383};
ram[34048] = {-9'd18,10'd383};
ram[34049] = {-9'd15,10'd386};
ram[34050] = {-9'd11,10'd389};
ram[34051] = {-9'd8,10'd392};
ram[34052] = {-9'd5,10'd395};
ram[34053] = {-9'd2,10'd398};
ram[34054] = {9'd1,-10'd399};
ram[34055] = {9'd4,-10'd396};
ram[34056] = {9'd7,-10'd393};
ram[34057] = {9'd10,-10'd390};
ram[34058] = {9'd14,-10'd387};
ram[34059] = {9'd17,-10'd384};
ram[34060] = {9'd20,-10'd381};
ram[34061] = {9'd23,-10'd377};
ram[34062] = {9'd26,-10'd374};
ram[34063] = {9'd29,-10'd371};
ram[34064] = {9'd32,-10'd368};
ram[34065] = {9'd36,-10'd365};
ram[34066] = {9'd39,-10'd362};
ram[34067] = {9'd42,-10'd359};
ram[34068] = {9'd45,-10'd355};
ram[34069] = {9'd48,-10'd352};
ram[34070] = {9'd51,-10'd349};
ram[34071] = {9'd54,-10'd346};
ram[34072] = {9'd58,-10'd343};
ram[34073] = {9'd61,-10'd340};
ram[34074] = {9'd64,-10'd337};
ram[34075] = {9'd67,-10'd334};
ram[34076] = {9'd70,-10'd330};
ram[34077] = {9'd73,-10'd327};
ram[34078] = {9'd76,-10'd324};
ram[34079] = {9'd80,-10'd321};
ram[34080] = {9'd83,-10'd318};
ram[34081] = {9'd86,-10'd315};
ram[34082] = {9'd89,-10'd312};
ram[34083] = {9'd92,-10'd308};
ram[34084] = {9'd95,-10'd305};
ram[34085] = {9'd98,-10'd302};
ram[34086] = {-9'd99,-10'd299};
ram[34087] = {-9'd96,-10'd296};
ram[34088] = {-9'd92,-10'd293};
ram[34089] = {-9'd89,-10'd290};
ram[34090] = {-9'd86,-10'd286};
ram[34091] = {-9'd83,-10'd283};
ram[34092] = {-9'd80,-10'd280};
ram[34093] = {-9'd77,-10'd277};
ram[34094] = {-9'd74,-10'd274};
ram[34095] = {-9'd70,-10'd271};
ram[34096] = {-9'd67,-10'd268};
ram[34097] = {-9'd64,-10'd264};
ram[34098] = {-9'd61,-10'd261};
ram[34099] = {-9'd58,-10'd258};
ram[34100] = {-9'd55,-10'd255};
ram[34101] = {-9'd52,-10'd252};
ram[34102] = {-9'd48,-10'd249};
ram[34103] = {-9'd45,-10'd246};
ram[34104] = {-9'd42,-10'd242};
ram[34105] = {-9'd39,-10'd239};
ram[34106] = {-9'd36,-10'd236};
ram[34107] = {-9'd33,-10'd233};
ram[34108] = {-9'd30,-10'd230};
ram[34109] = {-9'd26,-10'd227};
ram[34110] = {-9'd23,-10'd224};
ram[34111] = {-9'd20,-10'd220};
ram[34112] = {-9'd17,-10'd217};
ram[34113] = {-9'd14,-10'd214};
ram[34114] = {-9'd11,-10'd211};
ram[34115] = {-9'd8,-10'd208};
ram[34116] = {-9'd4,-10'd205};
ram[34117] = {-9'd1,-10'd202};
ram[34118] = {9'd2,-10'd198};
ram[34119] = {9'd5,-10'd195};
ram[34120] = {9'd8,-10'd192};
ram[34121] = {9'd11,-10'd189};
ram[34122] = {9'd14,-10'd186};
ram[34123] = {9'd18,-10'd183};
ram[34124] = {9'd21,-10'd180};
ram[34125] = {9'd24,-10'd176};
ram[34126] = {9'd27,-10'd173};
ram[34127] = {9'd30,-10'd170};
ram[34128] = {9'd33,-10'd167};
ram[34129] = {9'd36,-10'd164};
ram[34130] = {9'd40,-10'd161};
ram[34131] = {9'd43,-10'd158};
ram[34132] = {9'd46,-10'd154};
ram[34133] = {9'd49,-10'd151};
ram[34134] = {9'd52,-10'd148};
ram[34135] = {9'd55,-10'd145};
ram[34136] = {9'd58,-10'd142};
ram[34137] = {9'd62,-10'd139};
ram[34138] = {9'd65,-10'd136};
ram[34139] = {9'd68,-10'd132};
ram[34140] = {9'd71,-10'd129};
ram[34141] = {9'd74,-10'd126};
ram[34142] = {9'd77,-10'd123};
ram[34143] = {9'd80,-10'd120};
ram[34144] = {9'd84,-10'd117};
ram[34145] = {9'd87,-10'd114};
ram[34146] = {9'd90,-10'd110};
ram[34147] = {9'd93,-10'd107};
ram[34148] = {9'd96,-10'd104};
ram[34149] = {9'd99,-10'd101};
ram[34150] = {-9'd98,-10'd98};
ram[34151] = {-9'd95,-10'd95};
ram[34152] = {-9'd92,-10'd92};
ram[34153] = {-9'd88,-10'd88};
ram[34154] = {-9'd85,-10'd85};
ram[34155] = {-9'd82,-10'd82};
ram[34156] = {-9'd79,-10'd79};
ram[34157] = {-9'd76,-10'd76};
ram[34158] = {-9'd73,-10'd73};
ram[34159] = {-9'd70,-10'd70};
ram[34160] = {-9'd66,-10'd66};
ram[34161] = {-9'd63,-10'd63};
ram[34162] = {-9'd60,-10'd60};
ram[34163] = {-9'd57,-10'd57};
ram[34164] = {-9'd54,-10'd54};
ram[34165] = {-9'd51,-10'd51};
ram[34166] = {-9'd48,-10'd48};
ram[34167] = {-9'd44,-10'd44};
ram[34168] = {-9'd41,-10'd41};
ram[34169] = {-9'd38,-10'd38};
ram[34170] = {-9'd35,-10'd35};
ram[34171] = {-9'd32,-10'd32};
ram[34172] = {-9'd29,-10'd29};
ram[34173] = {-9'd26,-10'd26};
ram[34174] = {-9'd22,-10'd22};
ram[34175] = {-9'd19,-10'd19};
ram[34176] = {-9'd19,-10'd19};
ram[34177] = {-9'd16,-10'd16};
ram[34178] = {-9'd13,-10'd13};
ram[34179] = {-9'd10,-10'd10};
ram[34180] = {-9'd7,-10'd7};
ram[34181] = {-9'd4,-10'd4};
ram[34182] = {9'd0,10'd0};
ram[34183] = {9'd3,10'd3};
ram[34184] = {9'd6,10'd6};
ram[34185] = {9'd9,10'd9};
ram[34186] = {9'd12,10'd12};
ram[34187] = {9'd15,10'd15};
ram[34188] = {9'd18,10'd18};
ram[34189] = {9'd21,10'd21};
ram[34190] = {9'd25,10'd25};
ram[34191] = {9'd28,10'd28};
ram[34192] = {9'd31,10'd31};
ram[34193] = {9'd34,10'd34};
ram[34194] = {9'd37,10'd37};
ram[34195] = {9'd40,10'd40};
ram[34196] = {9'd43,10'd43};
ram[34197] = {9'd47,10'd47};
ram[34198] = {9'd50,10'd50};
ram[34199] = {9'd53,10'd53};
ram[34200] = {9'd56,10'd56};
ram[34201] = {9'd59,10'd59};
ram[34202] = {9'd62,10'd62};
ram[34203] = {9'd65,10'd65};
ram[34204] = {9'd69,10'd69};
ram[34205] = {9'd72,10'd72};
ram[34206] = {9'd75,10'd75};
ram[34207] = {9'd78,10'd78};
ram[34208] = {9'd81,10'd81};
ram[34209] = {9'd84,10'd84};
ram[34210] = {9'd87,10'd87};
ram[34211] = {9'd91,10'd91};
ram[34212] = {9'd94,10'd94};
ram[34213] = {9'd97,10'd97};
ram[34214] = {-9'd100,10'd100};
ram[34215] = {-9'd97,10'd103};
ram[34216] = {-9'd94,10'd106};
ram[34217] = {-9'd91,10'd109};
ram[34218] = {-9'd88,10'd113};
ram[34219] = {-9'd85,10'd116};
ram[34220] = {-9'd81,10'd119};
ram[34221] = {-9'd78,10'd122};
ram[34222] = {-9'd75,10'd125};
ram[34223] = {-9'd72,10'd128};
ram[34224] = {-9'd69,10'd131};
ram[34225] = {-9'd66,10'd135};
ram[34226] = {-9'd63,10'd138};
ram[34227] = {-9'd59,10'd141};
ram[34228] = {-9'd56,10'd144};
ram[34229] = {-9'd53,10'd147};
ram[34230] = {-9'd50,10'd150};
ram[34231] = {-9'd47,10'd153};
ram[34232] = {-9'd44,10'd157};
ram[34233] = {-9'd41,10'd160};
ram[34234] = {-9'd37,10'd163};
ram[34235] = {-9'd34,10'd166};
ram[34236] = {-9'd31,10'd169};
ram[34237] = {-9'd28,10'd172};
ram[34238] = {-9'd25,10'd175};
ram[34239] = {-9'd22,10'd179};
ram[34240] = {-9'd19,10'd182};
ram[34241] = {-9'd15,10'd185};
ram[34242] = {-9'd12,10'd188};
ram[34243] = {-9'd9,10'd191};
ram[34244] = {-9'd6,10'd194};
ram[34245] = {-9'd3,10'd197};
ram[34246] = {9'd0,10'd201};
ram[34247] = {9'd3,10'd204};
ram[34248] = {9'd7,10'd207};
ram[34249] = {9'd10,10'd210};
ram[34250] = {9'd13,10'd213};
ram[34251] = {9'd16,10'd216};
ram[34252] = {9'd19,10'd219};
ram[34253] = {9'd22,10'd223};
ram[34254] = {9'd25,10'd226};
ram[34255] = {9'd29,10'd229};
ram[34256] = {9'd32,10'd232};
ram[34257] = {9'd35,10'd235};
ram[34258] = {9'd38,10'd238};
ram[34259] = {9'd41,10'd241};
ram[34260] = {9'd44,10'd245};
ram[34261] = {9'd47,10'd248};
ram[34262] = {9'd51,10'd251};
ram[34263] = {9'd54,10'd254};
ram[34264] = {9'd57,10'd257};
ram[34265] = {9'd60,10'd260};
ram[34266] = {9'd63,10'd263};
ram[34267] = {9'd66,10'd267};
ram[34268] = {9'd69,10'd270};
ram[34269] = {9'd73,10'd273};
ram[34270] = {9'd76,10'd276};
ram[34271] = {9'd79,10'd279};
ram[34272] = {9'd82,10'd282};
ram[34273] = {9'd85,10'd285};
ram[34274] = {9'd88,10'd289};
ram[34275] = {9'd91,10'd292};
ram[34276] = {9'd95,10'd295};
ram[34277] = {9'd98,10'd298};
ram[34278] = {-9'd99,10'd301};
ram[34279] = {-9'd96,10'd304};
ram[34280] = {-9'd93,10'd307};
ram[34281] = {-9'd90,10'd311};
ram[34282] = {-9'd87,10'd314};
ram[34283] = {-9'd84,10'd317};
ram[34284] = {-9'd81,10'd320};
ram[34285] = {-9'd77,10'd323};
ram[34286] = {-9'd74,10'd326};
ram[34287] = {-9'd71,10'd329};
ram[34288] = {-9'd68,10'd333};
ram[34289] = {-9'd65,10'd336};
ram[34290] = {-9'd62,10'd339};
ram[34291] = {-9'd59,10'd342};
ram[34292] = {-9'd55,10'd345};
ram[34293] = {-9'd52,10'd348};
ram[34294] = {-9'd49,10'd351};
ram[34295] = {-9'd46,10'd354};
ram[34296] = {-9'd43,10'd358};
ram[34297] = {-9'd40,10'd361};
ram[34298] = {-9'd37,10'd364};
ram[34299] = {-9'd33,10'd367};
ram[34300] = {-9'd30,10'd370};
ram[34301] = {-9'd27,10'd373};
ram[34302] = {-9'd24,10'd376};
ram[34303] = {-9'd21,10'd380};
ram[34304] = {-9'd21,10'd380};
ram[34305] = {-9'd18,10'd383};
ram[34306] = {-9'd15,10'd386};
ram[34307] = {-9'd11,10'd389};
ram[34308] = {-9'd8,10'd392};
ram[34309] = {-9'd5,10'd395};
ram[34310] = {-9'd2,10'd398};
ram[34311] = {9'd1,-10'd399};
ram[34312] = {9'd4,-10'd396};
ram[34313] = {9'd7,-10'd393};
ram[34314] = {9'd10,-10'd390};
ram[34315] = {9'd14,-10'd387};
ram[34316] = {9'd17,-10'd384};
ram[34317] = {9'd20,-10'd381};
ram[34318] = {9'd23,-10'd377};
ram[34319] = {9'd26,-10'd374};
ram[34320] = {9'd29,-10'd371};
ram[34321] = {9'd32,-10'd368};
ram[34322] = {9'd36,-10'd365};
ram[34323] = {9'd39,-10'd362};
ram[34324] = {9'd42,-10'd359};
ram[34325] = {9'd45,-10'd355};
ram[34326] = {9'd48,-10'd352};
ram[34327] = {9'd51,-10'd349};
ram[34328] = {9'd54,-10'd346};
ram[34329] = {9'd58,-10'd343};
ram[34330] = {9'd61,-10'd340};
ram[34331] = {9'd64,-10'd337};
ram[34332] = {9'd67,-10'd334};
ram[34333] = {9'd70,-10'd330};
ram[34334] = {9'd73,-10'd327};
ram[34335] = {9'd76,-10'd324};
ram[34336] = {9'd80,-10'd321};
ram[34337] = {9'd83,-10'd318};
ram[34338] = {9'd86,-10'd315};
ram[34339] = {9'd89,-10'd312};
ram[34340] = {9'd92,-10'd308};
ram[34341] = {9'd95,-10'd305};
ram[34342] = {9'd98,-10'd302};
ram[34343] = {-9'd99,-10'd299};
ram[34344] = {-9'd96,-10'd296};
ram[34345] = {-9'd92,-10'd293};
ram[34346] = {-9'd89,-10'd290};
ram[34347] = {-9'd86,-10'd286};
ram[34348] = {-9'd83,-10'd283};
ram[34349] = {-9'd80,-10'd280};
ram[34350] = {-9'd77,-10'd277};
ram[34351] = {-9'd74,-10'd274};
ram[34352] = {-9'd70,-10'd271};
ram[34353] = {-9'd67,-10'd268};
ram[34354] = {-9'd64,-10'd264};
ram[34355] = {-9'd61,-10'd261};
ram[34356] = {-9'd58,-10'd258};
ram[34357] = {-9'd55,-10'd255};
ram[34358] = {-9'd52,-10'd252};
ram[34359] = {-9'd48,-10'd249};
ram[34360] = {-9'd45,-10'd246};
ram[34361] = {-9'd42,-10'd242};
ram[34362] = {-9'd39,-10'd239};
ram[34363] = {-9'd36,-10'd236};
ram[34364] = {-9'd33,-10'd233};
ram[34365] = {-9'd30,-10'd230};
ram[34366] = {-9'd26,-10'd227};
ram[34367] = {-9'd23,-10'd224};
ram[34368] = {-9'd20,-10'd220};
ram[34369] = {-9'd17,-10'd217};
ram[34370] = {-9'd14,-10'd214};
ram[34371] = {-9'd11,-10'd211};
ram[34372] = {-9'd8,-10'd208};
ram[34373] = {-9'd4,-10'd205};
ram[34374] = {-9'd1,-10'd202};
ram[34375] = {9'd2,-10'd198};
ram[34376] = {9'd5,-10'd195};
ram[34377] = {9'd8,-10'd192};
ram[34378] = {9'd11,-10'd189};
ram[34379] = {9'd14,-10'd186};
ram[34380] = {9'd18,-10'd183};
ram[34381] = {9'd21,-10'd180};
ram[34382] = {9'd24,-10'd176};
ram[34383] = {9'd27,-10'd173};
ram[34384] = {9'd30,-10'd170};
ram[34385] = {9'd33,-10'd167};
ram[34386] = {9'd36,-10'd164};
ram[34387] = {9'd40,-10'd161};
ram[34388] = {9'd43,-10'd158};
ram[34389] = {9'd46,-10'd154};
ram[34390] = {9'd49,-10'd151};
ram[34391] = {9'd52,-10'd148};
ram[34392] = {9'd55,-10'd145};
ram[34393] = {9'd58,-10'd142};
ram[34394] = {9'd62,-10'd139};
ram[34395] = {9'd65,-10'd136};
ram[34396] = {9'd68,-10'd132};
ram[34397] = {9'd71,-10'd129};
ram[34398] = {9'd74,-10'd126};
ram[34399] = {9'd77,-10'd123};
ram[34400] = {9'd80,-10'd120};
ram[34401] = {9'd84,-10'd117};
ram[34402] = {9'd87,-10'd114};
ram[34403] = {9'd90,-10'd110};
ram[34404] = {9'd93,-10'd107};
ram[34405] = {9'd96,-10'd104};
ram[34406] = {9'd99,-10'd101};
ram[34407] = {-9'd98,-10'd98};
ram[34408] = {-9'd95,-10'd95};
ram[34409] = {-9'd92,-10'd92};
ram[34410] = {-9'd88,-10'd88};
ram[34411] = {-9'd85,-10'd85};
ram[34412] = {-9'd82,-10'd82};
ram[34413] = {-9'd79,-10'd79};
ram[34414] = {-9'd76,-10'd76};
ram[34415] = {-9'd73,-10'd73};
ram[34416] = {-9'd70,-10'd70};
ram[34417] = {-9'd66,-10'd66};
ram[34418] = {-9'd63,-10'd63};
ram[34419] = {-9'd60,-10'd60};
ram[34420] = {-9'd57,-10'd57};
ram[34421] = {-9'd54,-10'd54};
ram[34422] = {-9'd51,-10'd51};
ram[34423] = {-9'd48,-10'd48};
ram[34424] = {-9'd44,-10'd44};
ram[34425] = {-9'd41,-10'd41};
ram[34426] = {-9'd38,-10'd38};
ram[34427] = {-9'd35,-10'd35};
ram[34428] = {-9'd32,-10'd32};
ram[34429] = {-9'd29,-10'd29};
ram[34430] = {-9'd26,-10'd26};
ram[34431] = {-9'd22,-10'd22};
ram[34432] = {-9'd22,-10'd22};
ram[34433] = {-9'd19,-10'd19};
ram[34434] = {-9'd16,-10'd16};
ram[34435] = {-9'd13,-10'd13};
ram[34436] = {-9'd10,-10'd10};
ram[34437] = {-9'd7,-10'd7};
ram[34438] = {-9'd4,-10'd4};
ram[34439] = {9'd0,10'd0};
ram[34440] = {9'd3,10'd3};
ram[34441] = {9'd6,10'd6};
ram[34442] = {9'd9,10'd9};
ram[34443] = {9'd12,10'd12};
ram[34444] = {9'd15,10'd15};
ram[34445] = {9'd18,10'd18};
ram[34446] = {9'd21,10'd21};
ram[34447] = {9'd25,10'd25};
ram[34448] = {9'd28,10'd28};
ram[34449] = {9'd31,10'd31};
ram[34450] = {9'd34,10'd34};
ram[34451] = {9'd37,10'd37};
ram[34452] = {9'd40,10'd40};
ram[34453] = {9'd43,10'd43};
ram[34454] = {9'd47,10'd47};
ram[34455] = {9'd50,10'd50};
ram[34456] = {9'd53,10'd53};
ram[34457] = {9'd56,10'd56};
ram[34458] = {9'd59,10'd59};
ram[34459] = {9'd62,10'd62};
ram[34460] = {9'd65,10'd65};
ram[34461] = {9'd69,10'd69};
ram[34462] = {9'd72,10'd72};
ram[34463] = {9'd75,10'd75};
ram[34464] = {9'd78,10'd78};
ram[34465] = {9'd81,10'd81};
ram[34466] = {9'd84,10'd84};
ram[34467] = {9'd87,10'd87};
ram[34468] = {9'd91,10'd91};
ram[34469] = {9'd94,10'd94};
ram[34470] = {9'd97,10'd97};
ram[34471] = {-9'd100,10'd100};
ram[34472] = {-9'd97,10'd103};
ram[34473] = {-9'd94,10'd106};
ram[34474] = {-9'd91,10'd109};
ram[34475] = {-9'd88,10'd113};
ram[34476] = {-9'd85,10'd116};
ram[34477] = {-9'd81,10'd119};
ram[34478] = {-9'd78,10'd122};
ram[34479] = {-9'd75,10'd125};
ram[34480] = {-9'd72,10'd128};
ram[34481] = {-9'd69,10'd131};
ram[34482] = {-9'd66,10'd135};
ram[34483] = {-9'd63,10'd138};
ram[34484] = {-9'd59,10'd141};
ram[34485] = {-9'd56,10'd144};
ram[34486] = {-9'd53,10'd147};
ram[34487] = {-9'd50,10'd150};
ram[34488] = {-9'd47,10'd153};
ram[34489] = {-9'd44,10'd157};
ram[34490] = {-9'd41,10'd160};
ram[34491] = {-9'd37,10'd163};
ram[34492] = {-9'd34,10'd166};
ram[34493] = {-9'd31,10'd169};
ram[34494] = {-9'd28,10'd172};
ram[34495] = {-9'd25,10'd175};
ram[34496] = {-9'd22,10'd179};
ram[34497] = {-9'd19,10'd182};
ram[34498] = {-9'd15,10'd185};
ram[34499] = {-9'd12,10'd188};
ram[34500] = {-9'd9,10'd191};
ram[34501] = {-9'd6,10'd194};
ram[34502] = {-9'd3,10'd197};
ram[34503] = {9'd0,10'd201};
ram[34504] = {9'd3,10'd204};
ram[34505] = {9'd7,10'd207};
ram[34506] = {9'd10,10'd210};
ram[34507] = {9'd13,10'd213};
ram[34508] = {9'd16,10'd216};
ram[34509] = {9'd19,10'd219};
ram[34510] = {9'd22,10'd223};
ram[34511] = {9'd25,10'd226};
ram[34512] = {9'd29,10'd229};
ram[34513] = {9'd32,10'd232};
ram[34514] = {9'd35,10'd235};
ram[34515] = {9'd38,10'd238};
ram[34516] = {9'd41,10'd241};
ram[34517] = {9'd44,10'd245};
ram[34518] = {9'd47,10'd248};
ram[34519] = {9'd51,10'd251};
ram[34520] = {9'd54,10'd254};
ram[34521] = {9'd57,10'd257};
ram[34522] = {9'd60,10'd260};
ram[34523] = {9'd63,10'd263};
ram[34524] = {9'd66,10'd267};
ram[34525] = {9'd69,10'd270};
ram[34526] = {9'd73,10'd273};
ram[34527] = {9'd76,10'd276};
ram[34528] = {9'd79,10'd279};
ram[34529] = {9'd82,10'd282};
ram[34530] = {9'd85,10'd285};
ram[34531] = {9'd88,10'd289};
ram[34532] = {9'd91,10'd292};
ram[34533] = {9'd95,10'd295};
ram[34534] = {9'd98,10'd298};
ram[34535] = {-9'd99,10'd301};
ram[34536] = {-9'd96,10'd304};
ram[34537] = {-9'd93,10'd307};
ram[34538] = {-9'd90,10'd311};
ram[34539] = {-9'd87,10'd314};
ram[34540] = {-9'd84,10'd317};
ram[34541] = {-9'd81,10'd320};
ram[34542] = {-9'd77,10'd323};
ram[34543] = {-9'd74,10'd326};
ram[34544] = {-9'd71,10'd329};
ram[34545] = {-9'd68,10'd333};
ram[34546] = {-9'd65,10'd336};
ram[34547] = {-9'd62,10'd339};
ram[34548] = {-9'd59,10'd342};
ram[34549] = {-9'd55,10'd345};
ram[34550] = {-9'd52,10'd348};
ram[34551] = {-9'd49,10'd351};
ram[34552] = {-9'd46,10'd354};
ram[34553] = {-9'd43,10'd358};
ram[34554] = {-9'd40,10'd361};
ram[34555] = {-9'd37,10'd364};
ram[34556] = {-9'd33,10'd367};
ram[34557] = {-9'd30,10'd370};
ram[34558] = {-9'd27,10'd373};
ram[34559] = {-9'd24,10'd376};
ram[34560] = {-9'd24,10'd376};
ram[34561] = {-9'd21,10'd380};
ram[34562] = {-9'd18,10'd383};
ram[34563] = {-9'd15,10'd386};
ram[34564] = {-9'd11,10'd389};
ram[34565] = {-9'd8,10'd392};
ram[34566] = {-9'd5,10'd395};
ram[34567] = {-9'd2,10'd398};
ram[34568] = {9'd1,-10'd399};
ram[34569] = {9'd4,-10'd396};
ram[34570] = {9'd7,-10'd393};
ram[34571] = {9'd10,-10'd390};
ram[34572] = {9'd14,-10'd387};
ram[34573] = {9'd17,-10'd384};
ram[34574] = {9'd20,-10'd381};
ram[34575] = {9'd23,-10'd377};
ram[34576] = {9'd26,-10'd374};
ram[34577] = {9'd29,-10'd371};
ram[34578] = {9'd32,-10'd368};
ram[34579] = {9'd36,-10'd365};
ram[34580] = {9'd39,-10'd362};
ram[34581] = {9'd42,-10'd359};
ram[34582] = {9'd45,-10'd355};
ram[34583] = {9'd48,-10'd352};
ram[34584] = {9'd51,-10'd349};
ram[34585] = {9'd54,-10'd346};
ram[34586] = {9'd58,-10'd343};
ram[34587] = {9'd61,-10'd340};
ram[34588] = {9'd64,-10'd337};
ram[34589] = {9'd67,-10'd334};
ram[34590] = {9'd70,-10'd330};
ram[34591] = {9'd73,-10'd327};
ram[34592] = {9'd76,-10'd324};
ram[34593] = {9'd80,-10'd321};
ram[34594] = {9'd83,-10'd318};
ram[34595] = {9'd86,-10'd315};
ram[34596] = {9'd89,-10'd312};
ram[34597] = {9'd92,-10'd308};
ram[34598] = {9'd95,-10'd305};
ram[34599] = {9'd98,-10'd302};
ram[34600] = {-9'd99,-10'd299};
ram[34601] = {-9'd96,-10'd296};
ram[34602] = {-9'd92,-10'd293};
ram[34603] = {-9'd89,-10'd290};
ram[34604] = {-9'd86,-10'd286};
ram[34605] = {-9'd83,-10'd283};
ram[34606] = {-9'd80,-10'd280};
ram[34607] = {-9'd77,-10'd277};
ram[34608] = {-9'd74,-10'd274};
ram[34609] = {-9'd70,-10'd271};
ram[34610] = {-9'd67,-10'd268};
ram[34611] = {-9'd64,-10'd264};
ram[34612] = {-9'd61,-10'd261};
ram[34613] = {-9'd58,-10'd258};
ram[34614] = {-9'd55,-10'd255};
ram[34615] = {-9'd52,-10'd252};
ram[34616] = {-9'd48,-10'd249};
ram[34617] = {-9'd45,-10'd246};
ram[34618] = {-9'd42,-10'd242};
ram[34619] = {-9'd39,-10'd239};
ram[34620] = {-9'd36,-10'd236};
ram[34621] = {-9'd33,-10'd233};
ram[34622] = {-9'd30,-10'd230};
ram[34623] = {-9'd26,-10'd227};
ram[34624] = {-9'd23,-10'd224};
ram[34625] = {-9'd20,-10'd220};
ram[34626] = {-9'd17,-10'd217};
ram[34627] = {-9'd14,-10'd214};
ram[34628] = {-9'd11,-10'd211};
ram[34629] = {-9'd8,-10'd208};
ram[34630] = {-9'd4,-10'd205};
ram[34631] = {-9'd1,-10'd202};
ram[34632] = {9'd2,-10'd198};
ram[34633] = {9'd5,-10'd195};
ram[34634] = {9'd8,-10'd192};
ram[34635] = {9'd11,-10'd189};
ram[34636] = {9'd14,-10'd186};
ram[34637] = {9'd18,-10'd183};
ram[34638] = {9'd21,-10'd180};
ram[34639] = {9'd24,-10'd176};
ram[34640] = {9'd27,-10'd173};
ram[34641] = {9'd30,-10'd170};
ram[34642] = {9'd33,-10'd167};
ram[34643] = {9'd36,-10'd164};
ram[34644] = {9'd40,-10'd161};
ram[34645] = {9'd43,-10'd158};
ram[34646] = {9'd46,-10'd154};
ram[34647] = {9'd49,-10'd151};
ram[34648] = {9'd52,-10'd148};
ram[34649] = {9'd55,-10'd145};
ram[34650] = {9'd58,-10'd142};
ram[34651] = {9'd62,-10'd139};
ram[34652] = {9'd65,-10'd136};
ram[34653] = {9'd68,-10'd132};
ram[34654] = {9'd71,-10'd129};
ram[34655] = {9'd74,-10'd126};
ram[34656] = {9'd77,-10'd123};
ram[34657] = {9'd80,-10'd120};
ram[34658] = {9'd84,-10'd117};
ram[34659] = {9'd87,-10'd114};
ram[34660] = {9'd90,-10'd110};
ram[34661] = {9'd93,-10'd107};
ram[34662] = {9'd96,-10'd104};
ram[34663] = {9'd99,-10'd101};
ram[34664] = {-9'd98,-10'd98};
ram[34665] = {-9'd95,-10'd95};
ram[34666] = {-9'd92,-10'd92};
ram[34667] = {-9'd88,-10'd88};
ram[34668] = {-9'd85,-10'd85};
ram[34669] = {-9'd82,-10'd82};
ram[34670] = {-9'd79,-10'd79};
ram[34671] = {-9'd76,-10'd76};
ram[34672] = {-9'd73,-10'd73};
ram[34673] = {-9'd70,-10'd70};
ram[34674] = {-9'd66,-10'd66};
ram[34675] = {-9'd63,-10'd63};
ram[34676] = {-9'd60,-10'd60};
ram[34677] = {-9'd57,-10'd57};
ram[34678] = {-9'd54,-10'd54};
ram[34679] = {-9'd51,-10'd51};
ram[34680] = {-9'd48,-10'd48};
ram[34681] = {-9'd44,-10'd44};
ram[34682] = {-9'd41,-10'd41};
ram[34683] = {-9'd38,-10'd38};
ram[34684] = {-9'd35,-10'd35};
ram[34685] = {-9'd32,-10'd32};
ram[34686] = {-9'd29,-10'd29};
ram[34687] = {-9'd26,-10'd26};
ram[34688] = {-9'd26,-10'd26};
ram[34689] = {-9'd22,-10'd22};
ram[34690] = {-9'd19,-10'd19};
ram[34691] = {-9'd16,-10'd16};
ram[34692] = {-9'd13,-10'd13};
ram[34693] = {-9'd10,-10'd10};
ram[34694] = {-9'd7,-10'd7};
ram[34695] = {-9'd4,-10'd4};
ram[34696] = {9'd0,10'd0};
ram[34697] = {9'd3,10'd3};
ram[34698] = {9'd6,10'd6};
ram[34699] = {9'd9,10'd9};
ram[34700] = {9'd12,10'd12};
ram[34701] = {9'd15,10'd15};
ram[34702] = {9'd18,10'd18};
ram[34703] = {9'd21,10'd21};
ram[34704] = {9'd25,10'd25};
ram[34705] = {9'd28,10'd28};
ram[34706] = {9'd31,10'd31};
ram[34707] = {9'd34,10'd34};
ram[34708] = {9'd37,10'd37};
ram[34709] = {9'd40,10'd40};
ram[34710] = {9'd43,10'd43};
ram[34711] = {9'd47,10'd47};
ram[34712] = {9'd50,10'd50};
ram[34713] = {9'd53,10'd53};
ram[34714] = {9'd56,10'd56};
ram[34715] = {9'd59,10'd59};
ram[34716] = {9'd62,10'd62};
ram[34717] = {9'd65,10'd65};
ram[34718] = {9'd69,10'd69};
ram[34719] = {9'd72,10'd72};
ram[34720] = {9'd75,10'd75};
ram[34721] = {9'd78,10'd78};
ram[34722] = {9'd81,10'd81};
ram[34723] = {9'd84,10'd84};
ram[34724] = {9'd87,10'd87};
ram[34725] = {9'd91,10'd91};
ram[34726] = {9'd94,10'd94};
ram[34727] = {9'd97,10'd97};
ram[34728] = {-9'd100,10'd100};
ram[34729] = {-9'd97,10'd103};
ram[34730] = {-9'd94,10'd106};
ram[34731] = {-9'd91,10'd109};
ram[34732] = {-9'd88,10'd113};
ram[34733] = {-9'd85,10'd116};
ram[34734] = {-9'd81,10'd119};
ram[34735] = {-9'd78,10'd122};
ram[34736] = {-9'd75,10'd125};
ram[34737] = {-9'd72,10'd128};
ram[34738] = {-9'd69,10'd131};
ram[34739] = {-9'd66,10'd135};
ram[34740] = {-9'd63,10'd138};
ram[34741] = {-9'd59,10'd141};
ram[34742] = {-9'd56,10'd144};
ram[34743] = {-9'd53,10'd147};
ram[34744] = {-9'd50,10'd150};
ram[34745] = {-9'd47,10'd153};
ram[34746] = {-9'd44,10'd157};
ram[34747] = {-9'd41,10'd160};
ram[34748] = {-9'd37,10'd163};
ram[34749] = {-9'd34,10'd166};
ram[34750] = {-9'd31,10'd169};
ram[34751] = {-9'd28,10'd172};
ram[34752] = {-9'd25,10'd175};
ram[34753] = {-9'd22,10'd179};
ram[34754] = {-9'd19,10'd182};
ram[34755] = {-9'd15,10'd185};
ram[34756] = {-9'd12,10'd188};
ram[34757] = {-9'd9,10'd191};
ram[34758] = {-9'd6,10'd194};
ram[34759] = {-9'd3,10'd197};
ram[34760] = {9'd0,10'd201};
ram[34761] = {9'd3,10'd204};
ram[34762] = {9'd7,10'd207};
ram[34763] = {9'd10,10'd210};
ram[34764] = {9'd13,10'd213};
ram[34765] = {9'd16,10'd216};
ram[34766] = {9'd19,10'd219};
ram[34767] = {9'd22,10'd223};
ram[34768] = {9'd25,10'd226};
ram[34769] = {9'd29,10'd229};
ram[34770] = {9'd32,10'd232};
ram[34771] = {9'd35,10'd235};
ram[34772] = {9'd38,10'd238};
ram[34773] = {9'd41,10'd241};
ram[34774] = {9'd44,10'd245};
ram[34775] = {9'd47,10'd248};
ram[34776] = {9'd51,10'd251};
ram[34777] = {9'd54,10'd254};
ram[34778] = {9'd57,10'd257};
ram[34779] = {9'd60,10'd260};
ram[34780] = {9'd63,10'd263};
ram[34781] = {9'd66,10'd267};
ram[34782] = {9'd69,10'd270};
ram[34783] = {9'd73,10'd273};
ram[34784] = {9'd76,10'd276};
ram[34785] = {9'd79,10'd279};
ram[34786] = {9'd82,10'd282};
ram[34787] = {9'd85,10'd285};
ram[34788] = {9'd88,10'd289};
ram[34789] = {9'd91,10'd292};
ram[34790] = {9'd95,10'd295};
ram[34791] = {9'd98,10'd298};
ram[34792] = {-9'd99,10'd301};
ram[34793] = {-9'd96,10'd304};
ram[34794] = {-9'd93,10'd307};
ram[34795] = {-9'd90,10'd311};
ram[34796] = {-9'd87,10'd314};
ram[34797] = {-9'd84,10'd317};
ram[34798] = {-9'd81,10'd320};
ram[34799] = {-9'd77,10'd323};
ram[34800] = {-9'd74,10'd326};
ram[34801] = {-9'd71,10'd329};
ram[34802] = {-9'd68,10'd333};
ram[34803] = {-9'd65,10'd336};
ram[34804] = {-9'd62,10'd339};
ram[34805] = {-9'd59,10'd342};
ram[34806] = {-9'd55,10'd345};
ram[34807] = {-9'd52,10'd348};
ram[34808] = {-9'd49,10'd351};
ram[34809] = {-9'd46,10'd354};
ram[34810] = {-9'd43,10'd358};
ram[34811] = {-9'd40,10'd361};
ram[34812] = {-9'd37,10'd364};
ram[34813] = {-9'd33,10'd367};
ram[34814] = {-9'd30,10'd370};
ram[34815] = {-9'd27,10'd373};
ram[34816] = {-9'd27,10'd373};
ram[34817] = {-9'd24,10'd376};
ram[34818] = {-9'd21,10'd380};
ram[34819] = {-9'd18,10'd383};
ram[34820] = {-9'd15,10'd386};
ram[34821] = {-9'd11,10'd389};
ram[34822] = {-9'd8,10'd392};
ram[34823] = {-9'd5,10'd395};
ram[34824] = {-9'd2,10'd398};
ram[34825] = {9'd1,-10'd399};
ram[34826] = {9'd4,-10'd396};
ram[34827] = {9'd7,-10'd393};
ram[34828] = {9'd10,-10'd390};
ram[34829] = {9'd14,-10'd387};
ram[34830] = {9'd17,-10'd384};
ram[34831] = {9'd20,-10'd381};
ram[34832] = {9'd23,-10'd377};
ram[34833] = {9'd26,-10'd374};
ram[34834] = {9'd29,-10'd371};
ram[34835] = {9'd32,-10'd368};
ram[34836] = {9'd36,-10'd365};
ram[34837] = {9'd39,-10'd362};
ram[34838] = {9'd42,-10'd359};
ram[34839] = {9'd45,-10'd355};
ram[34840] = {9'd48,-10'd352};
ram[34841] = {9'd51,-10'd349};
ram[34842] = {9'd54,-10'd346};
ram[34843] = {9'd58,-10'd343};
ram[34844] = {9'd61,-10'd340};
ram[34845] = {9'd64,-10'd337};
ram[34846] = {9'd67,-10'd334};
ram[34847] = {9'd70,-10'd330};
ram[34848] = {9'd73,-10'd327};
ram[34849] = {9'd76,-10'd324};
ram[34850] = {9'd80,-10'd321};
ram[34851] = {9'd83,-10'd318};
ram[34852] = {9'd86,-10'd315};
ram[34853] = {9'd89,-10'd312};
ram[34854] = {9'd92,-10'd308};
ram[34855] = {9'd95,-10'd305};
ram[34856] = {9'd98,-10'd302};
ram[34857] = {-9'd99,-10'd299};
ram[34858] = {-9'd96,-10'd296};
ram[34859] = {-9'd92,-10'd293};
ram[34860] = {-9'd89,-10'd290};
ram[34861] = {-9'd86,-10'd286};
ram[34862] = {-9'd83,-10'd283};
ram[34863] = {-9'd80,-10'd280};
ram[34864] = {-9'd77,-10'd277};
ram[34865] = {-9'd74,-10'd274};
ram[34866] = {-9'd70,-10'd271};
ram[34867] = {-9'd67,-10'd268};
ram[34868] = {-9'd64,-10'd264};
ram[34869] = {-9'd61,-10'd261};
ram[34870] = {-9'd58,-10'd258};
ram[34871] = {-9'd55,-10'd255};
ram[34872] = {-9'd52,-10'd252};
ram[34873] = {-9'd48,-10'd249};
ram[34874] = {-9'd45,-10'd246};
ram[34875] = {-9'd42,-10'd242};
ram[34876] = {-9'd39,-10'd239};
ram[34877] = {-9'd36,-10'd236};
ram[34878] = {-9'd33,-10'd233};
ram[34879] = {-9'd30,-10'd230};
ram[34880] = {-9'd26,-10'd227};
ram[34881] = {-9'd23,-10'd224};
ram[34882] = {-9'd20,-10'd220};
ram[34883] = {-9'd17,-10'd217};
ram[34884] = {-9'd14,-10'd214};
ram[34885] = {-9'd11,-10'd211};
ram[34886] = {-9'd8,-10'd208};
ram[34887] = {-9'd4,-10'd205};
ram[34888] = {-9'd1,-10'd202};
ram[34889] = {9'd2,-10'd198};
ram[34890] = {9'd5,-10'd195};
ram[34891] = {9'd8,-10'd192};
ram[34892] = {9'd11,-10'd189};
ram[34893] = {9'd14,-10'd186};
ram[34894] = {9'd18,-10'd183};
ram[34895] = {9'd21,-10'd180};
ram[34896] = {9'd24,-10'd176};
ram[34897] = {9'd27,-10'd173};
ram[34898] = {9'd30,-10'd170};
ram[34899] = {9'd33,-10'd167};
ram[34900] = {9'd36,-10'd164};
ram[34901] = {9'd40,-10'd161};
ram[34902] = {9'd43,-10'd158};
ram[34903] = {9'd46,-10'd154};
ram[34904] = {9'd49,-10'd151};
ram[34905] = {9'd52,-10'd148};
ram[34906] = {9'd55,-10'd145};
ram[34907] = {9'd58,-10'd142};
ram[34908] = {9'd62,-10'd139};
ram[34909] = {9'd65,-10'd136};
ram[34910] = {9'd68,-10'd132};
ram[34911] = {9'd71,-10'd129};
ram[34912] = {9'd74,-10'd126};
ram[34913] = {9'd77,-10'd123};
ram[34914] = {9'd80,-10'd120};
ram[34915] = {9'd84,-10'd117};
ram[34916] = {9'd87,-10'd114};
ram[34917] = {9'd90,-10'd110};
ram[34918] = {9'd93,-10'd107};
ram[34919] = {9'd96,-10'd104};
ram[34920] = {9'd99,-10'd101};
ram[34921] = {-9'd98,-10'd98};
ram[34922] = {-9'd95,-10'd95};
ram[34923] = {-9'd92,-10'd92};
ram[34924] = {-9'd88,-10'd88};
ram[34925] = {-9'd85,-10'd85};
ram[34926] = {-9'd82,-10'd82};
ram[34927] = {-9'd79,-10'd79};
ram[34928] = {-9'd76,-10'd76};
ram[34929] = {-9'd73,-10'd73};
ram[34930] = {-9'd70,-10'd70};
ram[34931] = {-9'd66,-10'd66};
ram[34932] = {-9'd63,-10'd63};
ram[34933] = {-9'd60,-10'd60};
ram[34934] = {-9'd57,-10'd57};
ram[34935] = {-9'd54,-10'd54};
ram[34936] = {-9'd51,-10'd51};
ram[34937] = {-9'd48,-10'd48};
ram[34938] = {-9'd44,-10'd44};
ram[34939] = {-9'd41,-10'd41};
ram[34940] = {-9'd38,-10'd38};
ram[34941] = {-9'd35,-10'd35};
ram[34942] = {-9'd32,-10'd32};
ram[34943] = {-9'd29,-10'd29};
ram[34944] = {-9'd29,-10'd29};
ram[34945] = {-9'd26,-10'd26};
ram[34946] = {-9'd22,-10'd22};
ram[34947] = {-9'd19,-10'd19};
ram[34948] = {-9'd16,-10'd16};
ram[34949] = {-9'd13,-10'd13};
ram[34950] = {-9'd10,-10'd10};
ram[34951] = {-9'd7,-10'd7};
ram[34952] = {-9'd4,-10'd4};
ram[34953] = {9'd0,10'd0};
ram[34954] = {9'd3,10'd3};
ram[34955] = {9'd6,10'd6};
ram[34956] = {9'd9,10'd9};
ram[34957] = {9'd12,10'd12};
ram[34958] = {9'd15,10'd15};
ram[34959] = {9'd18,10'd18};
ram[34960] = {9'd21,10'd21};
ram[34961] = {9'd25,10'd25};
ram[34962] = {9'd28,10'd28};
ram[34963] = {9'd31,10'd31};
ram[34964] = {9'd34,10'd34};
ram[34965] = {9'd37,10'd37};
ram[34966] = {9'd40,10'd40};
ram[34967] = {9'd43,10'd43};
ram[34968] = {9'd47,10'd47};
ram[34969] = {9'd50,10'd50};
ram[34970] = {9'd53,10'd53};
ram[34971] = {9'd56,10'd56};
ram[34972] = {9'd59,10'd59};
ram[34973] = {9'd62,10'd62};
ram[34974] = {9'd65,10'd65};
ram[34975] = {9'd69,10'd69};
ram[34976] = {9'd72,10'd72};
ram[34977] = {9'd75,10'd75};
ram[34978] = {9'd78,10'd78};
ram[34979] = {9'd81,10'd81};
ram[34980] = {9'd84,10'd84};
ram[34981] = {9'd87,10'd87};
ram[34982] = {9'd91,10'd91};
ram[34983] = {9'd94,10'd94};
ram[34984] = {9'd97,10'd97};
ram[34985] = {-9'd100,10'd100};
ram[34986] = {-9'd97,10'd103};
ram[34987] = {-9'd94,10'd106};
ram[34988] = {-9'd91,10'd109};
ram[34989] = {-9'd88,10'd113};
ram[34990] = {-9'd85,10'd116};
ram[34991] = {-9'd81,10'd119};
ram[34992] = {-9'd78,10'd122};
ram[34993] = {-9'd75,10'd125};
ram[34994] = {-9'd72,10'd128};
ram[34995] = {-9'd69,10'd131};
ram[34996] = {-9'd66,10'd135};
ram[34997] = {-9'd63,10'd138};
ram[34998] = {-9'd59,10'd141};
ram[34999] = {-9'd56,10'd144};
ram[35000] = {-9'd53,10'd147};
ram[35001] = {-9'd50,10'd150};
ram[35002] = {-9'd47,10'd153};
ram[35003] = {-9'd44,10'd157};
ram[35004] = {-9'd41,10'd160};
ram[35005] = {-9'd37,10'd163};
ram[35006] = {-9'd34,10'd166};
ram[35007] = {-9'd31,10'd169};
ram[35008] = {-9'd28,10'd172};
ram[35009] = {-9'd25,10'd175};
ram[35010] = {-9'd22,10'd179};
ram[35011] = {-9'd19,10'd182};
ram[35012] = {-9'd15,10'd185};
ram[35013] = {-9'd12,10'd188};
ram[35014] = {-9'd9,10'd191};
ram[35015] = {-9'd6,10'd194};
ram[35016] = {-9'd3,10'd197};
ram[35017] = {9'd0,10'd201};
ram[35018] = {9'd3,10'd204};
ram[35019] = {9'd7,10'd207};
ram[35020] = {9'd10,10'd210};
ram[35021] = {9'd13,10'd213};
ram[35022] = {9'd16,10'd216};
ram[35023] = {9'd19,10'd219};
ram[35024] = {9'd22,10'd223};
ram[35025] = {9'd25,10'd226};
ram[35026] = {9'd29,10'd229};
ram[35027] = {9'd32,10'd232};
ram[35028] = {9'd35,10'd235};
ram[35029] = {9'd38,10'd238};
ram[35030] = {9'd41,10'd241};
ram[35031] = {9'd44,10'd245};
ram[35032] = {9'd47,10'd248};
ram[35033] = {9'd51,10'd251};
ram[35034] = {9'd54,10'd254};
ram[35035] = {9'd57,10'd257};
ram[35036] = {9'd60,10'd260};
ram[35037] = {9'd63,10'd263};
ram[35038] = {9'd66,10'd267};
ram[35039] = {9'd69,10'd270};
ram[35040] = {9'd73,10'd273};
ram[35041] = {9'd76,10'd276};
ram[35042] = {9'd79,10'd279};
ram[35043] = {9'd82,10'd282};
ram[35044] = {9'd85,10'd285};
ram[35045] = {9'd88,10'd289};
ram[35046] = {9'd91,10'd292};
ram[35047] = {9'd95,10'd295};
ram[35048] = {9'd98,10'd298};
ram[35049] = {-9'd99,10'd301};
ram[35050] = {-9'd96,10'd304};
ram[35051] = {-9'd93,10'd307};
ram[35052] = {-9'd90,10'd311};
ram[35053] = {-9'd87,10'd314};
ram[35054] = {-9'd84,10'd317};
ram[35055] = {-9'd81,10'd320};
ram[35056] = {-9'd77,10'd323};
ram[35057] = {-9'd74,10'd326};
ram[35058] = {-9'd71,10'd329};
ram[35059] = {-9'd68,10'd333};
ram[35060] = {-9'd65,10'd336};
ram[35061] = {-9'd62,10'd339};
ram[35062] = {-9'd59,10'd342};
ram[35063] = {-9'd55,10'd345};
ram[35064] = {-9'd52,10'd348};
ram[35065] = {-9'd49,10'd351};
ram[35066] = {-9'd46,10'd354};
ram[35067] = {-9'd43,10'd358};
ram[35068] = {-9'd40,10'd361};
ram[35069] = {-9'd37,10'd364};
ram[35070] = {-9'd33,10'd367};
ram[35071] = {-9'd30,10'd370};
ram[35072] = {-9'd30,10'd370};
ram[35073] = {-9'd27,10'd373};
ram[35074] = {-9'd24,10'd376};
ram[35075] = {-9'd21,10'd380};
ram[35076] = {-9'd18,10'd383};
ram[35077] = {-9'd15,10'd386};
ram[35078] = {-9'd11,10'd389};
ram[35079] = {-9'd8,10'd392};
ram[35080] = {-9'd5,10'd395};
ram[35081] = {-9'd2,10'd398};
ram[35082] = {9'd1,-10'd399};
ram[35083] = {9'd4,-10'd396};
ram[35084] = {9'd7,-10'd393};
ram[35085] = {9'd10,-10'd390};
ram[35086] = {9'd14,-10'd387};
ram[35087] = {9'd17,-10'd384};
ram[35088] = {9'd20,-10'd381};
ram[35089] = {9'd23,-10'd377};
ram[35090] = {9'd26,-10'd374};
ram[35091] = {9'd29,-10'd371};
ram[35092] = {9'd32,-10'd368};
ram[35093] = {9'd36,-10'd365};
ram[35094] = {9'd39,-10'd362};
ram[35095] = {9'd42,-10'd359};
ram[35096] = {9'd45,-10'd355};
ram[35097] = {9'd48,-10'd352};
ram[35098] = {9'd51,-10'd349};
ram[35099] = {9'd54,-10'd346};
ram[35100] = {9'd58,-10'd343};
ram[35101] = {9'd61,-10'd340};
ram[35102] = {9'd64,-10'd337};
ram[35103] = {9'd67,-10'd334};
ram[35104] = {9'd70,-10'd330};
ram[35105] = {9'd73,-10'd327};
ram[35106] = {9'd76,-10'd324};
ram[35107] = {9'd80,-10'd321};
ram[35108] = {9'd83,-10'd318};
ram[35109] = {9'd86,-10'd315};
ram[35110] = {9'd89,-10'd312};
ram[35111] = {9'd92,-10'd308};
ram[35112] = {9'd95,-10'd305};
ram[35113] = {9'd98,-10'd302};
ram[35114] = {-9'd99,-10'd299};
ram[35115] = {-9'd96,-10'd296};
ram[35116] = {-9'd92,-10'd293};
ram[35117] = {-9'd89,-10'd290};
ram[35118] = {-9'd86,-10'd286};
ram[35119] = {-9'd83,-10'd283};
ram[35120] = {-9'd80,-10'd280};
ram[35121] = {-9'd77,-10'd277};
ram[35122] = {-9'd74,-10'd274};
ram[35123] = {-9'd70,-10'd271};
ram[35124] = {-9'd67,-10'd268};
ram[35125] = {-9'd64,-10'd264};
ram[35126] = {-9'd61,-10'd261};
ram[35127] = {-9'd58,-10'd258};
ram[35128] = {-9'd55,-10'd255};
ram[35129] = {-9'd52,-10'd252};
ram[35130] = {-9'd48,-10'd249};
ram[35131] = {-9'd45,-10'd246};
ram[35132] = {-9'd42,-10'd242};
ram[35133] = {-9'd39,-10'd239};
ram[35134] = {-9'd36,-10'd236};
ram[35135] = {-9'd33,-10'd233};
ram[35136] = {-9'd30,-10'd230};
ram[35137] = {-9'd26,-10'd227};
ram[35138] = {-9'd23,-10'd224};
ram[35139] = {-9'd20,-10'd220};
ram[35140] = {-9'd17,-10'd217};
ram[35141] = {-9'd14,-10'd214};
ram[35142] = {-9'd11,-10'd211};
ram[35143] = {-9'd8,-10'd208};
ram[35144] = {-9'd4,-10'd205};
ram[35145] = {-9'd1,-10'd202};
ram[35146] = {9'd2,-10'd198};
ram[35147] = {9'd5,-10'd195};
ram[35148] = {9'd8,-10'd192};
ram[35149] = {9'd11,-10'd189};
ram[35150] = {9'd14,-10'd186};
ram[35151] = {9'd18,-10'd183};
ram[35152] = {9'd21,-10'd180};
ram[35153] = {9'd24,-10'd176};
ram[35154] = {9'd27,-10'd173};
ram[35155] = {9'd30,-10'd170};
ram[35156] = {9'd33,-10'd167};
ram[35157] = {9'd36,-10'd164};
ram[35158] = {9'd40,-10'd161};
ram[35159] = {9'd43,-10'd158};
ram[35160] = {9'd46,-10'd154};
ram[35161] = {9'd49,-10'd151};
ram[35162] = {9'd52,-10'd148};
ram[35163] = {9'd55,-10'd145};
ram[35164] = {9'd58,-10'd142};
ram[35165] = {9'd62,-10'd139};
ram[35166] = {9'd65,-10'd136};
ram[35167] = {9'd68,-10'd132};
ram[35168] = {9'd71,-10'd129};
ram[35169] = {9'd74,-10'd126};
ram[35170] = {9'd77,-10'd123};
ram[35171] = {9'd80,-10'd120};
ram[35172] = {9'd84,-10'd117};
ram[35173] = {9'd87,-10'd114};
ram[35174] = {9'd90,-10'd110};
ram[35175] = {9'd93,-10'd107};
ram[35176] = {9'd96,-10'd104};
ram[35177] = {9'd99,-10'd101};
ram[35178] = {-9'd98,-10'd98};
ram[35179] = {-9'd95,-10'd95};
ram[35180] = {-9'd92,-10'd92};
ram[35181] = {-9'd88,-10'd88};
ram[35182] = {-9'd85,-10'd85};
ram[35183] = {-9'd82,-10'd82};
ram[35184] = {-9'd79,-10'd79};
ram[35185] = {-9'd76,-10'd76};
ram[35186] = {-9'd73,-10'd73};
ram[35187] = {-9'd70,-10'd70};
ram[35188] = {-9'd66,-10'd66};
ram[35189] = {-9'd63,-10'd63};
ram[35190] = {-9'd60,-10'd60};
ram[35191] = {-9'd57,-10'd57};
ram[35192] = {-9'd54,-10'd54};
ram[35193] = {-9'd51,-10'd51};
ram[35194] = {-9'd48,-10'd48};
ram[35195] = {-9'd44,-10'd44};
ram[35196] = {-9'd41,-10'd41};
ram[35197] = {-9'd38,-10'd38};
ram[35198] = {-9'd35,-10'd35};
ram[35199] = {-9'd32,-10'd32};
ram[35200] = {-9'd32,-10'd32};
ram[35201] = {-9'd29,-10'd29};
ram[35202] = {-9'd26,-10'd26};
ram[35203] = {-9'd22,-10'd22};
ram[35204] = {-9'd19,-10'd19};
ram[35205] = {-9'd16,-10'd16};
ram[35206] = {-9'd13,-10'd13};
ram[35207] = {-9'd10,-10'd10};
ram[35208] = {-9'd7,-10'd7};
ram[35209] = {-9'd4,-10'd4};
ram[35210] = {9'd0,10'd0};
ram[35211] = {9'd3,10'd3};
ram[35212] = {9'd6,10'd6};
ram[35213] = {9'd9,10'd9};
ram[35214] = {9'd12,10'd12};
ram[35215] = {9'd15,10'd15};
ram[35216] = {9'd18,10'd18};
ram[35217] = {9'd21,10'd21};
ram[35218] = {9'd25,10'd25};
ram[35219] = {9'd28,10'd28};
ram[35220] = {9'd31,10'd31};
ram[35221] = {9'd34,10'd34};
ram[35222] = {9'd37,10'd37};
ram[35223] = {9'd40,10'd40};
ram[35224] = {9'd43,10'd43};
ram[35225] = {9'd47,10'd47};
ram[35226] = {9'd50,10'd50};
ram[35227] = {9'd53,10'd53};
ram[35228] = {9'd56,10'd56};
ram[35229] = {9'd59,10'd59};
ram[35230] = {9'd62,10'd62};
ram[35231] = {9'd65,10'd65};
ram[35232] = {9'd69,10'd69};
ram[35233] = {9'd72,10'd72};
ram[35234] = {9'd75,10'd75};
ram[35235] = {9'd78,10'd78};
ram[35236] = {9'd81,10'd81};
ram[35237] = {9'd84,10'd84};
ram[35238] = {9'd87,10'd87};
ram[35239] = {9'd91,10'd91};
ram[35240] = {9'd94,10'd94};
ram[35241] = {9'd97,10'd97};
ram[35242] = {-9'd100,10'd100};
ram[35243] = {-9'd97,10'd103};
ram[35244] = {-9'd94,10'd106};
ram[35245] = {-9'd91,10'd109};
ram[35246] = {-9'd88,10'd113};
ram[35247] = {-9'd85,10'd116};
ram[35248] = {-9'd81,10'd119};
ram[35249] = {-9'd78,10'd122};
ram[35250] = {-9'd75,10'd125};
ram[35251] = {-9'd72,10'd128};
ram[35252] = {-9'd69,10'd131};
ram[35253] = {-9'd66,10'd135};
ram[35254] = {-9'd63,10'd138};
ram[35255] = {-9'd59,10'd141};
ram[35256] = {-9'd56,10'd144};
ram[35257] = {-9'd53,10'd147};
ram[35258] = {-9'd50,10'd150};
ram[35259] = {-9'd47,10'd153};
ram[35260] = {-9'd44,10'd157};
ram[35261] = {-9'd41,10'd160};
ram[35262] = {-9'd37,10'd163};
ram[35263] = {-9'd34,10'd166};
ram[35264] = {-9'd31,10'd169};
ram[35265] = {-9'd28,10'd172};
ram[35266] = {-9'd25,10'd175};
ram[35267] = {-9'd22,10'd179};
ram[35268] = {-9'd19,10'd182};
ram[35269] = {-9'd15,10'd185};
ram[35270] = {-9'd12,10'd188};
ram[35271] = {-9'd9,10'd191};
ram[35272] = {-9'd6,10'd194};
ram[35273] = {-9'd3,10'd197};
ram[35274] = {9'd0,10'd201};
ram[35275] = {9'd3,10'd204};
ram[35276] = {9'd7,10'd207};
ram[35277] = {9'd10,10'd210};
ram[35278] = {9'd13,10'd213};
ram[35279] = {9'd16,10'd216};
ram[35280] = {9'd19,10'd219};
ram[35281] = {9'd22,10'd223};
ram[35282] = {9'd25,10'd226};
ram[35283] = {9'd29,10'd229};
ram[35284] = {9'd32,10'd232};
ram[35285] = {9'd35,10'd235};
ram[35286] = {9'd38,10'd238};
ram[35287] = {9'd41,10'd241};
ram[35288] = {9'd44,10'd245};
ram[35289] = {9'd47,10'd248};
ram[35290] = {9'd51,10'd251};
ram[35291] = {9'd54,10'd254};
ram[35292] = {9'd57,10'd257};
ram[35293] = {9'd60,10'd260};
ram[35294] = {9'd63,10'd263};
ram[35295] = {9'd66,10'd267};
ram[35296] = {9'd69,10'd270};
ram[35297] = {9'd73,10'd273};
ram[35298] = {9'd76,10'd276};
ram[35299] = {9'd79,10'd279};
ram[35300] = {9'd82,10'd282};
ram[35301] = {9'd85,10'd285};
ram[35302] = {9'd88,10'd289};
ram[35303] = {9'd91,10'd292};
ram[35304] = {9'd95,10'd295};
ram[35305] = {9'd98,10'd298};
ram[35306] = {-9'd99,10'd301};
ram[35307] = {-9'd96,10'd304};
ram[35308] = {-9'd93,10'd307};
ram[35309] = {-9'd90,10'd311};
ram[35310] = {-9'd87,10'd314};
ram[35311] = {-9'd84,10'd317};
ram[35312] = {-9'd81,10'd320};
ram[35313] = {-9'd77,10'd323};
ram[35314] = {-9'd74,10'd326};
ram[35315] = {-9'd71,10'd329};
ram[35316] = {-9'd68,10'd333};
ram[35317] = {-9'd65,10'd336};
ram[35318] = {-9'd62,10'd339};
ram[35319] = {-9'd59,10'd342};
ram[35320] = {-9'd55,10'd345};
ram[35321] = {-9'd52,10'd348};
ram[35322] = {-9'd49,10'd351};
ram[35323] = {-9'd46,10'd354};
ram[35324] = {-9'd43,10'd358};
ram[35325] = {-9'd40,10'd361};
ram[35326] = {-9'd37,10'd364};
ram[35327] = {-9'd33,10'd367};
ram[35328] = {-9'd33,10'd367};
ram[35329] = {-9'd30,10'd370};
ram[35330] = {-9'd27,10'd373};
ram[35331] = {-9'd24,10'd376};
ram[35332] = {-9'd21,10'd380};
ram[35333] = {-9'd18,10'd383};
ram[35334] = {-9'd15,10'd386};
ram[35335] = {-9'd11,10'd389};
ram[35336] = {-9'd8,10'd392};
ram[35337] = {-9'd5,10'd395};
ram[35338] = {-9'd2,10'd398};
ram[35339] = {9'd1,-10'd399};
ram[35340] = {9'd4,-10'd396};
ram[35341] = {9'd7,-10'd393};
ram[35342] = {9'd10,-10'd390};
ram[35343] = {9'd14,-10'd387};
ram[35344] = {9'd17,-10'd384};
ram[35345] = {9'd20,-10'd381};
ram[35346] = {9'd23,-10'd377};
ram[35347] = {9'd26,-10'd374};
ram[35348] = {9'd29,-10'd371};
ram[35349] = {9'd32,-10'd368};
ram[35350] = {9'd36,-10'd365};
ram[35351] = {9'd39,-10'd362};
ram[35352] = {9'd42,-10'd359};
ram[35353] = {9'd45,-10'd355};
ram[35354] = {9'd48,-10'd352};
ram[35355] = {9'd51,-10'd349};
ram[35356] = {9'd54,-10'd346};
ram[35357] = {9'd58,-10'd343};
ram[35358] = {9'd61,-10'd340};
ram[35359] = {9'd64,-10'd337};
ram[35360] = {9'd67,-10'd334};
ram[35361] = {9'd70,-10'd330};
ram[35362] = {9'd73,-10'd327};
ram[35363] = {9'd76,-10'd324};
ram[35364] = {9'd80,-10'd321};
ram[35365] = {9'd83,-10'd318};
ram[35366] = {9'd86,-10'd315};
ram[35367] = {9'd89,-10'd312};
ram[35368] = {9'd92,-10'd308};
ram[35369] = {9'd95,-10'd305};
ram[35370] = {9'd98,-10'd302};
ram[35371] = {-9'd99,-10'd299};
ram[35372] = {-9'd96,-10'd296};
ram[35373] = {-9'd92,-10'd293};
ram[35374] = {-9'd89,-10'd290};
ram[35375] = {-9'd86,-10'd286};
ram[35376] = {-9'd83,-10'd283};
ram[35377] = {-9'd80,-10'd280};
ram[35378] = {-9'd77,-10'd277};
ram[35379] = {-9'd74,-10'd274};
ram[35380] = {-9'd70,-10'd271};
ram[35381] = {-9'd67,-10'd268};
ram[35382] = {-9'd64,-10'd264};
ram[35383] = {-9'd61,-10'd261};
ram[35384] = {-9'd58,-10'd258};
ram[35385] = {-9'd55,-10'd255};
ram[35386] = {-9'd52,-10'd252};
ram[35387] = {-9'd48,-10'd249};
ram[35388] = {-9'd45,-10'd246};
ram[35389] = {-9'd42,-10'd242};
ram[35390] = {-9'd39,-10'd239};
ram[35391] = {-9'd36,-10'd236};
ram[35392] = {-9'd33,-10'd233};
ram[35393] = {-9'd30,-10'd230};
ram[35394] = {-9'd26,-10'd227};
ram[35395] = {-9'd23,-10'd224};
ram[35396] = {-9'd20,-10'd220};
ram[35397] = {-9'd17,-10'd217};
ram[35398] = {-9'd14,-10'd214};
ram[35399] = {-9'd11,-10'd211};
ram[35400] = {-9'd8,-10'd208};
ram[35401] = {-9'd4,-10'd205};
ram[35402] = {-9'd1,-10'd202};
ram[35403] = {9'd2,-10'd198};
ram[35404] = {9'd5,-10'd195};
ram[35405] = {9'd8,-10'd192};
ram[35406] = {9'd11,-10'd189};
ram[35407] = {9'd14,-10'd186};
ram[35408] = {9'd18,-10'd183};
ram[35409] = {9'd21,-10'd180};
ram[35410] = {9'd24,-10'd176};
ram[35411] = {9'd27,-10'd173};
ram[35412] = {9'd30,-10'd170};
ram[35413] = {9'd33,-10'd167};
ram[35414] = {9'd36,-10'd164};
ram[35415] = {9'd40,-10'd161};
ram[35416] = {9'd43,-10'd158};
ram[35417] = {9'd46,-10'd154};
ram[35418] = {9'd49,-10'd151};
ram[35419] = {9'd52,-10'd148};
ram[35420] = {9'd55,-10'd145};
ram[35421] = {9'd58,-10'd142};
ram[35422] = {9'd62,-10'd139};
ram[35423] = {9'd65,-10'd136};
ram[35424] = {9'd68,-10'd132};
ram[35425] = {9'd71,-10'd129};
ram[35426] = {9'd74,-10'd126};
ram[35427] = {9'd77,-10'd123};
ram[35428] = {9'd80,-10'd120};
ram[35429] = {9'd84,-10'd117};
ram[35430] = {9'd87,-10'd114};
ram[35431] = {9'd90,-10'd110};
ram[35432] = {9'd93,-10'd107};
ram[35433] = {9'd96,-10'd104};
ram[35434] = {9'd99,-10'd101};
ram[35435] = {-9'd98,-10'd98};
ram[35436] = {-9'd95,-10'd95};
ram[35437] = {-9'd92,-10'd92};
ram[35438] = {-9'd88,-10'd88};
ram[35439] = {-9'd85,-10'd85};
ram[35440] = {-9'd82,-10'd82};
ram[35441] = {-9'd79,-10'd79};
ram[35442] = {-9'd76,-10'd76};
ram[35443] = {-9'd73,-10'd73};
ram[35444] = {-9'd70,-10'd70};
ram[35445] = {-9'd66,-10'd66};
ram[35446] = {-9'd63,-10'd63};
ram[35447] = {-9'd60,-10'd60};
ram[35448] = {-9'd57,-10'd57};
ram[35449] = {-9'd54,-10'd54};
ram[35450] = {-9'd51,-10'd51};
ram[35451] = {-9'd48,-10'd48};
ram[35452] = {-9'd44,-10'd44};
ram[35453] = {-9'd41,-10'd41};
ram[35454] = {-9'd38,-10'd38};
ram[35455] = {-9'd35,-10'd35};
ram[35456] = {-9'd35,-10'd35};
ram[35457] = {-9'd32,-10'd32};
ram[35458] = {-9'd29,-10'd29};
ram[35459] = {-9'd26,-10'd26};
ram[35460] = {-9'd22,-10'd22};
ram[35461] = {-9'd19,-10'd19};
ram[35462] = {-9'd16,-10'd16};
ram[35463] = {-9'd13,-10'd13};
ram[35464] = {-9'd10,-10'd10};
ram[35465] = {-9'd7,-10'd7};
ram[35466] = {-9'd4,-10'd4};
ram[35467] = {9'd0,10'd0};
ram[35468] = {9'd3,10'd3};
ram[35469] = {9'd6,10'd6};
ram[35470] = {9'd9,10'd9};
ram[35471] = {9'd12,10'd12};
ram[35472] = {9'd15,10'd15};
ram[35473] = {9'd18,10'd18};
ram[35474] = {9'd21,10'd21};
ram[35475] = {9'd25,10'd25};
ram[35476] = {9'd28,10'd28};
ram[35477] = {9'd31,10'd31};
ram[35478] = {9'd34,10'd34};
ram[35479] = {9'd37,10'd37};
ram[35480] = {9'd40,10'd40};
ram[35481] = {9'd43,10'd43};
ram[35482] = {9'd47,10'd47};
ram[35483] = {9'd50,10'd50};
ram[35484] = {9'd53,10'd53};
ram[35485] = {9'd56,10'd56};
ram[35486] = {9'd59,10'd59};
ram[35487] = {9'd62,10'd62};
ram[35488] = {9'd65,10'd65};
ram[35489] = {9'd69,10'd69};
ram[35490] = {9'd72,10'd72};
ram[35491] = {9'd75,10'd75};
ram[35492] = {9'd78,10'd78};
ram[35493] = {9'd81,10'd81};
ram[35494] = {9'd84,10'd84};
ram[35495] = {9'd87,10'd87};
ram[35496] = {9'd91,10'd91};
ram[35497] = {9'd94,10'd94};
ram[35498] = {9'd97,10'd97};
ram[35499] = {-9'd100,10'd100};
ram[35500] = {-9'd97,10'd103};
ram[35501] = {-9'd94,10'd106};
ram[35502] = {-9'd91,10'd109};
ram[35503] = {-9'd88,10'd113};
ram[35504] = {-9'd85,10'd116};
ram[35505] = {-9'd81,10'd119};
ram[35506] = {-9'd78,10'd122};
ram[35507] = {-9'd75,10'd125};
ram[35508] = {-9'd72,10'd128};
ram[35509] = {-9'd69,10'd131};
ram[35510] = {-9'd66,10'd135};
ram[35511] = {-9'd63,10'd138};
ram[35512] = {-9'd59,10'd141};
ram[35513] = {-9'd56,10'd144};
ram[35514] = {-9'd53,10'd147};
ram[35515] = {-9'd50,10'd150};
ram[35516] = {-9'd47,10'd153};
ram[35517] = {-9'd44,10'd157};
ram[35518] = {-9'd41,10'd160};
ram[35519] = {-9'd37,10'd163};
ram[35520] = {-9'd34,10'd166};
ram[35521] = {-9'd31,10'd169};
ram[35522] = {-9'd28,10'd172};
ram[35523] = {-9'd25,10'd175};
ram[35524] = {-9'd22,10'd179};
ram[35525] = {-9'd19,10'd182};
ram[35526] = {-9'd15,10'd185};
ram[35527] = {-9'd12,10'd188};
ram[35528] = {-9'd9,10'd191};
ram[35529] = {-9'd6,10'd194};
ram[35530] = {-9'd3,10'd197};
ram[35531] = {9'd0,10'd201};
ram[35532] = {9'd3,10'd204};
ram[35533] = {9'd7,10'd207};
ram[35534] = {9'd10,10'd210};
ram[35535] = {9'd13,10'd213};
ram[35536] = {9'd16,10'd216};
ram[35537] = {9'd19,10'd219};
ram[35538] = {9'd22,10'd223};
ram[35539] = {9'd25,10'd226};
ram[35540] = {9'd29,10'd229};
ram[35541] = {9'd32,10'd232};
ram[35542] = {9'd35,10'd235};
ram[35543] = {9'd38,10'd238};
ram[35544] = {9'd41,10'd241};
ram[35545] = {9'd44,10'd245};
ram[35546] = {9'd47,10'd248};
ram[35547] = {9'd51,10'd251};
ram[35548] = {9'd54,10'd254};
ram[35549] = {9'd57,10'd257};
ram[35550] = {9'd60,10'd260};
ram[35551] = {9'd63,10'd263};
ram[35552] = {9'd66,10'd267};
ram[35553] = {9'd69,10'd270};
ram[35554] = {9'd73,10'd273};
ram[35555] = {9'd76,10'd276};
ram[35556] = {9'd79,10'd279};
ram[35557] = {9'd82,10'd282};
ram[35558] = {9'd85,10'd285};
ram[35559] = {9'd88,10'd289};
ram[35560] = {9'd91,10'd292};
ram[35561] = {9'd95,10'd295};
ram[35562] = {9'd98,10'd298};
ram[35563] = {-9'd99,10'd301};
ram[35564] = {-9'd96,10'd304};
ram[35565] = {-9'd93,10'd307};
ram[35566] = {-9'd90,10'd311};
ram[35567] = {-9'd87,10'd314};
ram[35568] = {-9'd84,10'd317};
ram[35569] = {-9'd81,10'd320};
ram[35570] = {-9'd77,10'd323};
ram[35571] = {-9'd74,10'd326};
ram[35572] = {-9'd71,10'd329};
ram[35573] = {-9'd68,10'd333};
ram[35574] = {-9'd65,10'd336};
ram[35575] = {-9'd62,10'd339};
ram[35576] = {-9'd59,10'd342};
ram[35577] = {-9'd55,10'd345};
ram[35578] = {-9'd52,10'd348};
ram[35579] = {-9'd49,10'd351};
ram[35580] = {-9'd46,10'd354};
ram[35581] = {-9'd43,10'd358};
ram[35582] = {-9'd40,10'd361};
ram[35583] = {-9'd37,10'd364};
ram[35584] = {-9'd37,10'd364};
ram[35585] = {-9'd33,10'd367};
ram[35586] = {-9'd30,10'd370};
ram[35587] = {-9'd27,10'd373};
ram[35588] = {-9'd24,10'd376};
ram[35589] = {-9'd21,10'd380};
ram[35590] = {-9'd18,10'd383};
ram[35591] = {-9'd15,10'd386};
ram[35592] = {-9'd11,10'd389};
ram[35593] = {-9'd8,10'd392};
ram[35594] = {-9'd5,10'd395};
ram[35595] = {-9'd2,10'd398};
ram[35596] = {9'd1,-10'd399};
ram[35597] = {9'd4,-10'd396};
ram[35598] = {9'd7,-10'd393};
ram[35599] = {9'd10,-10'd390};
ram[35600] = {9'd14,-10'd387};
ram[35601] = {9'd17,-10'd384};
ram[35602] = {9'd20,-10'd381};
ram[35603] = {9'd23,-10'd377};
ram[35604] = {9'd26,-10'd374};
ram[35605] = {9'd29,-10'd371};
ram[35606] = {9'd32,-10'd368};
ram[35607] = {9'd36,-10'd365};
ram[35608] = {9'd39,-10'd362};
ram[35609] = {9'd42,-10'd359};
ram[35610] = {9'd45,-10'd355};
ram[35611] = {9'd48,-10'd352};
ram[35612] = {9'd51,-10'd349};
ram[35613] = {9'd54,-10'd346};
ram[35614] = {9'd58,-10'd343};
ram[35615] = {9'd61,-10'd340};
ram[35616] = {9'd64,-10'd337};
ram[35617] = {9'd67,-10'd334};
ram[35618] = {9'd70,-10'd330};
ram[35619] = {9'd73,-10'd327};
ram[35620] = {9'd76,-10'd324};
ram[35621] = {9'd80,-10'd321};
ram[35622] = {9'd83,-10'd318};
ram[35623] = {9'd86,-10'd315};
ram[35624] = {9'd89,-10'd312};
ram[35625] = {9'd92,-10'd308};
ram[35626] = {9'd95,-10'd305};
ram[35627] = {9'd98,-10'd302};
ram[35628] = {-9'd99,-10'd299};
ram[35629] = {-9'd96,-10'd296};
ram[35630] = {-9'd92,-10'd293};
ram[35631] = {-9'd89,-10'd290};
ram[35632] = {-9'd86,-10'd286};
ram[35633] = {-9'd83,-10'd283};
ram[35634] = {-9'd80,-10'd280};
ram[35635] = {-9'd77,-10'd277};
ram[35636] = {-9'd74,-10'd274};
ram[35637] = {-9'd70,-10'd271};
ram[35638] = {-9'd67,-10'd268};
ram[35639] = {-9'd64,-10'd264};
ram[35640] = {-9'd61,-10'd261};
ram[35641] = {-9'd58,-10'd258};
ram[35642] = {-9'd55,-10'd255};
ram[35643] = {-9'd52,-10'd252};
ram[35644] = {-9'd48,-10'd249};
ram[35645] = {-9'd45,-10'd246};
ram[35646] = {-9'd42,-10'd242};
ram[35647] = {-9'd39,-10'd239};
ram[35648] = {-9'd36,-10'd236};
ram[35649] = {-9'd33,-10'd233};
ram[35650] = {-9'd30,-10'd230};
ram[35651] = {-9'd26,-10'd227};
ram[35652] = {-9'd23,-10'd224};
ram[35653] = {-9'd20,-10'd220};
ram[35654] = {-9'd17,-10'd217};
ram[35655] = {-9'd14,-10'd214};
ram[35656] = {-9'd11,-10'd211};
ram[35657] = {-9'd8,-10'd208};
ram[35658] = {-9'd4,-10'd205};
ram[35659] = {-9'd1,-10'd202};
ram[35660] = {9'd2,-10'd198};
ram[35661] = {9'd5,-10'd195};
ram[35662] = {9'd8,-10'd192};
ram[35663] = {9'd11,-10'd189};
ram[35664] = {9'd14,-10'd186};
ram[35665] = {9'd18,-10'd183};
ram[35666] = {9'd21,-10'd180};
ram[35667] = {9'd24,-10'd176};
ram[35668] = {9'd27,-10'd173};
ram[35669] = {9'd30,-10'd170};
ram[35670] = {9'd33,-10'd167};
ram[35671] = {9'd36,-10'd164};
ram[35672] = {9'd40,-10'd161};
ram[35673] = {9'd43,-10'd158};
ram[35674] = {9'd46,-10'd154};
ram[35675] = {9'd49,-10'd151};
ram[35676] = {9'd52,-10'd148};
ram[35677] = {9'd55,-10'd145};
ram[35678] = {9'd58,-10'd142};
ram[35679] = {9'd62,-10'd139};
ram[35680] = {9'd65,-10'd136};
ram[35681] = {9'd68,-10'd132};
ram[35682] = {9'd71,-10'd129};
ram[35683] = {9'd74,-10'd126};
ram[35684] = {9'd77,-10'd123};
ram[35685] = {9'd80,-10'd120};
ram[35686] = {9'd84,-10'd117};
ram[35687] = {9'd87,-10'd114};
ram[35688] = {9'd90,-10'd110};
ram[35689] = {9'd93,-10'd107};
ram[35690] = {9'd96,-10'd104};
ram[35691] = {9'd99,-10'd101};
ram[35692] = {-9'd98,-10'd98};
ram[35693] = {-9'd95,-10'd95};
ram[35694] = {-9'd92,-10'd92};
ram[35695] = {-9'd88,-10'd88};
ram[35696] = {-9'd85,-10'd85};
ram[35697] = {-9'd82,-10'd82};
ram[35698] = {-9'd79,-10'd79};
ram[35699] = {-9'd76,-10'd76};
ram[35700] = {-9'd73,-10'd73};
ram[35701] = {-9'd70,-10'd70};
ram[35702] = {-9'd66,-10'd66};
ram[35703] = {-9'd63,-10'd63};
ram[35704] = {-9'd60,-10'd60};
ram[35705] = {-9'd57,-10'd57};
ram[35706] = {-9'd54,-10'd54};
ram[35707] = {-9'd51,-10'd51};
ram[35708] = {-9'd48,-10'd48};
ram[35709] = {-9'd44,-10'd44};
ram[35710] = {-9'd41,-10'd41};
ram[35711] = {-9'd38,-10'd38};
ram[35712] = {-9'd38,-10'd38};
ram[35713] = {-9'd35,-10'd35};
ram[35714] = {-9'd32,-10'd32};
ram[35715] = {-9'd29,-10'd29};
ram[35716] = {-9'd26,-10'd26};
ram[35717] = {-9'd22,-10'd22};
ram[35718] = {-9'd19,-10'd19};
ram[35719] = {-9'd16,-10'd16};
ram[35720] = {-9'd13,-10'd13};
ram[35721] = {-9'd10,-10'd10};
ram[35722] = {-9'd7,-10'd7};
ram[35723] = {-9'd4,-10'd4};
ram[35724] = {9'd0,10'd0};
ram[35725] = {9'd3,10'd3};
ram[35726] = {9'd6,10'd6};
ram[35727] = {9'd9,10'd9};
ram[35728] = {9'd12,10'd12};
ram[35729] = {9'd15,10'd15};
ram[35730] = {9'd18,10'd18};
ram[35731] = {9'd21,10'd21};
ram[35732] = {9'd25,10'd25};
ram[35733] = {9'd28,10'd28};
ram[35734] = {9'd31,10'd31};
ram[35735] = {9'd34,10'd34};
ram[35736] = {9'd37,10'd37};
ram[35737] = {9'd40,10'd40};
ram[35738] = {9'd43,10'd43};
ram[35739] = {9'd47,10'd47};
ram[35740] = {9'd50,10'd50};
ram[35741] = {9'd53,10'd53};
ram[35742] = {9'd56,10'd56};
ram[35743] = {9'd59,10'd59};
ram[35744] = {9'd62,10'd62};
ram[35745] = {9'd65,10'd65};
ram[35746] = {9'd69,10'd69};
ram[35747] = {9'd72,10'd72};
ram[35748] = {9'd75,10'd75};
ram[35749] = {9'd78,10'd78};
ram[35750] = {9'd81,10'd81};
ram[35751] = {9'd84,10'd84};
ram[35752] = {9'd87,10'd87};
ram[35753] = {9'd91,10'd91};
ram[35754] = {9'd94,10'd94};
ram[35755] = {9'd97,10'd97};
ram[35756] = {-9'd100,10'd100};
ram[35757] = {-9'd97,10'd103};
ram[35758] = {-9'd94,10'd106};
ram[35759] = {-9'd91,10'd109};
ram[35760] = {-9'd88,10'd113};
ram[35761] = {-9'd85,10'd116};
ram[35762] = {-9'd81,10'd119};
ram[35763] = {-9'd78,10'd122};
ram[35764] = {-9'd75,10'd125};
ram[35765] = {-9'd72,10'd128};
ram[35766] = {-9'd69,10'd131};
ram[35767] = {-9'd66,10'd135};
ram[35768] = {-9'd63,10'd138};
ram[35769] = {-9'd59,10'd141};
ram[35770] = {-9'd56,10'd144};
ram[35771] = {-9'd53,10'd147};
ram[35772] = {-9'd50,10'd150};
ram[35773] = {-9'd47,10'd153};
ram[35774] = {-9'd44,10'd157};
ram[35775] = {-9'd41,10'd160};
ram[35776] = {-9'd37,10'd163};
ram[35777] = {-9'd34,10'd166};
ram[35778] = {-9'd31,10'd169};
ram[35779] = {-9'd28,10'd172};
ram[35780] = {-9'd25,10'd175};
ram[35781] = {-9'd22,10'd179};
ram[35782] = {-9'd19,10'd182};
ram[35783] = {-9'd15,10'd185};
ram[35784] = {-9'd12,10'd188};
ram[35785] = {-9'd9,10'd191};
ram[35786] = {-9'd6,10'd194};
ram[35787] = {-9'd3,10'd197};
ram[35788] = {9'd0,10'd201};
ram[35789] = {9'd3,10'd204};
ram[35790] = {9'd7,10'd207};
ram[35791] = {9'd10,10'd210};
ram[35792] = {9'd13,10'd213};
ram[35793] = {9'd16,10'd216};
ram[35794] = {9'd19,10'd219};
ram[35795] = {9'd22,10'd223};
ram[35796] = {9'd25,10'd226};
ram[35797] = {9'd29,10'd229};
ram[35798] = {9'd32,10'd232};
ram[35799] = {9'd35,10'd235};
ram[35800] = {9'd38,10'd238};
ram[35801] = {9'd41,10'd241};
ram[35802] = {9'd44,10'd245};
ram[35803] = {9'd47,10'd248};
ram[35804] = {9'd51,10'd251};
ram[35805] = {9'd54,10'd254};
ram[35806] = {9'd57,10'd257};
ram[35807] = {9'd60,10'd260};
ram[35808] = {9'd63,10'd263};
ram[35809] = {9'd66,10'd267};
ram[35810] = {9'd69,10'd270};
ram[35811] = {9'd73,10'd273};
ram[35812] = {9'd76,10'd276};
ram[35813] = {9'd79,10'd279};
ram[35814] = {9'd82,10'd282};
ram[35815] = {9'd85,10'd285};
ram[35816] = {9'd88,10'd289};
ram[35817] = {9'd91,10'd292};
ram[35818] = {9'd95,10'd295};
ram[35819] = {9'd98,10'd298};
ram[35820] = {-9'd99,10'd301};
ram[35821] = {-9'd96,10'd304};
ram[35822] = {-9'd93,10'd307};
ram[35823] = {-9'd90,10'd311};
ram[35824] = {-9'd87,10'd314};
ram[35825] = {-9'd84,10'd317};
ram[35826] = {-9'd81,10'd320};
ram[35827] = {-9'd77,10'd323};
ram[35828] = {-9'd74,10'd326};
ram[35829] = {-9'd71,10'd329};
ram[35830] = {-9'd68,10'd333};
ram[35831] = {-9'd65,10'd336};
ram[35832] = {-9'd62,10'd339};
ram[35833] = {-9'd59,10'd342};
ram[35834] = {-9'd55,10'd345};
ram[35835] = {-9'd52,10'd348};
ram[35836] = {-9'd49,10'd351};
ram[35837] = {-9'd46,10'd354};
ram[35838] = {-9'd43,10'd358};
ram[35839] = {-9'd40,10'd361};
ram[35840] = {-9'd40,10'd361};
ram[35841] = {-9'd37,10'd364};
ram[35842] = {-9'd33,10'd367};
ram[35843] = {-9'd30,10'd370};
ram[35844] = {-9'd27,10'd373};
ram[35845] = {-9'd24,10'd376};
ram[35846] = {-9'd21,10'd380};
ram[35847] = {-9'd18,10'd383};
ram[35848] = {-9'd15,10'd386};
ram[35849] = {-9'd11,10'd389};
ram[35850] = {-9'd8,10'd392};
ram[35851] = {-9'd5,10'd395};
ram[35852] = {-9'd2,10'd398};
ram[35853] = {9'd1,-10'd399};
ram[35854] = {9'd4,-10'd396};
ram[35855] = {9'd7,-10'd393};
ram[35856] = {9'd10,-10'd390};
ram[35857] = {9'd14,-10'd387};
ram[35858] = {9'd17,-10'd384};
ram[35859] = {9'd20,-10'd381};
ram[35860] = {9'd23,-10'd377};
ram[35861] = {9'd26,-10'd374};
ram[35862] = {9'd29,-10'd371};
ram[35863] = {9'd32,-10'd368};
ram[35864] = {9'd36,-10'd365};
ram[35865] = {9'd39,-10'd362};
ram[35866] = {9'd42,-10'd359};
ram[35867] = {9'd45,-10'd355};
ram[35868] = {9'd48,-10'd352};
ram[35869] = {9'd51,-10'd349};
ram[35870] = {9'd54,-10'd346};
ram[35871] = {9'd58,-10'd343};
ram[35872] = {9'd61,-10'd340};
ram[35873] = {9'd64,-10'd337};
ram[35874] = {9'd67,-10'd334};
ram[35875] = {9'd70,-10'd330};
ram[35876] = {9'd73,-10'd327};
ram[35877] = {9'd76,-10'd324};
ram[35878] = {9'd80,-10'd321};
ram[35879] = {9'd83,-10'd318};
ram[35880] = {9'd86,-10'd315};
ram[35881] = {9'd89,-10'd312};
ram[35882] = {9'd92,-10'd308};
ram[35883] = {9'd95,-10'd305};
ram[35884] = {9'd98,-10'd302};
ram[35885] = {-9'd99,-10'd299};
ram[35886] = {-9'd96,-10'd296};
ram[35887] = {-9'd92,-10'd293};
ram[35888] = {-9'd89,-10'd290};
ram[35889] = {-9'd86,-10'd286};
ram[35890] = {-9'd83,-10'd283};
ram[35891] = {-9'd80,-10'd280};
ram[35892] = {-9'd77,-10'd277};
ram[35893] = {-9'd74,-10'd274};
ram[35894] = {-9'd70,-10'd271};
ram[35895] = {-9'd67,-10'd268};
ram[35896] = {-9'd64,-10'd264};
ram[35897] = {-9'd61,-10'd261};
ram[35898] = {-9'd58,-10'd258};
ram[35899] = {-9'd55,-10'd255};
ram[35900] = {-9'd52,-10'd252};
ram[35901] = {-9'd48,-10'd249};
ram[35902] = {-9'd45,-10'd246};
ram[35903] = {-9'd42,-10'd242};
ram[35904] = {-9'd39,-10'd239};
ram[35905] = {-9'd36,-10'd236};
ram[35906] = {-9'd33,-10'd233};
ram[35907] = {-9'd30,-10'd230};
ram[35908] = {-9'd26,-10'd227};
ram[35909] = {-9'd23,-10'd224};
ram[35910] = {-9'd20,-10'd220};
ram[35911] = {-9'd17,-10'd217};
ram[35912] = {-9'd14,-10'd214};
ram[35913] = {-9'd11,-10'd211};
ram[35914] = {-9'd8,-10'd208};
ram[35915] = {-9'd4,-10'd205};
ram[35916] = {-9'd1,-10'd202};
ram[35917] = {9'd2,-10'd198};
ram[35918] = {9'd5,-10'd195};
ram[35919] = {9'd8,-10'd192};
ram[35920] = {9'd11,-10'd189};
ram[35921] = {9'd14,-10'd186};
ram[35922] = {9'd18,-10'd183};
ram[35923] = {9'd21,-10'd180};
ram[35924] = {9'd24,-10'd176};
ram[35925] = {9'd27,-10'd173};
ram[35926] = {9'd30,-10'd170};
ram[35927] = {9'd33,-10'd167};
ram[35928] = {9'd36,-10'd164};
ram[35929] = {9'd40,-10'd161};
ram[35930] = {9'd43,-10'd158};
ram[35931] = {9'd46,-10'd154};
ram[35932] = {9'd49,-10'd151};
ram[35933] = {9'd52,-10'd148};
ram[35934] = {9'd55,-10'd145};
ram[35935] = {9'd58,-10'd142};
ram[35936] = {9'd62,-10'd139};
ram[35937] = {9'd65,-10'd136};
ram[35938] = {9'd68,-10'd132};
ram[35939] = {9'd71,-10'd129};
ram[35940] = {9'd74,-10'd126};
ram[35941] = {9'd77,-10'd123};
ram[35942] = {9'd80,-10'd120};
ram[35943] = {9'd84,-10'd117};
ram[35944] = {9'd87,-10'd114};
ram[35945] = {9'd90,-10'd110};
ram[35946] = {9'd93,-10'd107};
ram[35947] = {9'd96,-10'd104};
ram[35948] = {9'd99,-10'd101};
ram[35949] = {-9'd98,-10'd98};
ram[35950] = {-9'd95,-10'd95};
ram[35951] = {-9'd92,-10'd92};
ram[35952] = {-9'd88,-10'd88};
ram[35953] = {-9'd85,-10'd85};
ram[35954] = {-9'd82,-10'd82};
ram[35955] = {-9'd79,-10'd79};
ram[35956] = {-9'd76,-10'd76};
ram[35957] = {-9'd73,-10'd73};
ram[35958] = {-9'd70,-10'd70};
ram[35959] = {-9'd66,-10'd66};
ram[35960] = {-9'd63,-10'd63};
ram[35961] = {-9'd60,-10'd60};
ram[35962] = {-9'd57,-10'd57};
ram[35963] = {-9'd54,-10'd54};
ram[35964] = {-9'd51,-10'd51};
ram[35965] = {-9'd48,-10'd48};
ram[35966] = {-9'd44,-10'd44};
ram[35967] = {-9'd41,-10'd41};
ram[35968] = {-9'd41,-10'd41};
ram[35969] = {-9'd38,-10'd38};
ram[35970] = {-9'd35,-10'd35};
ram[35971] = {-9'd32,-10'd32};
ram[35972] = {-9'd29,-10'd29};
ram[35973] = {-9'd26,-10'd26};
ram[35974] = {-9'd22,-10'd22};
ram[35975] = {-9'd19,-10'd19};
ram[35976] = {-9'd16,-10'd16};
ram[35977] = {-9'd13,-10'd13};
ram[35978] = {-9'd10,-10'd10};
ram[35979] = {-9'd7,-10'd7};
ram[35980] = {-9'd4,-10'd4};
ram[35981] = {9'd0,10'd0};
ram[35982] = {9'd3,10'd3};
ram[35983] = {9'd6,10'd6};
ram[35984] = {9'd9,10'd9};
ram[35985] = {9'd12,10'd12};
ram[35986] = {9'd15,10'd15};
ram[35987] = {9'd18,10'd18};
ram[35988] = {9'd21,10'd21};
ram[35989] = {9'd25,10'd25};
ram[35990] = {9'd28,10'd28};
ram[35991] = {9'd31,10'd31};
ram[35992] = {9'd34,10'd34};
ram[35993] = {9'd37,10'd37};
ram[35994] = {9'd40,10'd40};
ram[35995] = {9'd43,10'd43};
ram[35996] = {9'd47,10'd47};
ram[35997] = {9'd50,10'd50};
ram[35998] = {9'd53,10'd53};
ram[35999] = {9'd56,10'd56};
ram[36000] = {9'd59,10'd59};
ram[36001] = {9'd62,10'd62};
ram[36002] = {9'd65,10'd65};
ram[36003] = {9'd69,10'd69};
ram[36004] = {9'd72,10'd72};
ram[36005] = {9'd75,10'd75};
ram[36006] = {9'd78,10'd78};
ram[36007] = {9'd81,10'd81};
ram[36008] = {9'd84,10'd84};
ram[36009] = {9'd87,10'd87};
ram[36010] = {9'd91,10'd91};
ram[36011] = {9'd94,10'd94};
ram[36012] = {9'd97,10'd97};
ram[36013] = {-9'd100,10'd100};
ram[36014] = {-9'd97,10'd103};
ram[36015] = {-9'd94,10'd106};
ram[36016] = {-9'd91,10'd109};
ram[36017] = {-9'd88,10'd113};
ram[36018] = {-9'd85,10'd116};
ram[36019] = {-9'd81,10'd119};
ram[36020] = {-9'd78,10'd122};
ram[36021] = {-9'd75,10'd125};
ram[36022] = {-9'd72,10'd128};
ram[36023] = {-9'd69,10'd131};
ram[36024] = {-9'd66,10'd135};
ram[36025] = {-9'd63,10'd138};
ram[36026] = {-9'd59,10'd141};
ram[36027] = {-9'd56,10'd144};
ram[36028] = {-9'd53,10'd147};
ram[36029] = {-9'd50,10'd150};
ram[36030] = {-9'd47,10'd153};
ram[36031] = {-9'd44,10'd157};
ram[36032] = {-9'd41,10'd160};
ram[36033] = {-9'd37,10'd163};
ram[36034] = {-9'd34,10'd166};
ram[36035] = {-9'd31,10'd169};
ram[36036] = {-9'd28,10'd172};
ram[36037] = {-9'd25,10'd175};
ram[36038] = {-9'd22,10'd179};
ram[36039] = {-9'd19,10'd182};
ram[36040] = {-9'd15,10'd185};
ram[36041] = {-9'd12,10'd188};
ram[36042] = {-9'd9,10'd191};
ram[36043] = {-9'd6,10'd194};
ram[36044] = {-9'd3,10'd197};
ram[36045] = {9'd0,10'd201};
ram[36046] = {9'd3,10'd204};
ram[36047] = {9'd7,10'd207};
ram[36048] = {9'd10,10'd210};
ram[36049] = {9'd13,10'd213};
ram[36050] = {9'd16,10'd216};
ram[36051] = {9'd19,10'd219};
ram[36052] = {9'd22,10'd223};
ram[36053] = {9'd25,10'd226};
ram[36054] = {9'd29,10'd229};
ram[36055] = {9'd32,10'd232};
ram[36056] = {9'd35,10'd235};
ram[36057] = {9'd38,10'd238};
ram[36058] = {9'd41,10'd241};
ram[36059] = {9'd44,10'd245};
ram[36060] = {9'd47,10'd248};
ram[36061] = {9'd51,10'd251};
ram[36062] = {9'd54,10'd254};
ram[36063] = {9'd57,10'd257};
ram[36064] = {9'd60,10'd260};
ram[36065] = {9'd63,10'd263};
ram[36066] = {9'd66,10'd267};
ram[36067] = {9'd69,10'd270};
ram[36068] = {9'd73,10'd273};
ram[36069] = {9'd76,10'd276};
ram[36070] = {9'd79,10'd279};
ram[36071] = {9'd82,10'd282};
ram[36072] = {9'd85,10'd285};
ram[36073] = {9'd88,10'd289};
ram[36074] = {9'd91,10'd292};
ram[36075] = {9'd95,10'd295};
ram[36076] = {9'd98,10'd298};
ram[36077] = {-9'd99,10'd301};
ram[36078] = {-9'd96,10'd304};
ram[36079] = {-9'd93,10'd307};
ram[36080] = {-9'd90,10'd311};
ram[36081] = {-9'd87,10'd314};
ram[36082] = {-9'd84,10'd317};
ram[36083] = {-9'd81,10'd320};
ram[36084] = {-9'd77,10'd323};
ram[36085] = {-9'd74,10'd326};
ram[36086] = {-9'd71,10'd329};
ram[36087] = {-9'd68,10'd333};
ram[36088] = {-9'd65,10'd336};
ram[36089] = {-9'd62,10'd339};
ram[36090] = {-9'd59,10'd342};
ram[36091] = {-9'd55,10'd345};
ram[36092] = {-9'd52,10'd348};
ram[36093] = {-9'd49,10'd351};
ram[36094] = {-9'd46,10'd354};
ram[36095] = {-9'd43,10'd358};
ram[36096] = {-9'd43,10'd358};
ram[36097] = {-9'd40,10'd361};
ram[36098] = {-9'd37,10'd364};
ram[36099] = {-9'd33,10'd367};
ram[36100] = {-9'd30,10'd370};
ram[36101] = {-9'd27,10'd373};
ram[36102] = {-9'd24,10'd376};
ram[36103] = {-9'd21,10'd380};
ram[36104] = {-9'd18,10'd383};
ram[36105] = {-9'd15,10'd386};
ram[36106] = {-9'd11,10'd389};
ram[36107] = {-9'd8,10'd392};
ram[36108] = {-9'd5,10'd395};
ram[36109] = {-9'd2,10'd398};
ram[36110] = {9'd1,-10'd399};
ram[36111] = {9'd4,-10'd396};
ram[36112] = {9'd7,-10'd393};
ram[36113] = {9'd10,-10'd390};
ram[36114] = {9'd14,-10'd387};
ram[36115] = {9'd17,-10'd384};
ram[36116] = {9'd20,-10'd381};
ram[36117] = {9'd23,-10'd377};
ram[36118] = {9'd26,-10'd374};
ram[36119] = {9'd29,-10'd371};
ram[36120] = {9'd32,-10'd368};
ram[36121] = {9'd36,-10'd365};
ram[36122] = {9'd39,-10'd362};
ram[36123] = {9'd42,-10'd359};
ram[36124] = {9'd45,-10'd355};
ram[36125] = {9'd48,-10'd352};
ram[36126] = {9'd51,-10'd349};
ram[36127] = {9'd54,-10'd346};
ram[36128] = {9'd58,-10'd343};
ram[36129] = {9'd61,-10'd340};
ram[36130] = {9'd64,-10'd337};
ram[36131] = {9'd67,-10'd334};
ram[36132] = {9'd70,-10'd330};
ram[36133] = {9'd73,-10'd327};
ram[36134] = {9'd76,-10'd324};
ram[36135] = {9'd80,-10'd321};
ram[36136] = {9'd83,-10'd318};
ram[36137] = {9'd86,-10'd315};
ram[36138] = {9'd89,-10'd312};
ram[36139] = {9'd92,-10'd308};
ram[36140] = {9'd95,-10'd305};
ram[36141] = {9'd98,-10'd302};
ram[36142] = {-9'd99,-10'd299};
ram[36143] = {-9'd96,-10'd296};
ram[36144] = {-9'd92,-10'd293};
ram[36145] = {-9'd89,-10'd290};
ram[36146] = {-9'd86,-10'd286};
ram[36147] = {-9'd83,-10'd283};
ram[36148] = {-9'd80,-10'd280};
ram[36149] = {-9'd77,-10'd277};
ram[36150] = {-9'd74,-10'd274};
ram[36151] = {-9'd70,-10'd271};
ram[36152] = {-9'd67,-10'd268};
ram[36153] = {-9'd64,-10'd264};
ram[36154] = {-9'd61,-10'd261};
ram[36155] = {-9'd58,-10'd258};
ram[36156] = {-9'd55,-10'd255};
ram[36157] = {-9'd52,-10'd252};
ram[36158] = {-9'd48,-10'd249};
ram[36159] = {-9'd45,-10'd246};
ram[36160] = {-9'd42,-10'd242};
ram[36161] = {-9'd39,-10'd239};
ram[36162] = {-9'd36,-10'd236};
ram[36163] = {-9'd33,-10'd233};
ram[36164] = {-9'd30,-10'd230};
ram[36165] = {-9'd26,-10'd227};
ram[36166] = {-9'd23,-10'd224};
ram[36167] = {-9'd20,-10'd220};
ram[36168] = {-9'd17,-10'd217};
ram[36169] = {-9'd14,-10'd214};
ram[36170] = {-9'd11,-10'd211};
ram[36171] = {-9'd8,-10'd208};
ram[36172] = {-9'd4,-10'd205};
ram[36173] = {-9'd1,-10'd202};
ram[36174] = {9'd2,-10'd198};
ram[36175] = {9'd5,-10'd195};
ram[36176] = {9'd8,-10'd192};
ram[36177] = {9'd11,-10'd189};
ram[36178] = {9'd14,-10'd186};
ram[36179] = {9'd18,-10'd183};
ram[36180] = {9'd21,-10'd180};
ram[36181] = {9'd24,-10'd176};
ram[36182] = {9'd27,-10'd173};
ram[36183] = {9'd30,-10'd170};
ram[36184] = {9'd33,-10'd167};
ram[36185] = {9'd36,-10'd164};
ram[36186] = {9'd40,-10'd161};
ram[36187] = {9'd43,-10'd158};
ram[36188] = {9'd46,-10'd154};
ram[36189] = {9'd49,-10'd151};
ram[36190] = {9'd52,-10'd148};
ram[36191] = {9'd55,-10'd145};
ram[36192] = {9'd58,-10'd142};
ram[36193] = {9'd62,-10'd139};
ram[36194] = {9'd65,-10'd136};
ram[36195] = {9'd68,-10'd132};
ram[36196] = {9'd71,-10'd129};
ram[36197] = {9'd74,-10'd126};
ram[36198] = {9'd77,-10'd123};
ram[36199] = {9'd80,-10'd120};
ram[36200] = {9'd84,-10'd117};
ram[36201] = {9'd87,-10'd114};
ram[36202] = {9'd90,-10'd110};
ram[36203] = {9'd93,-10'd107};
ram[36204] = {9'd96,-10'd104};
ram[36205] = {9'd99,-10'd101};
ram[36206] = {-9'd98,-10'd98};
ram[36207] = {-9'd95,-10'd95};
ram[36208] = {-9'd92,-10'd92};
ram[36209] = {-9'd88,-10'd88};
ram[36210] = {-9'd85,-10'd85};
ram[36211] = {-9'd82,-10'd82};
ram[36212] = {-9'd79,-10'd79};
ram[36213] = {-9'd76,-10'd76};
ram[36214] = {-9'd73,-10'd73};
ram[36215] = {-9'd70,-10'd70};
ram[36216] = {-9'd66,-10'd66};
ram[36217] = {-9'd63,-10'd63};
ram[36218] = {-9'd60,-10'd60};
ram[36219] = {-9'd57,-10'd57};
ram[36220] = {-9'd54,-10'd54};
ram[36221] = {-9'd51,-10'd51};
ram[36222] = {-9'd48,-10'd48};
ram[36223] = {-9'd44,-10'd44};
ram[36224] = {-9'd44,-10'd44};
ram[36225] = {-9'd41,-10'd41};
ram[36226] = {-9'd38,-10'd38};
ram[36227] = {-9'd35,-10'd35};
ram[36228] = {-9'd32,-10'd32};
ram[36229] = {-9'd29,-10'd29};
ram[36230] = {-9'd26,-10'd26};
ram[36231] = {-9'd22,-10'd22};
ram[36232] = {-9'd19,-10'd19};
ram[36233] = {-9'd16,-10'd16};
ram[36234] = {-9'd13,-10'd13};
ram[36235] = {-9'd10,-10'd10};
ram[36236] = {-9'd7,-10'd7};
ram[36237] = {-9'd4,-10'd4};
ram[36238] = {9'd0,10'd0};
ram[36239] = {9'd3,10'd3};
ram[36240] = {9'd6,10'd6};
ram[36241] = {9'd9,10'd9};
ram[36242] = {9'd12,10'd12};
ram[36243] = {9'd15,10'd15};
ram[36244] = {9'd18,10'd18};
ram[36245] = {9'd21,10'd21};
ram[36246] = {9'd25,10'd25};
ram[36247] = {9'd28,10'd28};
ram[36248] = {9'd31,10'd31};
ram[36249] = {9'd34,10'd34};
ram[36250] = {9'd37,10'd37};
ram[36251] = {9'd40,10'd40};
ram[36252] = {9'd43,10'd43};
ram[36253] = {9'd47,10'd47};
ram[36254] = {9'd50,10'd50};
ram[36255] = {9'd53,10'd53};
ram[36256] = {9'd56,10'd56};
ram[36257] = {9'd59,10'd59};
ram[36258] = {9'd62,10'd62};
ram[36259] = {9'd65,10'd65};
ram[36260] = {9'd69,10'd69};
ram[36261] = {9'd72,10'd72};
ram[36262] = {9'd75,10'd75};
ram[36263] = {9'd78,10'd78};
ram[36264] = {9'd81,10'd81};
ram[36265] = {9'd84,10'd84};
ram[36266] = {9'd87,10'd87};
ram[36267] = {9'd91,10'd91};
ram[36268] = {9'd94,10'd94};
ram[36269] = {9'd97,10'd97};
ram[36270] = {-9'd100,10'd100};
ram[36271] = {-9'd97,10'd103};
ram[36272] = {-9'd94,10'd106};
ram[36273] = {-9'd91,10'd109};
ram[36274] = {-9'd88,10'd113};
ram[36275] = {-9'd85,10'd116};
ram[36276] = {-9'd81,10'd119};
ram[36277] = {-9'd78,10'd122};
ram[36278] = {-9'd75,10'd125};
ram[36279] = {-9'd72,10'd128};
ram[36280] = {-9'd69,10'd131};
ram[36281] = {-9'd66,10'd135};
ram[36282] = {-9'd63,10'd138};
ram[36283] = {-9'd59,10'd141};
ram[36284] = {-9'd56,10'd144};
ram[36285] = {-9'd53,10'd147};
ram[36286] = {-9'd50,10'd150};
ram[36287] = {-9'd47,10'd153};
ram[36288] = {-9'd44,10'd157};
ram[36289] = {-9'd41,10'd160};
ram[36290] = {-9'd37,10'd163};
ram[36291] = {-9'd34,10'd166};
ram[36292] = {-9'd31,10'd169};
ram[36293] = {-9'd28,10'd172};
ram[36294] = {-9'd25,10'd175};
ram[36295] = {-9'd22,10'd179};
ram[36296] = {-9'd19,10'd182};
ram[36297] = {-9'd15,10'd185};
ram[36298] = {-9'd12,10'd188};
ram[36299] = {-9'd9,10'd191};
ram[36300] = {-9'd6,10'd194};
ram[36301] = {-9'd3,10'd197};
ram[36302] = {9'd0,10'd201};
ram[36303] = {9'd3,10'd204};
ram[36304] = {9'd7,10'd207};
ram[36305] = {9'd10,10'd210};
ram[36306] = {9'd13,10'd213};
ram[36307] = {9'd16,10'd216};
ram[36308] = {9'd19,10'd219};
ram[36309] = {9'd22,10'd223};
ram[36310] = {9'd25,10'd226};
ram[36311] = {9'd29,10'd229};
ram[36312] = {9'd32,10'd232};
ram[36313] = {9'd35,10'd235};
ram[36314] = {9'd38,10'd238};
ram[36315] = {9'd41,10'd241};
ram[36316] = {9'd44,10'd245};
ram[36317] = {9'd47,10'd248};
ram[36318] = {9'd51,10'd251};
ram[36319] = {9'd54,10'd254};
ram[36320] = {9'd57,10'd257};
ram[36321] = {9'd60,10'd260};
ram[36322] = {9'd63,10'd263};
ram[36323] = {9'd66,10'd267};
ram[36324] = {9'd69,10'd270};
ram[36325] = {9'd73,10'd273};
ram[36326] = {9'd76,10'd276};
ram[36327] = {9'd79,10'd279};
ram[36328] = {9'd82,10'd282};
ram[36329] = {9'd85,10'd285};
ram[36330] = {9'd88,10'd289};
ram[36331] = {9'd91,10'd292};
ram[36332] = {9'd95,10'd295};
ram[36333] = {9'd98,10'd298};
ram[36334] = {-9'd99,10'd301};
ram[36335] = {-9'd96,10'd304};
ram[36336] = {-9'd93,10'd307};
ram[36337] = {-9'd90,10'd311};
ram[36338] = {-9'd87,10'd314};
ram[36339] = {-9'd84,10'd317};
ram[36340] = {-9'd81,10'd320};
ram[36341] = {-9'd77,10'd323};
ram[36342] = {-9'd74,10'd326};
ram[36343] = {-9'd71,10'd329};
ram[36344] = {-9'd68,10'd333};
ram[36345] = {-9'd65,10'd336};
ram[36346] = {-9'd62,10'd339};
ram[36347] = {-9'd59,10'd342};
ram[36348] = {-9'd55,10'd345};
ram[36349] = {-9'd52,10'd348};
ram[36350] = {-9'd49,10'd351};
ram[36351] = {-9'd46,10'd354};
ram[36352] = {-9'd46,10'd354};
ram[36353] = {-9'd43,10'd358};
ram[36354] = {-9'd40,10'd361};
ram[36355] = {-9'd37,10'd364};
ram[36356] = {-9'd33,10'd367};
ram[36357] = {-9'd30,10'd370};
ram[36358] = {-9'd27,10'd373};
ram[36359] = {-9'd24,10'd376};
ram[36360] = {-9'd21,10'd380};
ram[36361] = {-9'd18,10'd383};
ram[36362] = {-9'd15,10'd386};
ram[36363] = {-9'd11,10'd389};
ram[36364] = {-9'd8,10'd392};
ram[36365] = {-9'd5,10'd395};
ram[36366] = {-9'd2,10'd398};
ram[36367] = {9'd1,-10'd399};
ram[36368] = {9'd4,-10'd396};
ram[36369] = {9'd7,-10'd393};
ram[36370] = {9'd10,-10'd390};
ram[36371] = {9'd14,-10'd387};
ram[36372] = {9'd17,-10'd384};
ram[36373] = {9'd20,-10'd381};
ram[36374] = {9'd23,-10'd377};
ram[36375] = {9'd26,-10'd374};
ram[36376] = {9'd29,-10'd371};
ram[36377] = {9'd32,-10'd368};
ram[36378] = {9'd36,-10'd365};
ram[36379] = {9'd39,-10'd362};
ram[36380] = {9'd42,-10'd359};
ram[36381] = {9'd45,-10'd355};
ram[36382] = {9'd48,-10'd352};
ram[36383] = {9'd51,-10'd349};
ram[36384] = {9'd54,-10'd346};
ram[36385] = {9'd58,-10'd343};
ram[36386] = {9'd61,-10'd340};
ram[36387] = {9'd64,-10'd337};
ram[36388] = {9'd67,-10'd334};
ram[36389] = {9'd70,-10'd330};
ram[36390] = {9'd73,-10'd327};
ram[36391] = {9'd76,-10'd324};
ram[36392] = {9'd80,-10'd321};
ram[36393] = {9'd83,-10'd318};
ram[36394] = {9'd86,-10'd315};
ram[36395] = {9'd89,-10'd312};
ram[36396] = {9'd92,-10'd308};
ram[36397] = {9'd95,-10'd305};
ram[36398] = {9'd98,-10'd302};
ram[36399] = {-9'd99,-10'd299};
ram[36400] = {-9'd96,-10'd296};
ram[36401] = {-9'd92,-10'd293};
ram[36402] = {-9'd89,-10'd290};
ram[36403] = {-9'd86,-10'd286};
ram[36404] = {-9'd83,-10'd283};
ram[36405] = {-9'd80,-10'd280};
ram[36406] = {-9'd77,-10'd277};
ram[36407] = {-9'd74,-10'd274};
ram[36408] = {-9'd70,-10'd271};
ram[36409] = {-9'd67,-10'd268};
ram[36410] = {-9'd64,-10'd264};
ram[36411] = {-9'd61,-10'd261};
ram[36412] = {-9'd58,-10'd258};
ram[36413] = {-9'd55,-10'd255};
ram[36414] = {-9'd52,-10'd252};
ram[36415] = {-9'd48,-10'd249};
ram[36416] = {-9'd45,-10'd246};
ram[36417] = {-9'd42,-10'd242};
ram[36418] = {-9'd39,-10'd239};
ram[36419] = {-9'd36,-10'd236};
ram[36420] = {-9'd33,-10'd233};
ram[36421] = {-9'd30,-10'd230};
ram[36422] = {-9'd26,-10'd227};
ram[36423] = {-9'd23,-10'd224};
ram[36424] = {-9'd20,-10'd220};
ram[36425] = {-9'd17,-10'd217};
ram[36426] = {-9'd14,-10'd214};
ram[36427] = {-9'd11,-10'd211};
ram[36428] = {-9'd8,-10'd208};
ram[36429] = {-9'd4,-10'd205};
ram[36430] = {-9'd1,-10'd202};
ram[36431] = {9'd2,-10'd198};
ram[36432] = {9'd5,-10'd195};
ram[36433] = {9'd8,-10'd192};
ram[36434] = {9'd11,-10'd189};
ram[36435] = {9'd14,-10'd186};
ram[36436] = {9'd18,-10'd183};
ram[36437] = {9'd21,-10'd180};
ram[36438] = {9'd24,-10'd176};
ram[36439] = {9'd27,-10'd173};
ram[36440] = {9'd30,-10'd170};
ram[36441] = {9'd33,-10'd167};
ram[36442] = {9'd36,-10'd164};
ram[36443] = {9'd40,-10'd161};
ram[36444] = {9'd43,-10'd158};
ram[36445] = {9'd46,-10'd154};
ram[36446] = {9'd49,-10'd151};
ram[36447] = {9'd52,-10'd148};
ram[36448] = {9'd55,-10'd145};
ram[36449] = {9'd58,-10'd142};
ram[36450] = {9'd62,-10'd139};
ram[36451] = {9'd65,-10'd136};
ram[36452] = {9'd68,-10'd132};
ram[36453] = {9'd71,-10'd129};
ram[36454] = {9'd74,-10'd126};
ram[36455] = {9'd77,-10'd123};
ram[36456] = {9'd80,-10'd120};
ram[36457] = {9'd84,-10'd117};
ram[36458] = {9'd87,-10'd114};
ram[36459] = {9'd90,-10'd110};
ram[36460] = {9'd93,-10'd107};
ram[36461] = {9'd96,-10'd104};
ram[36462] = {9'd99,-10'd101};
ram[36463] = {-9'd98,-10'd98};
ram[36464] = {-9'd95,-10'd95};
ram[36465] = {-9'd92,-10'd92};
ram[36466] = {-9'd88,-10'd88};
ram[36467] = {-9'd85,-10'd85};
ram[36468] = {-9'd82,-10'd82};
ram[36469] = {-9'd79,-10'd79};
ram[36470] = {-9'd76,-10'd76};
ram[36471] = {-9'd73,-10'd73};
ram[36472] = {-9'd70,-10'd70};
ram[36473] = {-9'd66,-10'd66};
ram[36474] = {-9'd63,-10'd63};
ram[36475] = {-9'd60,-10'd60};
ram[36476] = {-9'd57,-10'd57};
ram[36477] = {-9'd54,-10'd54};
ram[36478] = {-9'd51,-10'd51};
ram[36479] = {-9'd48,-10'd48};
ram[36480] = {-9'd48,-10'd48};
ram[36481] = {-9'd44,-10'd44};
ram[36482] = {-9'd41,-10'd41};
ram[36483] = {-9'd38,-10'd38};
ram[36484] = {-9'd35,-10'd35};
ram[36485] = {-9'd32,-10'd32};
ram[36486] = {-9'd29,-10'd29};
ram[36487] = {-9'd26,-10'd26};
ram[36488] = {-9'd22,-10'd22};
ram[36489] = {-9'd19,-10'd19};
ram[36490] = {-9'd16,-10'd16};
ram[36491] = {-9'd13,-10'd13};
ram[36492] = {-9'd10,-10'd10};
ram[36493] = {-9'd7,-10'd7};
ram[36494] = {-9'd4,-10'd4};
ram[36495] = {9'd0,10'd0};
ram[36496] = {9'd3,10'd3};
ram[36497] = {9'd6,10'd6};
ram[36498] = {9'd9,10'd9};
ram[36499] = {9'd12,10'd12};
ram[36500] = {9'd15,10'd15};
ram[36501] = {9'd18,10'd18};
ram[36502] = {9'd21,10'd21};
ram[36503] = {9'd25,10'd25};
ram[36504] = {9'd28,10'd28};
ram[36505] = {9'd31,10'd31};
ram[36506] = {9'd34,10'd34};
ram[36507] = {9'd37,10'd37};
ram[36508] = {9'd40,10'd40};
ram[36509] = {9'd43,10'd43};
ram[36510] = {9'd47,10'd47};
ram[36511] = {9'd50,10'd50};
ram[36512] = {9'd53,10'd53};
ram[36513] = {9'd56,10'd56};
ram[36514] = {9'd59,10'd59};
ram[36515] = {9'd62,10'd62};
ram[36516] = {9'd65,10'd65};
ram[36517] = {9'd69,10'd69};
ram[36518] = {9'd72,10'd72};
ram[36519] = {9'd75,10'd75};
ram[36520] = {9'd78,10'd78};
ram[36521] = {9'd81,10'd81};
ram[36522] = {9'd84,10'd84};
ram[36523] = {9'd87,10'd87};
ram[36524] = {9'd91,10'd91};
ram[36525] = {9'd94,10'd94};
ram[36526] = {9'd97,10'd97};
ram[36527] = {-9'd100,10'd100};
ram[36528] = {-9'd97,10'd103};
ram[36529] = {-9'd94,10'd106};
ram[36530] = {-9'd91,10'd109};
ram[36531] = {-9'd88,10'd113};
ram[36532] = {-9'd85,10'd116};
ram[36533] = {-9'd81,10'd119};
ram[36534] = {-9'd78,10'd122};
ram[36535] = {-9'd75,10'd125};
ram[36536] = {-9'd72,10'd128};
ram[36537] = {-9'd69,10'd131};
ram[36538] = {-9'd66,10'd135};
ram[36539] = {-9'd63,10'd138};
ram[36540] = {-9'd59,10'd141};
ram[36541] = {-9'd56,10'd144};
ram[36542] = {-9'd53,10'd147};
ram[36543] = {-9'd50,10'd150};
ram[36544] = {-9'd47,10'd153};
ram[36545] = {-9'd44,10'd157};
ram[36546] = {-9'd41,10'd160};
ram[36547] = {-9'd37,10'd163};
ram[36548] = {-9'd34,10'd166};
ram[36549] = {-9'd31,10'd169};
ram[36550] = {-9'd28,10'd172};
ram[36551] = {-9'd25,10'd175};
ram[36552] = {-9'd22,10'd179};
ram[36553] = {-9'd19,10'd182};
ram[36554] = {-9'd15,10'd185};
ram[36555] = {-9'd12,10'd188};
ram[36556] = {-9'd9,10'd191};
ram[36557] = {-9'd6,10'd194};
ram[36558] = {-9'd3,10'd197};
ram[36559] = {9'd0,10'd201};
ram[36560] = {9'd3,10'd204};
ram[36561] = {9'd7,10'd207};
ram[36562] = {9'd10,10'd210};
ram[36563] = {9'd13,10'd213};
ram[36564] = {9'd16,10'd216};
ram[36565] = {9'd19,10'd219};
ram[36566] = {9'd22,10'd223};
ram[36567] = {9'd25,10'd226};
ram[36568] = {9'd29,10'd229};
ram[36569] = {9'd32,10'd232};
ram[36570] = {9'd35,10'd235};
ram[36571] = {9'd38,10'd238};
ram[36572] = {9'd41,10'd241};
ram[36573] = {9'd44,10'd245};
ram[36574] = {9'd47,10'd248};
ram[36575] = {9'd51,10'd251};
ram[36576] = {9'd54,10'd254};
ram[36577] = {9'd57,10'd257};
ram[36578] = {9'd60,10'd260};
ram[36579] = {9'd63,10'd263};
ram[36580] = {9'd66,10'd267};
ram[36581] = {9'd69,10'd270};
ram[36582] = {9'd73,10'd273};
ram[36583] = {9'd76,10'd276};
ram[36584] = {9'd79,10'd279};
ram[36585] = {9'd82,10'd282};
ram[36586] = {9'd85,10'd285};
ram[36587] = {9'd88,10'd289};
ram[36588] = {9'd91,10'd292};
ram[36589] = {9'd95,10'd295};
ram[36590] = {9'd98,10'd298};
ram[36591] = {-9'd99,10'd301};
ram[36592] = {-9'd96,10'd304};
ram[36593] = {-9'd93,10'd307};
ram[36594] = {-9'd90,10'd311};
ram[36595] = {-9'd87,10'd314};
ram[36596] = {-9'd84,10'd317};
ram[36597] = {-9'd81,10'd320};
ram[36598] = {-9'd77,10'd323};
ram[36599] = {-9'd74,10'd326};
ram[36600] = {-9'd71,10'd329};
ram[36601] = {-9'd68,10'd333};
ram[36602] = {-9'd65,10'd336};
ram[36603] = {-9'd62,10'd339};
ram[36604] = {-9'd59,10'd342};
ram[36605] = {-9'd55,10'd345};
ram[36606] = {-9'd52,10'd348};
ram[36607] = {-9'd49,10'd351};
ram[36608] = {-9'd49,10'd351};
ram[36609] = {-9'd46,10'd354};
ram[36610] = {-9'd43,10'd358};
ram[36611] = {-9'd40,10'd361};
ram[36612] = {-9'd37,10'd364};
ram[36613] = {-9'd33,10'd367};
ram[36614] = {-9'd30,10'd370};
ram[36615] = {-9'd27,10'd373};
ram[36616] = {-9'd24,10'd376};
ram[36617] = {-9'd21,10'd380};
ram[36618] = {-9'd18,10'd383};
ram[36619] = {-9'd15,10'd386};
ram[36620] = {-9'd11,10'd389};
ram[36621] = {-9'd8,10'd392};
ram[36622] = {-9'd5,10'd395};
ram[36623] = {-9'd2,10'd398};
ram[36624] = {9'd1,-10'd399};
ram[36625] = {9'd4,-10'd396};
ram[36626] = {9'd7,-10'd393};
ram[36627] = {9'd10,-10'd390};
ram[36628] = {9'd14,-10'd387};
ram[36629] = {9'd17,-10'd384};
ram[36630] = {9'd20,-10'd381};
ram[36631] = {9'd23,-10'd377};
ram[36632] = {9'd26,-10'd374};
ram[36633] = {9'd29,-10'd371};
ram[36634] = {9'd32,-10'd368};
ram[36635] = {9'd36,-10'd365};
ram[36636] = {9'd39,-10'd362};
ram[36637] = {9'd42,-10'd359};
ram[36638] = {9'd45,-10'd355};
ram[36639] = {9'd48,-10'd352};
ram[36640] = {9'd51,-10'd349};
ram[36641] = {9'd54,-10'd346};
ram[36642] = {9'd58,-10'd343};
ram[36643] = {9'd61,-10'd340};
ram[36644] = {9'd64,-10'd337};
ram[36645] = {9'd67,-10'd334};
ram[36646] = {9'd70,-10'd330};
ram[36647] = {9'd73,-10'd327};
ram[36648] = {9'd76,-10'd324};
ram[36649] = {9'd80,-10'd321};
ram[36650] = {9'd83,-10'd318};
ram[36651] = {9'd86,-10'd315};
ram[36652] = {9'd89,-10'd312};
ram[36653] = {9'd92,-10'd308};
ram[36654] = {9'd95,-10'd305};
ram[36655] = {9'd98,-10'd302};
ram[36656] = {-9'd99,-10'd299};
ram[36657] = {-9'd96,-10'd296};
ram[36658] = {-9'd92,-10'd293};
ram[36659] = {-9'd89,-10'd290};
ram[36660] = {-9'd86,-10'd286};
ram[36661] = {-9'd83,-10'd283};
ram[36662] = {-9'd80,-10'd280};
ram[36663] = {-9'd77,-10'd277};
ram[36664] = {-9'd74,-10'd274};
ram[36665] = {-9'd70,-10'd271};
ram[36666] = {-9'd67,-10'd268};
ram[36667] = {-9'd64,-10'd264};
ram[36668] = {-9'd61,-10'd261};
ram[36669] = {-9'd58,-10'd258};
ram[36670] = {-9'd55,-10'd255};
ram[36671] = {-9'd52,-10'd252};
ram[36672] = {-9'd48,-10'd249};
ram[36673] = {-9'd45,-10'd246};
ram[36674] = {-9'd42,-10'd242};
ram[36675] = {-9'd39,-10'd239};
ram[36676] = {-9'd36,-10'd236};
ram[36677] = {-9'd33,-10'd233};
ram[36678] = {-9'd30,-10'd230};
ram[36679] = {-9'd26,-10'd227};
ram[36680] = {-9'd23,-10'd224};
ram[36681] = {-9'd20,-10'd220};
ram[36682] = {-9'd17,-10'd217};
ram[36683] = {-9'd14,-10'd214};
ram[36684] = {-9'd11,-10'd211};
ram[36685] = {-9'd8,-10'd208};
ram[36686] = {-9'd4,-10'd205};
ram[36687] = {-9'd1,-10'd202};
ram[36688] = {9'd2,-10'd198};
ram[36689] = {9'd5,-10'd195};
ram[36690] = {9'd8,-10'd192};
ram[36691] = {9'd11,-10'd189};
ram[36692] = {9'd14,-10'd186};
ram[36693] = {9'd18,-10'd183};
ram[36694] = {9'd21,-10'd180};
ram[36695] = {9'd24,-10'd176};
ram[36696] = {9'd27,-10'd173};
ram[36697] = {9'd30,-10'd170};
ram[36698] = {9'd33,-10'd167};
ram[36699] = {9'd36,-10'd164};
ram[36700] = {9'd40,-10'd161};
ram[36701] = {9'd43,-10'd158};
ram[36702] = {9'd46,-10'd154};
ram[36703] = {9'd49,-10'd151};
ram[36704] = {9'd52,-10'd148};
ram[36705] = {9'd55,-10'd145};
ram[36706] = {9'd58,-10'd142};
ram[36707] = {9'd62,-10'd139};
ram[36708] = {9'd65,-10'd136};
ram[36709] = {9'd68,-10'd132};
ram[36710] = {9'd71,-10'd129};
ram[36711] = {9'd74,-10'd126};
ram[36712] = {9'd77,-10'd123};
ram[36713] = {9'd80,-10'd120};
ram[36714] = {9'd84,-10'd117};
ram[36715] = {9'd87,-10'd114};
ram[36716] = {9'd90,-10'd110};
ram[36717] = {9'd93,-10'd107};
ram[36718] = {9'd96,-10'd104};
ram[36719] = {9'd99,-10'd101};
ram[36720] = {-9'd98,-10'd98};
ram[36721] = {-9'd95,-10'd95};
ram[36722] = {-9'd92,-10'd92};
ram[36723] = {-9'd88,-10'd88};
ram[36724] = {-9'd85,-10'd85};
ram[36725] = {-9'd82,-10'd82};
ram[36726] = {-9'd79,-10'd79};
ram[36727] = {-9'd76,-10'd76};
ram[36728] = {-9'd73,-10'd73};
ram[36729] = {-9'd70,-10'd70};
ram[36730] = {-9'd66,-10'd66};
ram[36731] = {-9'd63,-10'd63};
ram[36732] = {-9'd60,-10'd60};
ram[36733] = {-9'd57,-10'd57};
ram[36734] = {-9'd54,-10'd54};
ram[36735] = {-9'd51,-10'd51};
ram[36736] = {-9'd51,-10'd51};
ram[36737] = {-9'd48,-10'd48};
ram[36738] = {-9'd44,-10'd44};
ram[36739] = {-9'd41,-10'd41};
ram[36740] = {-9'd38,-10'd38};
ram[36741] = {-9'd35,-10'd35};
ram[36742] = {-9'd32,-10'd32};
ram[36743] = {-9'd29,-10'd29};
ram[36744] = {-9'd26,-10'd26};
ram[36745] = {-9'd22,-10'd22};
ram[36746] = {-9'd19,-10'd19};
ram[36747] = {-9'd16,-10'd16};
ram[36748] = {-9'd13,-10'd13};
ram[36749] = {-9'd10,-10'd10};
ram[36750] = {-9'd7,-10'd7};
ram[36751] = {-9'd4,-10'd4};
ram[36752] = {9'd0,10'd0};
ram[36753] = {9'd3,10'd3};
ram[36754] = {9'd6,10'd6};
ram[36755] = {9'd9,10'd9};
ram[36756] = {9'd12,10'd12};
ram[36757] = {9'd15,10'd15};
ram[36758] = {9'd18,10'd18};
ram[36759] = {9'd21,10'd21};
ram[36760] = {9'd25,10'd25};
ram[36761] = {9'd28,10'd28};
ram[36762] = {9'd31,10'd31};
ram[36763] = {9'd34,10'd34};
ram[36764] = {9'd37,10'd37};
ram[36765] = {9'd40,10'd40};
ram[36766] = {9'd43,10'd43};
ram[36767] = {9'd47,10'd47};
ram[36768] = {9'd50,10'd50};
ram[36769] = {9'd53,10'd53};
ram[36770] = {9'd56,10'd56};
ram[36771] = {9'd59,10'd59};
ram[36772] = {9'd62,10'd62};
ram[36773] = {9'd65,10'd65};
ram[36774] = {9'd69,10'd69};
ram[36775] = {9'd72,10'd72};
ram[36776] = {9'd75,10'd75};
ram[36777] = {9'd78,10'd78};
ram[36778] = {9'd81,10'd81};
ram[36779] = {9'd84,10'd84};
ram[36780] = {9'd87,10'd87};
ram[36781] = {9'd91,10'd91};
ram[36782] = {9'd94,10'd94};
ram[36783] = {9'd97,10'd97};
ram[36784] = {-9'd100,10'd100};
ram[36785] = {-9'd97,10'd103};
ram[36786] = {-9'd94,10'd106};
ram[36787] = {-9'd91,10'd109};
ram[36788] = {-9'd88,10'd113};
ram[36789] = {-9'd85,10'd116};
ram[36790] = {-9'd81,10'd119};
ram[36791] = {-9'd78,10'd122};
ram[36792] = {-9'd75,10'd125};
ram[36793] = {-9'd72,10'd128};
ram[36794] = {-9'd69,10'd131};
ram[36795] = {-9'd66,10'd135};
ram[36796] = {-9'd63,10'd138};
ram[36797] = {-9'd59,10'd141};
ram[36798] = {-9'd56,10'd144};
ram[36799] = {-9'd53,10'd147};
ram[36800] = {-9'd50,10'd150};
ram[36801] = {-9'd47,10'd153};
ram[36802] = {-9'd44,10'd157};
ram[36803] = {-9'd41,10'd160};
ram[36804] = {-9'd37,10'd163};
ram[36805] = {-9'd34,10'd166};
ram[36806] = {-9'd31,10'd169};
ram[36807] = {-9'd28,10'd172};
ram[36808] = {-9'd25,10'd175};
ram[36809] = {-9'd22,10'd179};
ram[36810] = {-9'd19,10'd182};
ram[36811] = {-9'd15,10'd185};
ram[36812] = {-9'd12,10'd188};
ram[36813] = {-9'd9,10'd191};
ram[36814] = {-9'd6,10'd194};
ram[36815] = {-9'd3,10'd197};
ram[36816] = {9'd0,10'd201};
ram[36817] = {9'd3,10'd204};
ram[36818] = {9'd7,10'd207};
ram[36819] = {9'd10,10'd210};
ram[36820] = {9'd13,10'd213};
ram[36821] = {9'd16,10'd216};
ram[36822] = {9'd19,10'd219};
ram[36823] = {9'd22,10'd223};
ram[36824] = {9'd25,10'd226};
ram[36825] = {9'd29,10'd229};
ram[36826] = {9'd32,10'd232};
ram[36827] = {9'd35,10'd235};
ram[36828] = {9'd38,10'd238};
ram[36829] = {9'd41,10'd241};
ram[36830] = {9'd44,10'd245};
ram[36831] = {9'd47,10'd248};
ram[36832] = {9'd51,10'd251};
ram[36833] = {9'd54,10'd254};
ram[36834] = {9'd57,10'd257};
ram[36835] = {9'd60,10'd260};
ram[36836] = {9'd63,10'd263};
ram[36837] = {9'd66,10'd267};
ram[36838] = {9'd69,10'd270};
ram[36839] = {9'd73,10'd273};
ram[36840] = {9'd76,10'd276};
ram[36841] = {9'd79,10'd279};
ram[36842] = {9'd82,10'd282};
ram[36843] = {9'd85,10'd285};
ram[36844] = {9'd88,10'd289};
ram[36845] = {9'd91,10'd292};
ram[36846] = {9'd95,10'd295};
ram[36847] = {9'd98,10'd298};
ram[36848] = {-9'd99,10'd301};
ram[36849] = {-9'd96,10'd304};
ram[36850] = {-9'd93,10'd307};
ram[36851] = {-9'd90,10'd311};
ram[36852] = {-9'd87,10'd314};
ram[36853] = {-9'd84,10'd317};
ram[36854] = {-9'd81,10'd320};
ram[36855] = {-9'd77,10'd323};
ram[36856] = {-9'd74,10'd326};
ram[36857] = {-9'd71,10'd329};
ram[36858] = {-9'd68,10'd333};
ram[36859] = {-9'd65,10'd336};
ram[36860] = {-9'd62,10'd339};
ram[36861] = {-9'd59,10'd342};
ram[36862] = {-9'd55,10'd345};
ram[36863] = {-9'd52,10'd348};
ram[36864] = {-9'd52,10'd348};
ram[36865] = {-9'd49,10'd351};
ram[36866] = {-9'd46,10'd354};
ram[36867] = {-9'd43,10'd358};
ram[36868] = {-9'd40,10'd361};
ram[36869] = {-9'd37,10'd364};
ram[36870] = {-9'd33,10'd367};
ram[36871] = {-9'd30,10'd370};
ram[36872] = {-9'd27,10'd373};
ram[36873] = {-9'd24,10'd376};
ram[36874] = {-9'd21,10'd380};
ram[36875] = {-9'd18,10'd383};
ram[36876] = {-9'd15,10'd386};
ram[36877] = {-9'd11,10'd389};
ram[36878] = {-9'd8,10'd392};
ram[36879] = {-9'd5,10'd395};
ram[36880] = {-9'd2,10'd398};
ram[36881] = {9'd1,-10'd399};
ram[36882] = {9'd4,-10'd396};
ram[36883] = {9'd7,-10'd393};
ram[36884] = {9'd10,-10'd390};
ram[36885] = {9'd14,-10'd387};
ram[36886] = {9'd17,-10'd384};
ram[36887] = {9'd20,-10'd381};
ram[36888] = {9'd23,-10'd377};
ram[36889] = {9'd26,-10'd374};
ram[36890] = {9'd29,-10'd371};
ram[36891] = {9'd32,-10'd368};
ram[36892] = {9'd36,-10'd365};
ram[36893] = {9'd39,-10'd362};
ram[36894] = {9'd42,-10'd359};
ram[36895] = {9'd45,-10'd355};
ram[36896] = {9'd48,-10'd352};
ram[36897] = {9'd51,-10'd349};
ram[36898] = {9'd54,-10'd346};
ram[36899] = {9'd58,-10'd343};
ram[36900] = {9'd61,-10'd340};
ram[36901] = {9'd64,-10'd337};
ram[36902] = {9'd67,-10'd334};
ram[36903] = {9'd70,-10'd330};
ram[36904] = {9'd73,-10'd327};
ram[36905] = {9'd76,-10'd324};
ram[36906] = {9'd80,-10'd321};
ram[36907] = {9'd83,-10'd318};
ram[36908] = {9'd86,-10'd315};
ram[36909] = {9'd89,-10'd312};
ram[36910] = {9'd92,-10'd308};
ram[36911] = {9'd95,-10'd305};
ram[36912] = {9'd98,-10'd302};
ram[36913] = {-9'd99,-10'd299};
ram[36914] = {-9'd96,-10'd296};
ram[36915] = {-9'd92,-10'd293};
ram[36916] = {-9'd89,-10'd290};
ram[36917] = {-9'd86,-10'd286};
ram[36918] = {-9'd83,-10'd283};
ram[36919] = {-9'd80,-10'd280};
ram[36920] = {-9'd77,-10'd277};
ram[36921] = {-9'd74,-10'd274};
ram[36922] = {-9'd70,-10'd271};
ram[36923] = {-9'd67,-10'd268};
ram[36924] = {-9'd64,-10'd264};
ram[36925] = {-9'd61,-10'd261};
ram[36926] = {-9'd58,-10'd258};
ram[36927] = {-9'd55,-10'd255};
ram[36928] = {-9'd52,-10'd252};
ram[36929] = {-9'd48,-10'd249};
ram[36930] = {-9'd45,-10'd246};
ram[36931] = {-9'd42,-10'd242};
ram[36932] = {-9'd39,-10'd239};
ram[36933] = {-9'd36,-10'd236};
ram[36934] = {-9'd33,-10'd233};
ram[36935] = {-9'd30,-10'd230};
ram[36936] = {-9'd26,-10'd227};
ram[36937] = {-9'd23,-10'd224};
ram[36938] = {-9'd20,-10'd220};
ram[36939] = {-9'd17,-10'd217};
ram[36940] = {-9'd14,-10'd214};
ram[36941] = {-9'd11,-10'd211};
ram[36942] = {-9'd8,-10'd208};
ram[36943] = {-9'd4,-10'd205};
ram[36944] = {-9'd1,-10'd202};
ram[36945] = {9'd2,-10'd198};
ram[36946] = {9'd5,-10'd195};
ram[36947] = {9'd8,-10'd192};
ram[36948] = {9'd11,-10'd189};
ram[36949] = {9'd14,-10'd186};
ram[36950] = {9'd18,-10'd183};
ram[36951] = {9'd21,-10'd180};
ram[36952] = {9'd24,-10'd176};
ram[36953] = {9'd27,-10'd173};
ram[36954] = {9'd30,-10'd170};
ram[36955] = {9'd33,-10'd167};
ram[36956] = {9'd36,-10'd164};
ram[36957] = {9'd40,-10'd161};
ram[36958] = {9'd43,-10'd158};
ram[36959] = {9'd46,-10'd154};
ram[36960] = {9'd49,-10'd151};
ram[36961] = {9'd52,-10'd148};
ram[36962] = {9'd55,-10'd145};
ram[36963] = {9'd58,-10'd142};
ram[36964] = {9'd62,-10'd139};
ram[36965] = {9'd65,-10'd136};
ram[36966] = {9'd68,-10'd132};
ram[36967] = {9'd71,-10'd129};
ram[36968] = {9'd74,-10'd126};
ram[36969] = {9'd77,-10'd123};
ram[36970] = {9'd80,-10'd120};
ram[36971] = {9'd84,-10'd117};
ram[36972] = {9'd87,-10'd114};
ram[36973] = {9'd90,-10'd110};
ram[36974] = {9'd93,-10'd107};
ram[36975] = {9'd96,-10'd104};
ram[36976] = {9'd99,-10'd101};
ram[36977] = {-9'd98,-10'd98};
ram[36978] = {-9'd95,-10'd95};
ram[36979] = {-9'd92,-10'd92};
ram[36980] = {-9'd88,-10'd88};
ram[36981] = {-9'd85,-10'd85};
ram[36982] = {-9'd82,-10'd82};
ram[36983] = {-9'd79,-10'd79};
ram[36984] = {-9'd76,-10'd76};
ram[36985] = {-9'd73,-10'd73};
ram[36986] = {-9'd70,-10'd70};
ram[36987] = {-9'd66,-10'd66};
ram[36988] = {-9'd63,-10'd63};
ram[36989] = {-9'd60,-10'd60};
ram[36990] = {-9'd57,-10'd57};
ram[36991] = {-9'd54,-10'd54};
ram[36992] = {-9'd54,-10'd54};
ram[36993] = {-9'd51,-10'd51};
ram[36994] = {-9'd48,-10'd48};
ram[36995] = {-9'd44,-10'd44};
ram[36996] = {-9'd41,-10'd41};
ram[36997] = {-9'd38,-10'd38};
ram[36998] = {-9'd35,-10'd35};
ram[36999] = {-9'd32,-10'd32};
ram[37000] = {-9'd29,-10'd29};
ram[37001] = {-9'd26,-10'd26};
ram[37002] = {-9'd22,-10'd22};
ram[37003] = {-9'd19,-10'd19};
ram[37004] = {-9'd16,-10'd16};
ram[37005] = {-9'd13,-10'd13};
ram[37006] = {-9'd10,-10'd10};
ram[37007] = {-9'd7,-10'd7};
ram[37008] = {-9'd4,-10'd4};
ram[37009] = {9'd0,10'd0};
ram[37010] = {9'd3,10'd3};
ram[37011] = {9'd6,10'd6};
ram[37012] = {9'd9,10'd9};
ram[37013] = {9'd12,10'd12};
ram[37014] = {9'd15,10'd15};
ram[37015] = {9'd18,10'd18};
ram[37016] = {9'd21,10'd21};
ram[37017] = {9'd25,10'd25};
ram[37018] = {9'd28,10'd28};
ram[37019] = {9'd31,10'd31};
ram[37020] = {9'd34,10'd34};
ram[37021] = {9'd37,10'd37};
ram[37022] = {9'd40,10'd40};
ram[37023] = {9'd43,10'd43};
ram[37024] = {9'd47,10'd47};
ram[37025] = {9'd50,10'd50};
ram[37026] = {9'd53,10'd53};
ram[37027] = {9'd56,10'd56};
ram[37028] = {9'd59,10'd59};
ram[37029] = {9'd62,10'd62};
ram[37030] = {9'd65,10'd65};
ram[37031] = {9'd69,10'd69};
ram[37032] = {9'd72,10'd72};
ram[37033] = {9'd75,10'd75};
ram[37034] = {9'd78,10'd78};
ram[37035] = {9'd81,10'd81};
ram[37036] = {9'd84,10'd84};
ram[37037] = {9'd87,10'd87};
ram[37038] = {9'd91,10'd91};
ram[37039] = {9'd94,10'd94};
ram[37040] = {9'd97,10'd97};
ram[37041] = {-9'd100,10'd100};
ram[37042] = {-9'd97,10'd103};
ram[37043] = {-9'd94,10'd106};
ram[37044] = {-9'd91,10'd109};
ram[37045] = {-9'd88,10'd113};
ram[37046] = {-9'd85,10'd116};
ram[37047] = {-9'd81,10'd119};
ram[37048] = {-9'd78,10'd122};
ram[37049] = {-9'd75,10'd125};
ram[37050] = {-9'd72,10'd128};
ram[37051] = {-9'd69,10'd131};
ram[37052] = {-9'd66,10'd135};
ram[37053] = {-9'd63,10'd138};
ram[37054] = {-9'd59,10'd141};
ram[37055] = {-9'd56,10'd144};
ram[37056] = {-9'd53,10'd147};
ram[37057] = {-9'd50,10'd150};
ram[37058] = {-9'd47,10'd153};
ram[37059] = {-9'd44,10'd157};
ram[37060] = {-9'd41,10'd160};
ram[37061] = {-9'd37,10'd163};
ram[37062] = {-9'd34,10'd166};
ram[37063] = {-9'd31,10'd169};
ram[37064] = {-9'd28,10'd172};
ram[37065] = {-9'd25,10'd175};
ram[37066] = {-9'd22,10'd179};
ram[37067] = {-9'd19,10'd182};
ram[37068] = {-9'd15,10'd185};
ram[37069] = {-9'd12,10'd188};
ram[37070] = {-9'd9,10'd191};
ram[37071] = {-9'd6,10'd194};
ram[37072] = {-9'd3,10'd197};
ram[37073] = {9'd0,10'd201};
ram[37074] = {9'd3,10'd204};
ram[37075] = {9'd7,10'd207};
ram[37076] = {9'd10,10'd210};
ram[37077] = {9'd13,10'd213};
ram[37078] = {9'd16,10'd216};
ram[37079] = {9'd19,10'd219};
ram[37080] = {9'd22,10'd223};
ram[37081] = {9'd25,10'd226};
ram[37082] = {9'd29,10'd229};
ram[37083] = {9'd32,10'd232};
ram[37084] = {9'd35,10'd235};
ram[37085] = {9'd38,10'd238};
ram[37086] = {9'd41,10'd241};
ram[37087] = {9'd44,10'd245};
ram[37088] = {9'd47,10'd248};
ram[37089] = {9'd51,10'd251};
ram[37090] = {9'd54,10'd254};
ram[37091] = {9'd57,10'd257};
ram[37092] = {9'd60,10'd260};
ram[37093] = {9'd63,10'd263};
ram[37094] = {9'd66,10'd267};
ram[37095] = {9'd69,10'd270};
ram[37096] = {9'd73,10'd273};
ram[37097] = {9'd76,10'd276};
ram[37098] = {9'd79,10'd279};
ram[37099] = {9'd82,10'd282};
ram[37100] = {9'd85,10'd285};
ram[37101] = {9'd88,10'd289};
ram[37102] = {9'd91,10'd292};
ram[37103] = {9'd95,10'd295};
ram[37104] = {9'd98,10'd298};
ram[37105] = {-9'd99,10'd301};
ram[37106] = {-9'd96,10'd304};
ram[37107] = {-9'd93,10'd307};
ram[37108] = {-9'd90,10'd311};
ram[37109] = {-9'd87,10'd314};
ram[37110] = {-9'd84,10'd317};
ram[37111] = {-9'd81,10'd320};
ram[37112] = {-9'd77,10'd323};
ram[37113] = {-9'd74,10'd326};
ram[37114] = {-9'd71,10'd329};
ram[37115] = {-9'd68,10'd333};
ram[37116] = {-9'd65,10'd336};
ram[37117] = {-9'd62,10'd339};
ram[37118] = {-9'd59,10'd342};
ram[37119] = {-9'd55,10'd345};
ram[37120] = {-9'd55,10'd345};
ram[37121] = {-9'd52,10'd348};
ram[37122] = {-9'd49,10'd351};
ram[37123] = {-9'd46,10'd354};
ram[37124] = {-9'd43,10'd358};
ram[37125] = {-9'd40,10'd361};
ram[37126] = {-9'd37,10'd364};
ram[37127] = {-9'd33,10'd367};
ram[37128] = {-9'd30,10'd370};
ram[37129] = {-9'd27,10'd373};
ram[37130] = {-9'd24,10'd376};
ram[37131] = {-9'd21,10'd380};
ram[37132] = {-9'd18,10'd383};
ram[37133] = {-9'd15,10'd386};
ram[37134] = {-9'd11,10'd389};
ram[37135] = {-9'd8,10'd392};
ram[37136] = {-9'd5,10'd395};
ram[37137] = {-9'd2,10'd398};
ram[37138] = {9'd1,-10'd399};
ram[37139] = {9'd4,-10'd396};
ram[37140] = {9'd7,-10'd393};
ram[37141] = {9'd10,-10'd390};
ram[37142] = {9'd14,-10'd387};
ram[37143] = {9'd17,-10'd384};
ram[37144] = {9'd20,-10'd381};
ram[37145] = {9'd23,-10'd377};
ram[37146] = {9'd26,-10'd374};
ram[37147] = {9'd29,-10'd371};
ram[37148] = {9'd32,-10'd368};
ram[37149] = {9'd36,-10'd365};
ram[37150] = {9'd39,-10'd362};
ram[37151] = {9'd42,-10'd359};
ram[37152] = {9'd45,-10'd355};
ram[37153] = {9'd48,-10'd352};
ram[37154] = {9'd51,-10'd349};
ram[37155] = {9'd54,-10'd346};
ram[37156] = {9'd58,-10'd343};
ram[37157] = {9'd61,-10'd340};
ram[37158] = {9'd64,-10'd337};
ram[37159] = {9'd67,-10'd334};
ram[37160] = {9'd70,-10'd330};
ram[37161] = {9'd73,-10'd327};
ram[37162] = {9'd76,-10'd324};
ram[37163] = {9'd80,-10'd321};
ram[37164] = {9'd83,-10'd318};
ram[37165] = {9'd86,-10'd315};
ram[37166] = {9'd89,-10'd312};
ram[37167] = {9'd92,-10'd308};
ram[37168] = {9'd95,-10'd305};
ram[37169] = {9'd98,-10'd302};
ram[37170] = {-9'd99,-10'd299};
ram[37171] = {-9'd96,-10'd296};
ram[37172] = {-9'd92,-10'd293};
ram[37173] = {-9'd89,-10'd290};
ram[37174] = {-9'd86,-10'd286};
ram[37175] = {-9'd83,-10'd283};
ram[37176] = {-9'd80,-10'd280};
ram[37177] = {-9'd77,-10'd277};
ram[37178] = {-9'd74,-10'd274};
ram[37179] = {-9'd70,-10'd271};
ram[37180] = {-9'd67,-10'd268};
ram[37181] = {-9'd64,-10'd264};
ram[37182] = {-9'd61,-10'd261};
ram[37183] = {-9'd58,-10'd258};
ram[37184] = {-9'd55,-10'd255};
ram[37185] = {-9'd52,-10'd252};
ram[37186] = {-9'd48,-10'd249};
ram[37187] = {-9'd45,-10'd246};
ram[37188] = {-9'd42,-10'd242};
ram[37189] = {-9'd39,-10'd239};
ram[37190] = {-9'd36,-10'd236};
ram[37191] = {-9'd33,-10'd233};
ram[37192] = {-9'd30,-10'd230};
ram[37193] = {-9'd26,-10'd227};
ram[37194] = {-9'd23,-10'd224};
ram[37195] = {-9'd20,-10'd220};
ram[37196] = {-9'd17,-10'd217};
ram[37197] = {-9'd14,-10'd214};
ram[37198] = {-9'd11,-10'd211};
ram[37199] = {-9'd8,-10'd208};
ram[37200] = {-9'd4,-10'd205};
ram[37201] = {-9'd1,-10'd202};
ram[37202] = {9'd2,-10'd198};
ram[37203] = {9'd5,-10'd195};
ram[37204] = {9'd8,-10'd192};
ram[37205] = {9'd11,-10'd189};
ram[37206] = {9'd14,-10'd186};
ram[37207] = {9'd18,-10'd183};
ram[37208] = {9'd21,-10'd180};
ram[37209] = {9'd24,-10'd176};
ram[37210] = {9'd27,-10'd173};
ram[37211] = {9'd30,-10'd170};
ram[37212] = {9'd33,-10'd167};
ram[37213] = {9'd36,-10'd164};
ram[37214] = {9'd40,-10'd161};
ram[37215] = {9'd43,-10'd158};
ram[37216] = {9'd46,-10'd154};
ram[37217] = {9'd49,-10'd151};
ram[37218] = {9'd52,-10'd148};
ram[37219] = {9'd55,-10'd145};
ram[37220] = {9'd58,-10'd142};
ram[37221] = {9'd62,-10'd139};
ram[37222] = {9'd65,-10'd136};
ram[37223] = {9'd68,-10'd132};
ram[37224] = {9'd71,-10'd129};
ram[37225] = {9'd74,-10'd126};
ram[37226] = {9'd77,-10'd123};
ram[37227] = {9'd80,-10'd120};
ram[37228] = {9'd84,-10'd117};
ram[37229] = {9'd87,-10'd114};
ram[37230] = {9'd90,-10'd110};
ram[37231] = {9'd93,-10'd107};
ram[37232] = {9'd96,-10'd104};
ram[37233] = {9'd99,-10'd101};
ram[37234] = {-9'd98,-10'd98};
ram[37235] = {-9'd95,-10'd95};
ram[37236] = {-9'd92,-10'd92};
ram[37237] = {-9'd88,-10'd88};
ram[37238] = {-9'd85,-10'd85};
ram[37239] = {-9'd82,-10'd82};
ram[37240] = {-9'd79,-10'd79};
ram[37241] = {-9'd76,-10'd76};
ram[37242] = {-9'd73,-10'd73};
ram[37243] = {-9'd70,-10'd70};
ram[37244] = {-9'd66,-10'd66};
ram[37245] = {-9'd63,-10'd63};
ram[37246] = {-9'd60,-10'd60};
ram[37247] = {-9'd57,-10'd57};
ram[37248] = {-9'd57,-10'd57};
ram[37249] = {-9'd54,-10'd54};
ram[37250] = {-9'd51,-10'd51};
ram[37251] = {-9'd48,-10'd48};
ram[37252] = {-9'd44,-10'd44};
ram[37253] = {-9'd41,-10'd41};
ram[37254] = {-9'd38,-10'd38};
ram[37255] = {-9'd35,-10'd35};
ram[37256] = {-9'd32,-10'd32};
ram[37257] = {-9'd29,-10'd29};
ram[37258] = {-9'd26,-10'd26};
ram[37259] = {-9'd22,-10'd22};
ram[37260] = {-9'd19,-10'd19};
ram[37261] = {-9'd16,-10'd16};
ram[37262] = {-9'd13,-10'd13};
ram[37263] = {-9'd10,-10'd10};
ram[37264] = {-9'd7,-10'd7};
ram[37265] = {-9'd4,-10'd4};
ram[37266] = {9'd0,10'd0};
ram[37267] = {9'd3,10'd3};
ram[37268] = {9'd6,10'd6};
ram[37269] = {9'd9,10'd9};
ram[37270] = {9'd12,10'd12};
ram[37271] = {9'd15,10'd15};
ram[37272] = {9'd18,10'd18};
ram[37273] = {9'd21,10'd21};
ram[37274] = {9'd25,10'd25};
ram[37275] = {9'd28,10'd28};
ram[37276] = {9'd31,10'd31};
ram[37277] = {9'd34,10'd34};
ram[37278] = {9'd37,10'd37};
ram[37279] = {9'd40,10'd40};
ram[37280] = {9'd43,10'd43};
ram[37281] = {9'd47,10'd47};
ram[37282] = {9'd50,10'd50};
ram[37283] = {9'd53,10'd53};
ram[37284] = {9'd56,10'd56};
ram[37285] = {9'd59,10'd59};
ram[37286] = {9'd62,10'd62};
ram[37287] = {9'd65,10'd65};
ram[37288] = {9'd69,10'd69};
ram[37289] = {9'd72,10'd72};
ram[37290] = {9'd75,10'd75};
ram[37291] = {9'd78,10'd78};
ram[37292] = {9'd81,10'd81};
ram[37293] = {9'd84,10'd84};
ram[37294] = {9'd87,10'd87};
ram[37295] = {9'd91,10'd91};
ram[37296] = {9'd94,10'd94};
ram[37297] = {9'd97,10'd97};
ram[37298] = {-9'd100,10'd100};
ram[37299] = {-9'd97,10'd103};
ram[37300] = {-9'd94,10'd106};
ram[37301] = {-9'd91,10'd109};
ram[37302] = {-9'd88,10'd113};
ram[37303] = {-9'd85,10'd116};
ram[37304] = {-9'd81,10'd119};
ram[37305] = {-9'd78,10'd122};
ram[37306] = {-9'd75,10'd125};
ram[37307] = {-9'd72,10'd128};
ram[37308] = {-9'd69,10'd131};
ram[37309] = {-9'd66,10'd135};
ram[37310] = {-9'd63,10'd138};
ram[37311] = {-9'd59,10'd141};
ram[37312] = {-9'd56,10'd144};
ram[37313] = {-9'd53,10'd147};
ram[37314] = {-9'd50,10'd150};
ram[37315] = {-9'd47,10'd153};
ram[37316] = {-9'd44,10'd157};
ram[37317] = {-9'd41,10'd160};
ram[37318] = {-9'd37,10'd163};
ram[37319] = {-9'd34,10'd166};
ram[37320] = {-9'd31,10'd169};
ram[37321] = {-9'd28,10'd172};
ram[37322] = {-9'd25,10'd175};
ram[37323] = {-9'd22,10'd179};
ram[37324] = {-9'd19,10'd182};
ram[37325] = {-9'd15,10'd185};
ram[37326] = {-9'd12,10'd188};
ram[37327] = {-9'd9,10'd191};
ram[37328] = {-9'd6,10'd194};
ram[37329] = {-9'd3,10'd197};
ram[37330] = {9'd0,10'd201};
ram[37331] = {9'd3,10'd204};
ram[37332] = {9'd7,10'd207};
ram[37333] = {9'd10,10'd210};
ram[37334] = {9'd13,10'd213};
ram[37335] = {9'd16,10'd216};
ram[37336] = {9'd19,10'd219};
ram[37337] = {9'd22,10'd223};
ram[37338] = {9'd25,10'd226};
ram[37339] = {9'd29,10'd229};
ram[37340] = {9'd32,10'd232};
ram[37341] = {9'd35,10'd235};
ram[37342] = {9'd38,10'd238};
ram[37343] = {9'd41,10'd241};
ram[37344] = {9'd44,10'd245};
ram[37345] = {9'd47,10'd248};
ram[37346] = {9'd51,10'd251};
ram[37347] = {9'd54,10'd254};
ram[37348] = {9'd57,10'd257};
ram[37349] = {9'd60,10'd260};
ram[37350] = {9'd63,10'd263};
ram[37351] = {9'd66,10'd267};
ram[37352] = {9'd69,10'd270};
ram[37353] = {9'd73,10'd273};
ram[37354] = {9'd76,10'd276};
ram[37355] = {9'd79,10'd279};
ram[37356] = {9'd82,10'd282};
ram[37357] = {9'd85,10'd285};
ram[37358] = {9'd88,10'd289};
ram[37359] = {9'd91,10'd292};
ram[37360] = {9'd95,10'd295};
ram[37361] = {9'd98,10'd298};
ram[37362] = {-9'd99,10'd301};
ram[37363] = {-9'd96,10'd304};
ram[37364] = {-9'd93,10'd307};
ram[37365] = {-9'd90,10'd311};
ram[37366] = {-9'd87,10'd314};
ram[37367] = {-9'd84,10'd317};
ram[37368] = {-9'd81,10'd320};
ram[37369] = {-9'd77,10'd323};
ram[37370] = {-9'd74,10'd326};
ram[37371] = {-9'd71,10'd329};
ram[37372] = {-9'd68,10'd333};
ram[37373] = {-9'd65,10'd336};
ram[37374] = {-9'd62,10'd339};
ram[37375] = {-9'd59,10'd342};
ram[37376] = {-9'd59,10'd342};
ram[37377] = {-9'd55,10'd345};
ram[37378] = {-9'd52,10'd348};
ram[37379] = {-9'd49,10'd351};
ram[37380] = {-9'd46,10'd354};
ram[37381] = {-9'd43,10'd358};
ram[37382] = {-9'd40,10'd361};
ram[37383] = {-9'd37,10'd364};
ram[37384] = {-9'd33,10'd367};
ram[37385] = {-9'd30,10'd370};
ram[37386] = {-9'd27,10'd373};
ram[37387] = {-9'd24,10'd376};
ram[37388] = {-9'd21,10'd380};
ram[37389] = {-9'd18,10'd383};
ram[37390] = {-9'd15,10'd386};
ram[37391] = {-9'd11,10'd389};
ram[37392] = {-9'd8,10'd392};
ram[37393] = {-9'd5,10'd395};
ram[37394] = {-9'd2,10'd398};
ram[37395] = {9'd1,-10'd399};
ram[37396] = {9'd4,-10'd396};
ram[37397] = {9'd7,-10'd393};
ram[37398] = {9'd10,-10'd390};
ram[37399] = {9'd14,-10'd387};
ram[37400] = {9'd17,-10'd384};
ram[37401] = {9'd20,-10'd381};
ram[37402] = {9'd23,-10'd377};
ram[37403] = {9'd26,-10'd374};
ram[37404] = {9'd29,-10'd371};
ram[37405] = {9'd32,-10'd368};
ram[37406] = {9'd36,-10'd365};
ram[37407] = {9'd39,-10'd362};
ram[37408] = {9'd42,-10'd359};
ram[37409] = {9'd45,-10'd355};
ram[37410] = {9'd48,-10'd352};
ram[37411] = {9'd51,-10'd349};
ram[37412] = {9'd54,-10'd346};
ram[37413] = {9'd58,-10'd343};
ram[37414] = {9'd61,-10'd340};
ram[37415] = {9'd64,-10'd337};
ram[37416] = {9'd67,-10'd334};
ram[37417] = {9'd70,-10'd330};
ram[37418] = {9'd73,-10'd327};
ram[37419] = {9'd76,-10'd324};
ram[37420] = {9'd80,-10'd321};
ram[37421] = {9'd83,-10'd318};
ram[37422] = {9'd86,-10'd315};
ram[37423] = {9'd89,-10'd312};
ram[37424] = {9'd92,-10'd308};
ram[37425] = {9'd95,-10'd305};
ram[37426] = {9'd98,-10'd302};
ram[37427] = {-9'd99,-10'd299};
ram[37428] = {-9'd96,-10'd296};
ram[37429] = {-9'd92,-10'd293};
ram[37430] = {-9'd89,-10'd290};
ram[37431] = {-9'd86,-10'd286};
ram[37432] = {-9'd83,-10'd283};
ram[37433] = {-9'd80,-10'd280};
ram[37434] = {-9'd77,-10'd277};
ram[37435] = {-9'd74,-10'd274};
ram[37436] = {-9'd70,-10'd271};
ram[37437] = {-9'd67,-10'd268};
ram[37438] = {-9'd64,-10'd264};
ram[37439] = {-9'd61,-10'd261};
ram[37440] = {-9'd58,-10'd258};
ram[37441] = {-9'd55,-10'd255};
ram[37442] = {-9'd52,-10'd252};
ram[37443] = {-9'd48,-10'd249};
ram[37444] = {-9'd45,-10'd246};
ram[37445] = {-9'd42,-10'd242};
ram[37446] = {-9'd39,-10'd239};
ram[37447] = {-9'd36,-10'd236};
ram[37448] = {-9'd33,-10'd233};
ram[37449] = {-9'd30,-10'd230};
ram[37450] = {-9'd26,-10'd227};
ram[37451] = {-9'd23,-10'd224};
ram[37452] = {-9'd20,-10'd220};
ram[37453] = {-9'd17,-10'd217};
ram[37454] = {-9'd14,-10'd214};
ram[37455] = {-9'd11,-10'd211};
ram[37456] = {-9'd8,-10'd208};
ram[37457] = {-9'd4,-10'd205};
ram[37458] = {-9'd1,-10'd202};
ram[37459] = {9'd2,-10'd198};
ram[37460] = {9'd5,-10'd195};
ram[37461] = {9'd8,-10'd192};
ram[37462] = {9'd11,-10'd189};
ram[37463] = {9'd14,-10'd186};
ram[37464] = {9'd18,-10'd183};
ram[37465] = {9'd21,-10'd180};
ram[37466] = {9'd24,-10'd176};
ram[37467] = {9'd27,-10'd173};
ram[37468] = {9'd30,-10'd170};
ram[37469] = {9'd33,-10'd167};
ram[37470] = {9'd36,-10'd164};
ram[37471] = {9'd40,-10'd161};
ram[37472] = {9'd43,-10'd158};
ram[37473] = {9'd46,-10'd154};
ram[37474] = {9'd49,-10'd151};
ram[37475] = {9'd52,-10'd148};
ram[37476] = {9'd55,-10'd145};
ram[37477] = {9'd58,-10'd142};
ram[37478] = {9'd62,-10'd139};
ram[37479] = {9'd65,-10'd136};
ram[37480] = {9'd68,-10'd132};
ram[37481] = {9'd71,-10'd129};
ram[37482] = {9'd74,-10'd126};
ram[37483] = {9'd77,-10'd123};
ram[37484] = {9'd80,-10'd120};
ram[37485] = {9'd84,-10'd117};
ram[37486] = {9'd87,-10'd114};
ram[37487] = {9'd90,-10'd110};
ram[37488] = {9'd93,-10'd107};
ram[37489] = {9'd96,-10'd104};
ram[37490] = {9'd99,-10'd101};
ram[37491] = {-9'd98,-10'd98};
ram[37492] = {-9'd95,-10'd95};
ram[37493] = {-9'd92,-10'd92};
ram[37494] = {-9'd88,-10'd88};
ram[37495] = {-9'd85,-10'd85};
ram[37496] = {-9'd82,-10'd82};
ram[37497] = {-9'd79,-10'd79};
ram[37498] = {-9'd76,-10'd76};
ram[37499] = {-9'd73,-10'd73};
ram[37500] = {-9'd70,-10'd70};
ram[37501] = {-9'd66,-10'd66};
ram[37502] = {-9'd63,-10'd63};
ram[37503] = {-9'd60,-10'd60};
ram[37504] = {-9'd60,-10'd60};
ram[37505] = {-9'd57,-10'd57};
ram[37506] = {-9'd54,-10'd54};
ram[37507] = {-9'd51,-10'd51};
ram[37508] = {-9'd48,-10'd48};
ram[37509] = {-9'd44,-10'd44};
ram[37510] = {-9'd41,-10'd41};
ram[37511] = {-9'd38,-10'd38};
ram[37512] = {-9'd35,-10'd35};
ram[37513] = {-9'd32,-10'd32};
ram[37514] = {-9'd29,-10'd29};
ram[37515] = {-9'd26,-10'd26};
ram[37516] = {-9'd22,-10'd22};
ram[37517] = {-9'd19,-10'd19};
ram[37518] = {-9'd16,-10'd16};
ram[37519] = {-9'd13,-10'd13};
ram[37520] = {-9'd10,-10'd10};
ram[37521] = {-9'd7,-10'd7};
ram[37522] = {-9'd4,-10'd4};
ram[37523] = {9'd0,10'd0};
ram[37524] = {9'd3,10'd3};
ram[37525] = {9'd6,10'd6};
ram[37526] = {9'd9,10'd9};
ram[37527] = {9'd12,10'd12};
ram[37528] = {9'd15,10'd15};
ram[37529] = {9'd18,10'd18};
ram[37530] = {9'd21,10'd21};
ram[37531] = {9'd25,10'd25};
ram[37532] = {9'd28,10'd28};
ram[37533] = {9'd31,10'd31};
ram[37534] = {9'd34,10'd34};
ram[37535] = {9'd37,10'd37};
ram[37536] = {9'd40,10'd40};
ram[37537] = {9'd43,10'd43};
ram[37538] = {9'd47,10'd47};
ram[37539] = {9'd50,10'd50};
ram[37540] = {9'd53,10'd53};
ram[37541] = {9'd56,10'd56};
ram[37542] = {9'd59,10'd59};
ram[37543] = {9'd62,10'd62};
ram[37544] = {9'd65,10'd65};
ram[37545] = {9'd69,10'd69};
ram[37546] = {9'd72,10'd72};
ram[37547] = {9'd75,10'd75};
ram[37548] = {9'd78,10'd78};
ram[37549] = {9'd81,10'd81};
ram[37550] = {9'd84,10'd84};
ram[37551] = {9'd87,10'd87};
ram[37552] = {9'd91,10'd91};
ram[37553] = {9'd94,10'd94};
ram[37554] = {9'd97,10'd97};
ram[37555] = {-9'd100,10'd100};
ram[37556] = {-9'd97,10'd103};
ram[37557] = {-9'd94,10'd106};
ram[37558] = {-9'd91,10'd109};
ram[37559] = {-9'd88,10'd113};
ram[37560] = {-9'd85,10'd116};
ram[37561] = {-9'd81,10'd119};
ram[37562] = {-9'd78,10'd122};
ram[37563] = {-9'd75,10'd125};
ram[37564] = {-9'd72,10'd128};
ram[37565] = {-9'd69,10'd131};
ram[37566] = {-9'd66,10'd135};
ram[37567] = {-9'd63,10'd138};
ram[37568] = {-9'd59,10'd141};
ram[37569] = {-9'd56,10'd144};
ram[37570] = {-9'd53,10'd147};
ram[37571] = {-9'd50,10'd150};
ram[37572] = {-9'd47,10'd153};
ram[37573] = {-9'd44,10'd157};
ram[37574] = {-9'd41,10'd160};
ram[37575] = {-9'd37,10'd163};
ram[37576] = {-9'd34,10'd166};
ram[37577] = {-9'd31,10'd169};
ram[37578] = {-9'd28,10'd172};
ram[37579] = {-9'd25,10'd175};
ram[37580] = {-9'd22,10'd179};
ram[37581] = {-9'd19,10'd182};
ram[37582] = {-9'd15,10'd185};
ram[37583] = {-9'd12,10'd188};
ram[37584] = {-9'd9,10'd191};
ram[37585] = {-9'd6,10'd194};
ram[37586] = {-9'd3,10'd197};
ram[37587] = {9'd0,10'd201};
ram[37588] = {9'd3,10'd204};
ram[37589] = {9'd7,10'd207};
ram[37590] = {9'd10,10'd210};
ram[37591] = {9'd13,10'd213};
ram[37592] = {9'd16,10'd216};
ram[37593] = {9'd19,10'd219};
ram[37594] = {9'd22,10'd223};
ram[37595] = {9'd25,10'd226};
ram[37596] = {9'd29,10'd229};
ram[37597] = {9'd32,10'd232};
ram[37598] = {9'd35,10'd235};
ram[37599] = {9'd38,10'd238};
ram[37600] = {9'd41,10'd241};
ram[37601] = {9'd44,10'd245};
ram[37602] = {9'd47,10'd248};
ram[37603] = {9'd51,10'd251};
ram[37604] = {9'd54,10'd254};
ram[37605] = {9'd57,10'd257};
ram[37606] = {9'd60,10'd260};
ram[37607] = {9'd63,10'd263};
ram[37608] = {9'd66,10'd267};
ram[37609] = {9'd69,10'd270};
ram[37610] = {9'd73,10'd273};
ram[37611] = {9'd76,10'd276};
ram[37612] = {9'd79,10'd279};
ram[37613] = {9'd82,10'd282};
ram[37614] = {9'd85,10'd285};
ram[37615] = {9'd88,10'd289};
ram[37616] = {9'd91,10'd292};
ram[37617] = {9'd95,10'd295};
ram[37618] = {9'd98,10'd298};
ram[37619] = {-9'd99,10'd301};
ram[37620] = {-9'd96,10'd304};
ram[37621] = {-9'd93,10'd307};
ram[37622] = {-9'd90,10'd311};
ram[37623] = {-9'd87,10'd314};
ram[37624] = {-9'd84,10'd317};
ram[37625] = {-9'd81,10'd320};
ram[37626] = {-9'd77,10'd323};
ram[37627] = {-9'd74,10'd326};
ram[37628] = {-9'd71,10'd329};
ram[37629] = {-9'd68,10'd333};
ram[37630] = {-9'd65,10'd336};
ram[37631] = {-9'd62,10'd339};
ram[37632] = {-9'd62,10'd339};
ram[37633] = {-9'd59,10'd342};
ram[37634] = {-9'd55,10'd345};
ram[37635] = {-9'd52,10'd348};
ram[37636] = {-9'd49,10'd351};
ram[37637] = {-9'd46,10'd354};
ram[37638] = {-9'd43,10'd358};
ram[37639] = {-9'd40,10'd361};
ram[37640] = {-9'd37,10'd364};
ram[37641] = {-9'd33,10'd367};
ram[37642] = {-9'd30,10'd370};
ram[37643] = {-9'd27,10'd373};
ram[37644] = {-9'd24,10'd376};
ram[37645] = {-9'd21,10'd380};
ram[37646] = {-9'd18,10'd383};
ram[37647] = {-9'd15,10'd386};
ram[37648] = {-9'd11,10'd389};
ram[37649] = {-9'd8,10'd392};
ram[37650] = {-9'd5,10'd395};
ram[37651] = {-9'd2,10'd398};
ram[37652] = {9'd1,-10'd399};
ram[37653] = {9'd4,-10'd396};
ram[37654] = {9'd7,-10'd393};
ram[37655] = {9'd10,-10'd390};
ram[37656] = {9'd14,-10'd387};
ram[37657] = {9'd17,-10'd384};
ram[37658] = {9'd20,-10'd381};
ram[37659] = {9'd23,-10'd377};
ram[37660] = {9'd26,-10'd374};
ram[37661] = {9'd29,-10'd371};
ram[37662] = {9'd32,-10'd368};
ram[37663] = {9'd36,-10'd365};
ram[37664] = {9'd39,-10'd362};
ram[37665] = {9'd42,-10'd359};
ram[37666] = {9'd45,-10'd355};
ram[37667] = {9'd48,-10'd352};
ram[37668] = {9'd51,-10'd349};
ram[37669] = {9'd54,-10'd346};
ram[37670] = {9'd58,-10'd343};
ram[37671] = {9'd61,-10'd340};
ram[37672] = {9'd64,-10'd337};
ram[37673] = {9'd67,-10'd334};
ram[37674] = {9'd70,-10'd330};
ram[37675] = {9'd73,-10'd327};
ram[37676] = {9'd76,-10'd324};
ram[37677] = {9'd80,-10'd321};
ram[37678] = {9'd83,-10'd318};
ram[37679] = {9'd86,-10'd315};
ram[37680] = {9'd89,-10'd312};
ram[37681] = {9'd92,-10'd308};
ram[37682] = {9'd95,-10'd305};
ram[37683] = {9'd98,-10'd302};
ram[37684] = {-9'd99,-10'd299};
ram[37685] = {-9'd96,-10'd296};
ram[37686] = {-9'd92,-10'd293};
ram[37687] = {-9'd89,-10'd290};
ram[37688] = {-9'd86,-10'd286};
ram[37689] = {-9'd83,-10'd283};
ram[37690] = {-9'd80,-10'd280};
ram[37691] = {-9'd77,-10'd277};
ram[37692] = {-9'd74,-10'd274};
ram[37693] = {-9'd70,-10'd271};
ram[37694] = {-9'd67,-10'd268};
ram[37695] = {-9'd64,-10'd264};
ram[37696] = {-9'd61,-10'd261};
ram[37697] = {-9'd58,-10'd258};
ram[37698] = {-9'd55,-10'd255};
ram[37699] = {-9'd52,-10'd252};
ram[37700] = {-9'd48,-10'd249};
ram[37701] = {-9'd45,-10'd246};
ram[37702] = {-9'd42,-10'd242};
ram[37703] = {-9'd39,-10'd239};
ram[37704] = {-9'd36,-10'd236};
ram[37705] = {-9'd33,-10'd233};
ram[37706] = {-9'd30,-10'd230};
ram[37707] = {-9'd26,-10'd227};
ram[37708] = {-9'd23,-10'd224};
ram[37709] = {-9'd20,-10'd220};
ram[37710] = {-9'd17,-10'd217};
ram[37711] = {-9'd14,-10'd214};
ram[37712] = {-9'd11,-10'd211};
ram[37713] = {-9'd8,-10'd208};
ram[37714] = {-9'd4,-10'd205};
ram[37715] = {-9'd1,-10'd202};
ram[37716] = {9'd2,-10'd198};
ram[37717] = {9'd5,-10'd195};
ram[37718] = {9'd8,-10'd192};
ram[37719] = {9'd11,-10'd189};
ram[37720] = {9'd14,-10'd186};
ram[37721] = {9'd18,-10'd183};
ram[37722] = {9'd21,-10'd180};
ram[37723] = {9'd24,-10'd176};
ram[37724] = {9'd27,-10'd173};
ram[37725] = {9'd30,-10'd170};
ram[37726] = {9'd33,-10'd167};
ram[37727] = {9'd36,-10'd164};
ram[37728] = {9'd40,-10'd161};
ram[37729] = {9'd43,-10'd158};
ram[37730] = {9'd46,-10'd154};
ram[37731] = {9'd49,-10'd151};
ram[37732] = {9'd52,-10'd148};
ram[37733] = {9'd55,-10'd145};
ram[37734] = {9'd58,-10'd142};
ram[37735] = {9'd62,-10'd139};
ram[37736] = {9'd65,-10'd136};
ram[37737] = {9'd68,-10'd132};
ram[37738] = {9'd71,-10'd129};
ram[37739] = {9'd74,-10'd126};
ram[37740] = {9'd77,-10'd123};
ram[37741] = {9'd80,-10'd120};
ram[37742] = {9'd84,-10'd117};
ram[37743] = {9'd87,-10'd114};
ram[37744] = {9'd90,-10'd110};
ram[37745] = {9'd93,-10'd107};
ram[37746] = {9'd96,-10'd104};
ram[37747] = {9'd99,-10'd101};
ram[37748] = {-9'd98,-10'd98};
ram[37749] = {-9'd95,-10'd95};
ram[37750] = {-9'd92,-10'd92};
ram[37751] = {-9'd88,-10'd88};
ram[37752] = {-9'd85,-10'd85};
ram[37753] = {-9'd82,-10'd82};
ram[37754] = {-9'd79,-10'd79};
ram[37755] = {-9'd76,-10'd76};
ram[37756] = {-9'd73,-10'd73};
ram[37757] = {-9'd70,-10'd70};
ram[37758] = {-9'd66,-10'd66};
ram[37759] = {-9'd63,-10'd63};
ram[37760] = {-9'd63,-10'd63};
ram[37761] = {-9'd60,-10'd60};
ram[37762] = {-9'd57,-10'd57};
ram[37763] = {-9'd54,-10'd54};
ram[37764] = {-9'd51,-10'd51};
ram[37765] = {-9'd48,-10'd48};
ram[37766] = {-9'd44,-10'd44};
ram[37767] = {-9'd41,-10'd41};
ram[37768] = {-9'd38,-10'd38};
ram[37769] = {-9'd35,-10'd35};
ram[37770] = {-9'd32,-10'd32};
ram[37771] = {-9'd29,-10'd29};
ram[37772] = {-9'd26,-10'd26};
ram[37773] = {-9'd22,-10'd22};
ram[37774] = {-9'd19,-10'd19};
ram[37775] = {-9'd16,-10'd16};
ram[37776] = {-9'd13,-10'd13};
ram[37777] = {-9'd10,-10'd10};
ram[37778] = {-9'd7,-10'd7};
ram[37779] = {-9'd4,-10'd4};
ram[37780] = {9'd0,10'd0};
ram[37781] = {9'd3,10'd3};
ram[37782] = {9'd6,10'd6};
ram[37783] = {9'd9,10'd9};
ram[37784] = {9'd12,10'd12};
ram[37785] = {9'd15,10'd15};
ram[37786] = {9'd18,10'd18};
ram[37787] = {9'd21,10'd21};
ram[37788] = {9'd25,10'd25};
ram[37789] = {9'd28,10'd28};
ram[37790] = {9'd31,10'd31};
ram[37791] = {9'd34,10'd34};
ram[37792] = {9'd37,10'd37};
ram[37793] = {9'd40,10'd40};
ram[37794] = {9'd43,10'd43};
ram[37795] = {9'd47,10'd47};
ram[37796] = {9'd50,10'd50};
ram[37797] = {9'd53,10'd53};
ram[37798] = {9'd56,10'd56};
ram[37799] = {9'd59,10'd59};
ram[37800] = {9'd62,10'd62};
ram[37801] = {9'd65,10'd65};
ram[37802] = {9'd69,10'd69};
ram[37803] = {9'd72,10'd72};
ram[37804] = {9'd75,10'd75};
ram[37805] = {9'd78,10'd78};
ram[37806] = {9'd81,10'd81};
ram[37807] = {9'd84,10'd84};
ram[37808] = {9'd87,10'd87};
ram[37809] = {9'd91,10'd91};
ram[37810] = {9'd94,10'd94};
ram[37811] = {9'd97,10'd97};
ram[37812] = {-9'd100,10'd100};
ram[37813] = {-9'd97,10'd103};
ram[37814] = {-9'd94,10'd106};
ram[37815] = {-9'd91,10'd109};
ram[37816] = {-9'd88,10'd113};
ram[37817] = {-9'd85,10'd116};
ram[37818] = {-9'd81,10'd119};
ram[37819] = {-9'd78,10'd122};
ram[37820] = {-9'd75,10'd125};
ram[37821] = {-9'd72,10'd128};
ram[37822] = {-9'd69,10'd131};
ram[37823] = {-9'd66,10'd135};
ram[37824] = {-9'd63,10'd138};
ram[37825] = {-9'd59,10'd141};
ram[37826] = {-9'd56,10'd144};
ram[37827] = {-9'd53,10'd147};
ram[37828] = {-9'd50,10'd150};
ram[37829] = {-9'd47,10'd153};
ram[37830] = {-9'd44,10'd157};
ram[37831] = {-9'd41,10'd160};
ram[37832] = {-9'd37,10'd163};
ram[37833] = {-9'd34,10'd166};
ram[37834] = {-9'd31,10'd169};
ram[37835] = {-9'd28,10'd172};
ram[37836] = {-9'd25,10'd175};
ram[37837] = {-9'd22,10'd179};
ram[37838] = {-9'd19,10'd182};
ram[37839] = {-9'd15,10'd185};
ram[37840] = {-9'd12,10'd188};
ram[37841] = {-9'd9,10'd191};
ram[37842] = {-9'd6,10'd194};
ram[37843] = {-9'd3,10'd197};
ram[37844] = {9'd0,10'd201};
ram[37845] = {9'd3,10'd204};
ram[37846] = {9'd7,10'd207};
ram[37847] = {9'd10,10'd210};
ram[37848] = {9'd13,10'd213};
ram[37849] = {9'd16,10'd216};
ram[37850] = {9'd19,10'd219};
ram[37851] = {9'd22,10'd223};
ram[37852] = {9'd25,10'd226};
ram[37853] = {9'd29,10'd229};
ram[37854] = {9'd32,10'd232};
ram[37855] = {9'd35,10'd235};
ram[37856] = {9'd38,10'd238};
ram[37857] = {9'd41,10'd241};
ram[37858] = {9'd44,10'd245};
ram[37859] = {9'd47,10'd248};
ram[37860] = {9'd51,10'd251};
ram[37861] = {9'd54,10'd254};
ram[37862] = {9'd57,10'd257};
ram[37863] = {9'd60,10'd260};
ram[37864] = {9'd63,10'd263};
ram[37865] = {9'd66,10'd267};
ram[37866] = {9'd69,10'd270};
ram[37867] = {9'd73,10'd273};
ram[37868] = {9'd76,10'd276};
ram[37869] = {9'd79,10'd279};
ram[37870] = {9'd82,10'd282};
ram[37871] = {9'd85,10'd285};
ram[37872] = {9'd88,10'd289};
ram[37873] = {9'd91,10'd292};
ram[37874] = {9'd95,10'd295};
ram[37875] = {9'd98,10'd298};
ram[37876] = {-9'd99,10'd301};
ram[37877] = {-9'd96,10'd304};
ram[37878] = {-9'd93,10'd307};
ram[37879] = {-9'd90,10'd311};
ram[37880] = {-9'd87,10'd314};
ram[37881] = {-9'd84,10'd317};
ram[37882] = {-9'd81,10'd320};
ram[37883] = {-9'd77,10'd323};
ram[37884] = {-9'd74,10'd326};
ram[37885] = {-9'd71,10'd329};
ram[37886] = {-9'd68,10'd333};
ram[37887] = {-9'd65,10'd336};
ram[37888] = {-9'd65,10'd336};
ram[37889] = {-9'd62,10'd339};
ram[37890] = {-9'd59,10'd342};
ram[37891] = {-9'd55,10'd345};
ram[37892] = {-9'd52,10'd348};
ram[37893] = {-9'd49,10'd351};
ram[37894] = {-9'd46,10'd354};
ram[37895] = {-9'd43,10'd358};
ram[37896] = {-9'd40,10'd361};
ram[37897] = {-9'd37,10'd364};
ram[37898] = {-9'd33,10'd367};
ram[37899] = {-9'd30,10'd370};
ram[37900] = {-9'd27,10'd373};
ram[37901] = {-9'd24,10'd376};
ram[37902] = {-9'd21,10'd380};
ram[37903] = {-9'd18,10'd383};
ram[37904] = {-9'd15,10'd386};
ram[37905] = {-9'd11,10'd389};
ram[37906] = {-9'd8,10'd392};
ram[37907] = {-9'd5,10'd395};
ram[37908] = {-9'd2,10'd398};
ram[37909] = {9'd1,-10'd399};
ram[37910] = {9'd4,-10'd396};
ram[37911] = {9'd7,-10'd393};
ram[37912] = {9'd10,-10'd390};
ram[37913] = {9'd14,-10'd387};
ram[37914] = {9'd17,-10'd384};
ram[37915] = {9'd20,-10'd381};
ram[37916] = {9'd23,-10'd377};
ram[37917] = {9'd26,-10'd374};
ram[37918] = {9'd29,-10'd371};
ram[37919] = {9'd32,-10'd368};
ram[37920] = {9'd36,-10'd365};
ram[37921] = {9'd39,-10'd362};
ram[37922] = {9'd42,-10'd359};
ram[37923] = {9'd45,-10'd355};
ram[37924] = {9'd48,-10'd352};
ram[37925] = {9'd51,-10'd349};
ram[37926] = {9'd54,-10'd346};
ram[37927] = {9'd58,-10'd343};
ram[37928] = {9'd61,-10'd340};
ram[37929] = {9'd64,-10'd337};
ram[37930] = {9'd67,-10'd334};
ram[37931] = {9'd70,-10'd330};
ram[37932] = {9'd73,-10'd327};
ram[37933] = {9'd76,-10'd324};
ram[37934] = {9'd80,-10'd321};
ram[37935] = {9'd83,-10'd318};
ram[37936] = {9'd86,-10'd315};
ram[37937] = {9'd89,-10'd312};
ram[37938] = {9'd92,-10'd308};
ram[37939] = {9'd95,-10'd305};
ram[37940] = {9'd98,-10'd302};
ram[37941] = {-9'd99,-10'd299};
ram[37942] = {-9'd96,-10'd296};
ram[37943] = {-9'd92,-10'd293};
ram[37944] = {-9'd89,-10'd290};
ram[37945] = {-9'd86,-10'd286};
ram[37946] = {-9'd83,-10'd283};
ram[37947] = {-9'd80,-10'd280};
ram[37948] = {-9'd77,-10'd277};
ram[37949] = {-9'd74,-10'd274};
ram[37950] = {-9'd70,-10'd271};
ram[37951] = {-9'd67,-10'd268};
ram[37952] = {-9'd64,-10'd264};
ram[37953] = {-9'd61,-10'd261};
ram[37954] = {-9'd58,-10'd258};
ram[37955] = {-9'd55,-10'd255};
ram[37956] = {-9'd52,-10'd252};
ram[37957] = {-9'd48,-10'd249};
ram[37958] = {-9'd45,-10'd246};
ram[37959] = {-9'd42,-10'd242};
ram[37960] = {-9'd39,-10'd239};
ram[37961] = {-9'd36,-10'd236};
ram[37962] = {-9'd33,-10'd233};
ram[37963] = {-9'd30,-10'd230};
ram[37964] = {-9'd26,-10'd227};
ram[37965] = {-9'd23,-10'd224};
ram[37966] = {-9'd20,-10'd220};
ram[37967] = {-9'd17,-10'd217};
ram[37968] = {-9'd14,-10'd214};
ram[37969] = {-9'd11,-10'd211};
ram[37970] = {-9'd8,-10'd208};
ram[37971] = {-9'd4,-10'd205};
ram[37972] = {-9'd1,-10'd202};
ram[37973] = {9'd2,-10'd198};
ram[37974] = {9'd5,-10'd195};
ram[37975] = {9'd8,-10'd192};
ram[37976] = {9'd11,-10'd189};
ram[37977] = {9'd14,-10'd186};
ram[37978] = {9'd18,-10'd183};
ram[37979] = {9'd21,-10'd180};
ram[37980] = {9'd24,-10'd176};
ram[37981] = {9'd27,-10'd173};
ram[37982] = {9'd30,-10'd170};
ram[37983] = {9'd33,-10'd167};
ram[37984] = {9'd36,-10'd164};
ram[37985] = {9'd40,-10'd161};
ram[37986] = {9'd43,-10'd158};
ram[37987] = {9'd46,-10'd154};
ram[37988] = {9'd49,-10'd151};
ram[37989] = {9'd52,-10'd148};
ram[37990] = {9'd55,-10'd145};
ram[37991] = {9'd58,-10'd142};
ram[37992] = {9'd62,-10'd139};
ram[37993] = {9'd65,-10'd136};
ram[37994] = {9'd68,-10'd132};
ram[37995] = {9'd71,-10'd129};
ram[37996] = {9'd74,-10'd126};
ram[37997] = {9'd77,-10'd123};
ram[37998] = {9'd80,-10'd120};
ram[37999] = {9'd84,-10'd117};
ram[38000] = {9'd87,-10'd114};
ram[38001] = {9'd90,-10'd110};
ram[38002] = {9'd93,-10'd107};
ram[38003] = {9'd96,-10'd104};
ram[38004] = {9'd99,-10'd101};
ram[38005] = {-9'd98,-10'd98};
ram[38006] = {-9'd95,-10'd95};
ram[38007] = {-9'd92,-10'd92};
ram[38008] = {-9'd88,-10'd88};
ram[38009] = {-9'd85,-10'd85};
ram[38010] = {-9'd82,-10'd82};
ram[38011] = {-9'd79,-10'd79};
ram[38012] = {-9'd76,-10'd76};
ram[38013] = {-9'd73,-10'd73};
ram[38014] = {-9'd70,-10'd70};
ram[38015] = {-9'd66,-10'd66};
ram[38016] = {-9'd66,-10'd66};
ram[38017] = {-9'd63,-10'd63};
ram[38018] = {-9'd60,-10'd60};
ram[38019] = {-9'd57,-10'd57};
ram[38020] = {-9'd54,-10'd54};
ram[38021] = {-9'd51,-10'd51};
ram[38022] = {-9'd48,-10'd48};
ram[38023] = {-9'd44,-10'd44};
ram[38024] = {-9'd41,-10'd41};
ram[38025] = {-9'd38,-10'd38};
ram[38026] = {-9'd35,-10'd35};
ram[38027] = {-9'd32,-10'd32};
ram[38028] = {-9'd29,-10'd29};
ram[38029] = {-9'd26,-10'd26};
ram[38030] = {-9'd22,-10'd22};
ram[38031] = {-9'd19,-10'd19};
ram[38032] = {-9'd16,-10'd16};
ram[38033] = {-9'd13,-10'd13};
ram[38034] = {-9'd10,-10'd10};
ram[38035] = {-9'd7,-10'd7};
ram[38036] = {-9'd4,-10'd4};
ram[38037] = {9'd0,10'd0};
ram[38038] = {9'd3,10'd3};
ram[38039] = {9'd6,10'd6};
ram[38040] = {9'd9,10'd9};
ram[38041] = {9'd12,10'd12};
ram[38042] = {9'd15,10'd15};
ram[38043] = {9'd18,10'd18};
ram[38044] = {9'd21,10'd21};
ram[38045] = {9'd25,10'd25};
ram[38046] = {9'd28,10'd28};
ram[38047] = {9'd31,10'd31};
ram[38048] = {9'd34,10'd34};
ram[38049] = {9'd37,10'd37};
ram[38050] = {9'd40,10'd40};
ram[38051] = {9'd43,10'd43};
ram[38052] = {9'd47,10'd47};
ram[38053] = {9'd50,10'd50};
ram[38054] = {9'd53,10'd53};
ram[38055] = {9'd56,10'd56};
ram[38056] = {9'd59,10'd59};
ram[38057] = {9'd62,10'd62};
ram[38058] = {9'd65,10'd65};
ram[38059] = {9'd69,10'd69};
ram[38060] = {9'd72,10'd72};
ram[38061] = {9'd75,10'd75};
ram[38062] = {9'd78,10'd78};
ram[38063] = {9'd81,10'd81};
ram[38064] = {9'd84,10'd84};
ram[38065] = {9'd87,10'd87};
ram[38066] = {9'd91,10'd91};
ram[38067] = {9'd94,10'd94};
ram[38068] = {9'd97,10'd97};
ram[38069] = {-9'd100,10'd100};
ram[38070] = {-9'd97,10'd103};
ram[38071] = {-9'd94,10'd106};
ram[38072] = {-9'd91,10'd109};
ram[38073] = {-9'd88,10'd113};
ram[38074] = {-9'd85,10'd116};
ram[38075] = {-9'd81,10'd119};
ram[38076] = {-9'd78,10'd122};
ram[38077] = {-9'd75,10'd125};
ram[38078] = {-9'd72,10'd128};
ram[38079] = {-9'd69,10'd131};
ram[38080] = {-9'd66,10'd135};
ram[38081] = {-9'd63,10'd138};
ram[38082] = {-9'd59,10'd141};
ram[38083] = {-9'd56,10'd144};
ram[38084] = {-9'd53,10'd147};
ram[38085] = {-9'd50,10'd150};
ram[38086] = {-9'd47,10'd153};
ram[38087] = {-9'd44,10'd157};
ram[38088] = {-9'd41,10'd160};
ram[38089] = {-9'd37,10'd163};
ram[38090] = {-9'd34,10'd166};
ram[38091] = {-9'd31,10'd169};
ram[38092] = {-9'd28,10'd172};
ram[38093] = {-9'd25,10'd175};
ram[38094] = {-9'd22,10'd179};
ram[38095] = {-9'd19,10'd182};
ram[38096] = {-9'd15,10'd185};
ram[38097] = {-9'd12,10'd188};
ram[38098] = {-9'd9,10'd191};
ram[38099] = {-9'd6,10'd194};
ram[38100] = {-9'd3,10'd197};
ram[38101] = {9'd0,10'd201};
ram[38102] = {9'd3,10'd204};
ram[38103] = {9'd7,10'd207};
ram[38104] = {9'd10,10'd210};
ram[38105] = {9'd13,10'd213};
ram[38106] = {9'd16,10'd216};
ram[38107] = {9'd19,10'd219};
ram[38108] = {9'd22,10'd223};
ram[38109] = {9'd25,10'd226};
ram[38110] = {9'd29,10'd229};
ram[38111] = {9'd32,10'd232};
ram[38112] = {9'd35,10'd235};
ram[38113] = {9'd38,10'd238};
ram[38114] = {9'd41,10'd241};
ram[38115] = {9'd44,10'd245};
ram[38116] = {9'd47,10'd248};
ram[38117] = {9'd51,10'd251};
ram[38118] = {9'd54,10'd254};
ram[38119] = {9'd57,10'd257};
ram[38120] = {9'd60,10'd260};
ram[38121] = {9'd63,10'd263};
ram[38122] = {9'd66,10'd267};
ram[38123] = {9'd69,10'd270};
ram[38124] = {9'd73,10'd273};
ram[38125] = {9'd76,10'd276};
ram[38126] = {9'd79,10'd279};
ram[38127] = {9'd82,10'd282};
ram[38128] = {9'd85,10'd285};
ram[38129] = {9'd88,10'd289};
ram[38130] = {9'd91,10'd292};
ram[38131] = {9'd95,10'd295};
ram[38132] = {9'd98,10'd298};
ram[38133] = {-9'd99,10'd301};
ram[38134] = {-9'd96,10'd304};
ram[38135] = {-9'd93,10'd307};
ram[38136] = {-9'd90,10'd311};
ram[38137] = {-9'd87,10'd314};
ram[38138] = {-9'd84,10'd317};
ram[38139] = {-9'd81,10'd320};
ram[38140] = {-9'd77,10'd323};
ram[38141] = {-9'd74,10'd326};
ram[38142] = {-9'd71,10'd329};
ram[38143] = {-9'd68,10'd333};
ram[38144] = {-9'd68,10'd333};
ram[38145] = {-9'd65,10'd336};
ram[38146] = {-9'd62,10'd339};
ram[38147] = {-9'd59,10'd342};
ram[38148] = {-9'd55,10'd345};
ram[38149] = {-9'd52,10'd348};
ram[38150] = {-9'd49,10'd351};
ram[38151] = {-9'd46,10'd354};
ram[38152] = {-9'd43,10'd358};
ram[38153] = {-9'd40,10'd361};
ram[38154] = {-9'd37,10'd364};
ram[38155] = {-9'd33,10'd367};
ram[38156] = {-9'd30,10'd370};
ram[38157] = {-9'd27,10'd373};
ram[38158] = {-9'd24,10'd376};
ram[38159] = {-9'd21,10'd380};
ram[38160] = {-9'd18,10'd383};
ram[38161] = {-9'd15,10'd386};
ram[38162] = {-9'd11,10'd389};
ram[38163] = {-9'd8,10'd392};
ram[38164] = {-9'd5,10'd395};
ram[38165] = {-9'd2,10'd398};
ram[38166] = {9'd1,-10'd399};
ram[38167] = {9'd4,-10'd396};
ram[38168] = {9'd7,-10'd393};
ram[38169] = {9'd10,-10'd390};
ram[38170] = {9'd14,-10'd387};
ram[38171] = {9'd17,-10'd384};
ram[38172] = {9'd20,-10'd381};
ram[38173] = {9'd23,-10'd377};
ram[38174] = {9'd26,-10'd374};
ram[38175] = {9'd29,-10'd371};
ram[38176] = {9'd32,-10'd368};
ram[38177] = {9'd36,-10'd365};
ram[38178] = {9'd39,-10'd362};
ram[38179] = {9'd42,-10'd359};
ram[38180] = {9'd45,-10'd355};
ram[38181] = {9'd48,-10'd352};
ram[38182] = {9'd51,-10'd349};
ram[38183] = {9'd54,-10'd346};
ram[38184] = {9'd58,-10'd343};
ram[38185] = {9'd61,-10'd340};
ram[38186] = {9'd64,-10'd337};
ram[38187] = {9'd67,-10'd334};
ram[38188] = {9'd70,-10'd330};
ram[38189] = {9'd73,-10'd327};
ram[38190] = {9'd76,-10'd324};
ram[38191] = {9'd80,-10'd321};
ram[38192] = {9'd83,-10'd318};
ram[38193] = {9'd86,-10'd315};
ram[38194] = {9'd89,-10'd312};
ram[38195] = {9'd92,-10'd308};
ram[38196] = {9'd95,-10'd305};
ram[38197] = {9'd98,-10'd302};
ram[38198] = {-9'd99,-10'd299};
ram[38199] = {-9'd96,-10'd296};
ram[38200] = {-9'd92,-10'd293};
ram[38201] = {-9'd89,-10'd290};
ram[38202] = {-9'd86,-10'd286};
ram[38203] = {-9'd83,-10'd283};
ram[38204] = {-9'd80,-10'd280};
ram[38205] = {-9'd77,-10'd277};
ram[38206] = {-9'd74,-10'd274};
ram[38207] = {-9'd70,-10'd271};
ram[38208] = {-9'd67,-10'd268};
ram[38209] = {-9'd64,-10'd264};
ram[38210] = {-9'd61,-10'd261};
ram[38211] = {-9'd58,-10'd258};
ram[38212] = {-9'd55,-10'd255};
ram[38213] = {-9'd52,-10'd252};
ram[38214] = {-9'd48,-10'd249};
ram[38215] = {-9'd45,-10'd246};
ram[38216] = {-9'd42,-10'd242};
ram[38217] = {-9'd39,-10'd239};
ram[38218] = {-9'd36,-10'd236};
ram[38219] = {-9'd33,-10'd233};
ram[38220] = {-9'd30,-10'd230};
ram[38221] = {-9'd26,-10'd227};
ram[38222] = {-9'd23,-10'd224};
ram[38223] = {-9'd20,-10'd220};
ram[38224] = {-9'd17,-10'd217};
ram[38225] = {-9'd14,-10'd214};
ram[38226] = {-9'd11,-10'd211};
ram[38227] = {-9'd8,-10'd208};
ram[38228] = {-9'd4,-10'd205};
ram[38229] = {-9'd1,-10'd202};
ram[38230] = {9'd2,-10'd198};
ram[38231] = {9'd5,-10'd195};
ram[38232] = {9'd8,-10'd192};
ram[38233] = {9'd11,-10'd189};
ram[38234] = {9'd14,-10'd186};
ram[38235] = {9'd18,-10'd183};
ram[38236] = {9'd21,-10'd180};
ram[38237] = {9'd24,-10'd176};
ram[38238] = {9'd27,-10'd173};
ram[38239] = {9'd30,-10'd170};
ram[38240] = {9'd33,-10'd167};
ram[38241] = {9'd36,-10'd164};
ram[38242] = {9'd40,-10'd161};
ram[38243] = {9'd43,-10'd158};
ram[38244] = {9'd46,-10'd154};
ram[38245] = {9'd49,-10'd151};
ram[38246] = {9'd52,-10'd148};
ram[38247] = {9'd55,-10'd145};
ram[38248] = {9'd58,-10'd142};
ram[38249] = {9'd62,-10'd139};
ram[38250] = {9'd65,-10'd136};
ram[38251] = {9'd68,-10'd132};
ram[38252] = {9'd71,-10'd129};
ram[38253] = {9'd74,-10'd126};
ram[38254] = {9'd77,-10'd123};
ram[38255] = {9'd80,-10'd120};
ram[38256] = {9'd84,-10'd117};
ram[38257] = {9'd87,-10'd114};
ram[38258] = {9'd90,-10'd110};
ram[38259] = {9'd93,-10'd107};
ram[38260] = {9'd96,-10'd104};
ram[38261] = {9'd99,-10'd101};
ram[38262] = {-9'd98,-10'd98};
ram[38263] = {-9'd95,-10'd95};
ram[38264] = {-9'd92,-10'd92};
ram[38265] = {-9'd88,-10'd88};
ram[38266] = {-9'd85,-10'd85};
ram[38267] = {-9'd82,-10'd82};
ram[38268] = {-9'd79,-10'd79};
ram[38269] = {-9'd76,-10'd76};
ram[38270] = {-9'd73,-10'd73};
ram[38271] = {-9'd70,-10'd70};
ram[38272] = {-9'd70,-10'd70};
ram[38273] = {-9'd66,-10'd66};
ram[38274] = {-9'd63,-10'd63};
ram[38275] = {-9'd60,-10'd60};
ram[38276] = {-9'd57,-10'd57};
ram[38277] = {-9'd54,-10'd54};
ram[38278] = {-9'd51,-10'd51};
ram[38279] = {-9'd48,-10'd48};
ram[38280] = {-9'd44,-10'd44};
ram[38281] = {-9'd41,-10'd41};
ram[38282] = {-9'd38,-10'd38};
ram[38283] = {-9'd35,-10'd35};
ram[38284] = {-9'd32,-10'd32};
ram[38285] = {-9'd29,-10'd29};
ram[38286] = {-9'd26,-10'd26};
ram[38287] = {-9'd22,-10'd22};
ram[38288] = {-9'd19,-10'd19};
ram[38289] = {-9'd16,-10'd16};
ram[38290] = {-9'd13,-10'd13};
ram[38291] = {-9'd10,-10'd10};
ram[38292] = {-9'd7,-10'd7};
ram[38293] = {-9'd4,-10'd4};
ram[38294] = {9'd0,10'd0};
ram[38295] = {9'd3,10'd3};
ram[38296] = {9'd6,10'd6};
ram[38297] = {9'd9,10'd9};
ram[38298] = {9'd12,10'd12};
ram[38299] = {9'd15,10'd15};
ram[38300] = {9'd18,10'd18};
ram[38301] = {9'd21,10'd21};
ram[38302] = {9'd25,10'd25};
ram[38303] = {9'd28,10'd28};
ram[38304] = {9'd31,10'd31};
ram[38305] = {9'd34,10'd34};
ram[38306] = {9'd37,10'd37};
ram[38307] = {9'd40,10'd40};
ram[38308] = {9'd43,10'd43};
ram[38309] = {9'd47,10'd47};
ram[38310] = {9'd50,10'd50};
ram[38311] = {9'd53,10'd53};
ram[38312] = {9'd56,10'd56};
ram[38313] = {9'd59,10'd59};
ram[38314] = {9'd62,10'd62};
ram[38315] = {9'd65,10'd65};
ram[38316] = {9'd69,10'd69};
ram[38317] = {9'd72,10'd72};
ram[38318] = {9'd75,10'd75};
ram[38319] = {9'd78,10'd78};
ram[38320] = {9'd81,10'd81};
ram[38321] = {9'd84,10'd84};
ram[38322] = {9'd87,10'd87};
ram[38323] = {9'd91,10'd91};
ram[38324] = {9'd94,10'd94};
ram[38325] = {9'd97,10'd97};
ram[38326] = {-9'd100,10'd100};
ram[38327] = {-9'd97,10'd103};
ram[38328] = {-9'd94,10'd106};
ram[38329] = {-9'd91,10'd109};
ram[38330] = {-9'd88,10'd113};
ram[38331] = {-9'd85,10'd116};
ram[38332] = {-9'd81,10'd119};
ram[38333] = {-9'd78,10'd122};
ram[38334] = {-9'd75,10'd125};
ram[38335] = {-9'd72,10'd128};
ram[38336] = {-9'd69,10'd131};
ram[38337] = {-9'd66,10'd135};
ram[38338] = {-9'd63,10'd138};
ram[38339] = {-9'd59,10'd141};
ram[38340] = {-9'd56,10'd144};
ram[38341] = {-9'd53,10'd147};
ram[38342] = {-9'd50,10'd150};
ram[38343] = {-9'd47,10'd153};
ram[38344] = {-9'd44,10'd157};
ram[38345] = {-9'd41,10'd160};
ram[38346] = {-9'd37,10'd163};
ram[38347] = {-9'd34,10'd166};
ram[38348] = {-9'd31,10'd169};
ram[38349] = {-9'd28,10'd172};
ram[38350] = {-9'd25,10'd175};
ram[38351] = {-9'd22,10'd179};
ram[38352] = {-9'd19,10'd182};
ram[38353] = {-9'd15,10'd185};
ram[38354] = {-9'd12,10'd188};
ram[38355] = {-9'd9,10'd191};
ram[38356] = {-9'd6,10'd194};
ram[38357] = {-9'd3,10'd197};
ram[38358] = {9'd0,10'd201};
ram[38359] = {9'd3,10'd204};
ram[38360] = {9'd7,10'd207};
ram[38361] = {9'd10,10'd210};
ram[38362] = {9'd13,10'd213};
ram[38363] = {9'd16,10'd216};
ram[38364] = {9'd19,10'd219};
ram[38365] = {9'd22,10'd223};
ram[38366] = {9'd25,10'd226};
ram[38367] = {9'd29,10'd229};
ram[38368] = {9'd32,10'd232};
ram[38369] = {9'd35,10'd235};
ram[38370] = {9'd38,10'd238};
ram[38371] = {9'd41,10'd241};
ram[38372] = {9'd44,10'd245};
ram[38373] = {9'd47,10'd248};
ram[38374] = {9'd51,10'd251};
ram[38375] = {9'd54,10'd254};
ram[38376] = {9'd57,10'd257};
ram[38377] = {9'd60,10'd260};
ram[38378] = {9'd63,10'd263};
ram[38379] = {9'd66,10'd267};
ram[38380] = {9'd69,10'd270};
ram[38381] = {9'd73,10'd273};
ram[38382] = {9'd76,10'd276};
ram[38383] = {9'd79,10'd279};
ram[38384] = {9'd82,10'd282};
ram[38385] = {9'd85,10'd285};
ram[38386] = {9'd88,10'd289};
ram[38387] = {9'd91,10'd292};
ram[38388] = {9'd95,10'd295};
ram[38389] = {9'd98,10'd298};
ram[38390] = {-9'd99,10'd301};
ram[38391] = {-9'd96,10'd304};
ram[38392] = {-9'd93,10'd307};
ram[38393] = {-9'd90,10'd311};
ram[38394] = {-9'd87,10'd314};
ram[38395] = {-9'd84,10'd317};
ram[38396] = {-9'd81,10'd320};
ram[38397] = {-9'd77,10'd323};
ram[38398] = {-9'd74,10'd326};
ram[38399] = {-9'd71,10'd329};
ram[38400] = {-9'd71,10'd329};
ram[38401] = {-9'd68,10'd333};
ram[38402] = {-9'd65,10'd336};
ram[38403] = {-9'd62,10'd339};
ram[38404] = {-9'd59,10'd342};
ram[38405] = {-9'd55,10'd345};
ram[38406] = {-9'd52,10'd348};
ram[38407] = {-9'd49,10'd351};
ram[38408] = {-9'd46,10'd354};
ram[38409] = {-9'd43,10'd358};
ram[38410] = {-9'd40,10'd361};
ram[38411] = {-9'd37,10'd364};
ram[38412] = {-9'd33,10'd367};
ram[38413] = {-9'd30,10'd370};
ram[38414] = {-9'd27,10'd373};
ram[38415] = {-9'd24,10'd376};
ram[38416] = {-9'd21,10'd380};
ram[38417] = {-9'd18,10'd383};
ram[38418] = {-9'd15,10'd386};
ram[38419] = {-9'd11,10'd389};
ram[38420] = {-9'd8,10'd392};
ram[38421] = {-9'd5,10'd395};
ram[38422] = {-9'd2,10'd398};
ram[38423] = {9'd1,-10'd399};
ram[38424] = {9'd4,-10'd396};
ram[38425] = {9'd7,-10'd393};
ram[38426] = {9'd10,-10'd390};
ram[38427] = {9'd14,-10'd387};
ram[38428] = {9'd17,-10'd384};
ram[38429] = {9'd20,-10'd381};
ram[38430] = {9'd23,-10'd377};
ram[38431] = {9'd26,-10'd374};
ram[38432] = {9'd29,-10'd371};
ram[38433] = {9'd32,-10'd368};
ram[38434] = {9'd36,-10'd365};
ram[38435] = {9'd39,-10'd362};
ram[38436] = {9'd42,-10'd359};
ram[38437] = {9'd45,-10'd355};
ram[38438] = {9'd48,-10'd352};
ram[38439] = {9'd51,-10'd349};
ram[38440] = {9'd54,-10'd346};
ram[38441] = {9'd58,-10'd343};
ram[38442] = {9'd61,-10'd340};
ram[38443] = {9'd64,-10'd337};
ram[38444] = {9'd67,-10'd334};
ram[38445] = {9'd70,-10'd330};
ram[38446] = {9'd73,-10'd327};
ram[38447] = {9'd76,-10'd324};
ram[38448] = {9'd80,-10'd321};
ram[38449] = {9'd83,-10'd318};
ram[38450] = {9'd86,-10'd315};
ram[38451] = {9'd89,-10'd312};
ram[38452] = {9'd92,-10'd308};
ram[38453] = {9'd95,-10'd305};
ram[38454] = {9'd98,-10'd302};
ram[38455] = {-9'd99,-10'd299};
ram[38456] = {-9'd96,-10'd296};
ram[38457] = {-9'd92,-10'd293};
ram[38458] = {-9'd89,-10'd290};
ram[38459] = {-9'd86,-10'd286};
ram[38460] = {-9'd83,-10'd283};
ram[38461] = {-9'd80,-10'd280};
ram[38462] = {-9'd77,-10'd277};
ram[38463] = {-9'd74,-10'd274};
ram[38464] = {-9'd70,-10'd271};
ram[38465] = {-9'd67,-10'd268};
ram[38466] = {-9'd64,-10'd264};
ram[38467] = {-9'd61,-10'd261};
ram[38468] = {-9'd58,-10'd258};
ram[38469] = {-9'd55,-10'd255};
ram[38470] = {-9'd52,-10'd252};
ram[38471] = {-9'd48,-10'd249};
ram[38472] = {-9'd45,-10'd246};
ram[38473] = {-9'd42,-10'd242};
ram[38474] = {-9'd39,-10'd239};
ram[38475] = {-9'd36,-10'd236};
ram[38476] = {-9'd33,-10'd233};
ram[38477] = {-9'd30,-10'd230};
ram[38478] = {-9'd26,-10'd227};
ram[38479] = {-9'd23,-10'd224};
ram[38480] = {-9'd20,-10'd220};
ram[38481] = {-9'd17,-10'd217};
ram[38482] = {-9'd14,-10'd214};
ram[38483] = {-9'd11,-10'd211};
ram[38484] = {-9'd8,-10'd208};
ram[38485] = {-9'd4,-10'd205};
ram[38486] = {-9'd1,-10'd202};
ram[38487] = {9'd2,-10'd198};
ram[38488] = {9'd5,-10'd195};
ram[38489] = {9'd8,-10'd192};
ram[38490] = {9'd11,-10'd189};
ram[38491] = {9'd14,-10'd186};
ram[38492] = {9'd18,-10'd183};
ram[38493] = {9'd21,-10'd180};
ram[38494] = {9'd24,-10'd176};
ram[38495] = {9'd27,-10'd173};
ram[38496] = {9'd30,-10'd170};
ram[38497] = {9'd33,-10'd167};
ram[38498] = {9'd36,-10'd164};
ram[38499] = {9'd40,-10'd161};
ram[38500] = {9'd43,-10'd158};
ram[38501] = {9'd46,-10'd154};
ram[38502] = {9'd49,-10'd151};
ram[38503] = {9'd52,-10'd148};
ram[38504] = {9'd55,-10'd145};
ram[38505] = {9'd58,-10'd142};
ram[38506] = {9'd62,-10'd139};
ram[38507] = {9'd65,-10'd136};
ram[38508] = {9'd68,-10'd132};
ram[38509] = {9'd71,-10'd129};
ram[38510] = {9'd74,-10'd126};
ram[38511] = {9'd77,-10'd123};
ram[38512] = {9'd80,-10'd120};
ram[38513] = {9'd84,-10'd117};
ram[38514] = {9'd87,-10'd114};
ram[38515] = {9'd90,-10'd110};
ram[38516] = {9'd93,-10'd107};
ram[38517] = {9'd96,-10'd104};
ram[38518] = {9'd99,-10'd101};
ram[38519] = {-9'd98,-10'd98};
ram[38520] = {-9'd95,-10'd95};
ram[38521] = {-9'd92,-10'd92};
ram[38522] = {-9'd88,-10'd88};
ram[38523] = {-9'd85,-10'd85};
ram[38524] = {-9'd82,-10'd82};
ram[38525] = {-9'd79,-10'd79};
ram[38526] = {-9'd76,-10'd76};
ram[38527] = {-9'd73,-10'd73};
ram[38528] = {-9'd73,-10'd73};
ram[38529] = {-9'd70,-10'd70};
ram[38530] = {-9'd66,-10'd66};
ram[38531] = {-9'd63,-10'd63};
ram[38532] = {-9'd60,-10'd60};
ram[38533] = {-9'd57,-10'd57};
ram[38534] = {-9'd54,-10'd54};
ram[38535] = {-9'd51,-10'd51};
ram[38536] = {-9'd48,-10'd48};
ram[38537] = {-9'd44,-10'd44};
ram[38538] = {-9'd41,-10'd41};
ram[38539] = {-9'd38,-10'd38};
ram[38540] = {-9'd35,-10'd35};
ram[38541] = {-9'd32,-10'd32};
ram[38542] = {-9'd29,-10'd29};
ram[38543] = {-9'd26,-10'd26};
ram[38544] = {-9'd22,-10'd22};
ram[38545] = {-9'd19,-10'd19};
ram[38546] = {-9'd16,-10'd16};
ram[38547] = {-9'd13,-10'd13};
ram[38548] = {-9'd10,-10'd10};
ram[38549] = {-9'd7,-10'd7};
ram[38550] = {-9'd4,-10'd4};
ram[38551] = {9'd0,10'd0};
ram[38552] = {9'd3,10'd3};
ram[38553] = {9'd6,10'd6};
ram[38554] = {9'd9,10'd9};
ram[38555] = {9'd12,10'd12};
ram[38556] = {9'd15,10'd15};
ram[38557] = {9'd18,10'd18};
ram[38558] = {9'd21,10'd21};
ram[38559] = {9'd25,10'd25};
ram[38560] = {9'd28,10'd28};
ram[38561] = {9'd31,10'd31};
ram[38562] = {9'd34,10'd34};
ram[38563] = {9'd37,10'd37};
ram[38564] = {9'd40,10'd40};
ram[38565] = {9'd43,10'd43};
ram[38566] = {9'd47,10'd47};
ram[38567] = {9'd50,10'd50};
ram[38568] = {9'd53,10'd53};
ram[38569] = {9'd56,10'd56};
ram[38570] = {9'd59,10'd59};
ram[38571] = {9'd62,10'd62};
ram[38572] = {9'd65,10'd65};
ram[38573] = {9'd69,10'd69};
ram[38574] = {9'd72,10'd72};
ram[38575] = {9'd75,10'd75};
ram[38576] = {9'd78,10'd78};
ram[38577] = {9'd81,10'd81};
ram[38578] = {9'd84,10'd84};
ram[38579] = {9'd87,10'd87};
ram[38580] = {9'd91,10'd91};
ram[38581] = {9'd94,10'd94};
ram[38582] = {9'd97,10'd97};
ram[38583] = {-9'd100,10'd100};
ram[38584] = {-9'd97,10'd103};
ram[38585] = {-9'd94,10'd106};
ram[38586] = {-9'd91,10'd109};
ram[38587] = {-9'd88,10'd113};
ram[38588] = {-9'd85,10'd116};
ram[38589] = {-9'd81,10'd119};
ram[38590] = {-9'd78,10'd122};
ram[38591] = {-9'd75,10'd125};
ram[38592] = {-9'd72,10'd128};
ram[38593] = {-9'd69,10'd131};
ram[38594] = {-9'd66,10'd135};
ram[38595] = {-9'd63,10'd138};
ram[38596] = {-9'd59,10'd141};
ram[38597] = {-9'd56,10'd144};
ram[38598] = {-9'd53,10'd147};
ram[38599] = {-9'd50,10'd150};
ram[38600] = {-9'd47,10'd153};
ram[38601] = {-9'd44,10'd157};
ram[38602] = {-9'd41,10'd160};
ram[38603] = {-9'd37,10'd163};
ram[38604] = {-9'd34,10'd166};
ram[38605] = {-9'd31,10'd169};
ram[38606] = {-9'd28,10'd172};
ram[38607] = {-9'd25,10'd175};
ram[38608] = {-9'd22,10'd179};
ram[38609] = {-9'd19,10'd182};
ram[38610] = {-9'd15,10'd185};
ram[38611] = {-9'd12,10'd188};
ram[38612] = {-9'd9,10'd191};
ram[38613] = {-9'd6,10'd194};
ram[38614] = {-9'd3,10'd197};
ram[38615] = {9'd0,10'd201};
ram[38616] = {9'd3,10'd204};
ram[38617] = {9'd7,10'd207};
ram[38618] = {9'd10,10'd210};
ram[38619] = {9'd13,10'd213};
ram[38620] = {9'd16,10'd216};
ram[38621] = {9'd19,10'd219};
ram[38622] = {9'd22,10'd223};
ram[38623] = {9'd25,10'd226};
ram[38624] = {9'd29,10'd229};
ram[38625] = {9'd32,10'd232};
ram[38626] = {9'd35,10'd235};
ram[38627] = {9'd38,10'd238};
ram[38628] = {9'd41,10'd241};
ram[38629] = {9'd44,10'd245};
ram[38630] = {9'd47,10'd248};
ram[38631] = {9'd51,10'd251};
ram[38632] = {9'd54,10'd254};
ram[38633] = {9'd57,10'd257};
ram[38634] = {9'd60,10'd260};
ram[38635] = {9'd63,10'd263};
ram[38636] = {9'd66,10'd267};
ram[38637] = {9'd69,10'd270};
ram[38638] = {9'd73,10'd273};
ram[38639] = {9'd76,10'd276};
ram[38640] = {9'd79,10'd279};
ram[38641] = {9'd82,10'd282};
ram[38642] = {9'd85,10'd285};
ram[38643] = {9'd88,10'd289};
ram[38644] = {9'd91,10'd292};
ram[38645] = {9'd95,10'd295};
ram[38646] = {9'd98,10'd298};
ram[38647] = {-9'd99,10'd301};
ram[38648] = {-9'd96,10'd304};
ram[38649] = {-9'd93,10'd307};
ram[38650] = {-9'd90,10'd311};
ram[38651] = {-9'd87,10'd314};
ram[38652] = {-9'd84,10'd317};
ram[38653] = {-9'd81,10'd320};
ram[38654] = {-9'd77,10'd323};
ram[38655] = {-9'd74,10'd326};
ram[38656] = {-9'd74,10'd326};
ram[38657] = {-9'd71,10'd329};
ram[38658] = {-9'd68,10'd333};
ram[38659] = {-9'd65,10'd336};
ram[38660] = {-9'd62,10'd339};
ram[38661] = {-9'd59,10'd342};
ram[38662] = {-9'd55,10'd345};
ram[38663] = {-9'd52,10'd348};
ram[38664] = {-9'd49,10'd351};
ram[38665] = {-9'd46,10'd354};
ram[38666] = {-9'd43,10'd358};
ram[38667] = {-9'd40,10'd361};
ram[38668] = {-9'd37,10'd364};
ram[38669] = {-9'd33,10'd367};
ram[38670] = {-9'd30,10'd370};
ram[38671] = {-9'd27,10'd373};
ram[38672] = {-9'd24,10'd376};
ram[38673] = {-9'd21,10'd380};
ram[38674] = {-9'd18,10'd383};
ram[38675] = {-9'd15,10'd386};
ram[38676] = {-9'd11,10'd389};
ram[38677] = {-9'd8,10'd392};
ram[38678] = {-9'd5,10'd395};
ram[38679] = {-9'd2,10'd398};
ram[38680] = {9'd1,-10'd399};
ram[38681] = {9'd4,-10'd396};
ram[38682] = {9'd7,-10'd393};
ram[38683] = {9'd10,-10'd390};
ram[38684] = {9'd14,-10'd387};
ram[38685] = {9'd17,-10'd384};
ram[38686] = {9'd20,-10'd381};
ram[38687] = {9'd23,-10'd377};
ram[38688] = {9'd26,-10'd374};
ram[38689] = {9'd29,-10'd371};
ram[38690] = {9'd32,-10'd368};
ram[38691] = {9'd36,-10'd365};
ram[38692] = {9'd39,-10'd362};
ram[38693] = {9'd42,-10'd359};
ram[38694] = {9'd45,-10'd355};
ram[38695] = {9'd48,-10'd352};
ram[38696] = {9'd51,-10'd349};
ram[38697] = {9'd54,-10'd346};
ram[38698] = {9'd58,-10'd343};
ram[38699] = {9'd61,-10'd340};
ram[38700] = {9'd64,-10'd337};
ram[38701] = {9'd67,-10'd334};
ram[38702] = {9'd70,-10'd330};
ram[38703] = {9'd73,-10'd327};
ram[38704] = {9'd76,-10'd324};
ram[38705] = {9'd80,-10'd321};
ram[38706] = {9'd83,-10'd318};
ram[38707] = {9'd86,-10'd315};
ram[38708] = {9'd89,-10'd312};
ram[38709] = {9'd92,-10'd308};
ram[38710] = {9'd95,-10'd305};
ram[38711] = {9'd98,-10'd302};
ram[38712] = {-9'd99,-10'd299};
ram[38713] = {-9'd96,-10'd296};
ram[38714] = {-9'd92,-10'd293};
ram[38715] = {-9'd89,-10'd290};
ram[38716] = {-9'd86,-10'd286};
ram[38717] = {-9'd83,-10'd283};
ram[38718] = {-9'd80,-10'd280};
ram[38719] = {-9'd77,-10'd277};
ram[38720] = {-9'd74,-10'd274};
ram[38721] = {-9'd70,-10'd271};
ram[38722] = {-9'd67,-10'd268};
ram[38723] = {-9'd64,-10'd264};
ram[38724] = {-9'd61,-10'd261};
ram[38725] = {-9'd58,-10'd258};
ram[38726] = {-9'd55,-10'd255};
ram[38727] = {-9'd52,-10'd252};
ram[38728] = {-9'd48,-10'd249};
ram[38729] = {-9'd45,-10'd246};
ram[38730] = {-9'd42,-10'd242};
ram[38731] = {-9'd39,-10'd239};
ram[38732] = {-9'd36,-10'd236};
ram[38733] = {-9'd33,-10'd233};
ram[38734] = {-9'd30,-10'd230};
ram[38735] = {-9'd26,-10'd227};
ram[38736] = {-9'd23,-10'd224};
ram[38737] = {-9'd20,-10'd220};
ram[38738] = {-9'd17,-10'd217};
ram[38739] = {-9'd14,-10'd214};
ram[38740] = {-9'd11,-10'd211};
ram[38741] = {-9'd8,-10'd208};
ram[38742] = {-9'd4,-10'd205};
ram[38743] = {-9'd1,-10'd202};
ram[38744] = {9'd2,-10'd198};
ram[38745] = {9'd5,-10'd195};
ram[38746] = {9'd8,-10'd192};
ram[38747] = {9'd11,-10'd189};
ram[38748] = {9'd14,-10'd186};
ram[38749] = {9'd18,-10'd183};
ram[38750] = {9'd21,-10'd180};
ram[38751] = {9'd24,-10'd176};
ram[38752] = {9'd27,-10'd173};
ram[38753] = {9'd30,-10'd170};
ram[38754] = {9'd33,-10'd167};
ram[38755] = {9'd36,-10'd164};
ram[38756] = {9'd40,-10'd161};
ram[38757] = {9'd43,-10'd158};
ram[38758] = {9'd46,-10'd154};
ram[38759] = {9'd49,-10'd151};
ram[38760] = {9'd52,-10'd148};
ram[38761] = {9'd55,-10'd145};
ram[38762] = {9'd58,-10'd142};
ram[38763] = {9'd62,-10'd139};
ram[38764] = {9'd65,-10'd136};
ram[38765] = {9'd68,-10'd132};
ram[38766] = {9'd71,-10'd129};
ram[38767] = {9'd74,-10'd126};
ram[38768] = {9'd77,-10'd123};
ram[38769] = {9'd80,-10'd120};
ram[38770] = {9'd84,-10'd117};
ram[38771] = {9'd87,-10'd114};
ram[38772] = {9'd90,-10'd110};
ram[38773] = {9'd93,-10'd107};
ram[38774] = {9'd96,-10'd104};
ram[38775] = {9'd99,-10'd101};
ram[38776] = {-9'd98,-10'd98};
ram[38777] = {-9'd95,-10'd95};
ram[38778] = {-9'd92,-10'd92};
ram[38779] = {-9'd88,-10'd88};
ram[38780] = {-9'd85,-10'd85};
ram[38781] = {-9'd82,-10'd82};
ram[38782] = {-9'd79,-10'd79};
ram[38783] = {-9'd76,-10'd76};
ram[38784] = {-9'd76,-10'd76};
ram[38785] = {-9'd73,-10'd73};
ram[38786] = {-9'd70,-10'd70};
ram[38787] = {-9'd66,-10'd66};
ram[38788] = {-9'd63,-10'd63};
ram[38789] = {-9'd60,-10'd60};
ram[38790] = {-9'd57,-10'd57};
ram[38791] = {-9'd54,-10'd54};
ram[38792] = {-9'd51,-10'd51};
ram[38793] = {-9'd48,-10'd48};
ram[38794] = {-9'd44,-10'd44};
ram[38795] = {-9'd41,-10'd41};
ram[38796] = {-9'd38,-10'd38};
ram[38797] = {-9'd35,-10'd35};
ram[38798] = {-9'd32,-10'd32};
ram[38799] = {-9'd29,-10'd29};
ram[38800] = {-9'd26,-10'd26};
ram[38801] = {-9'd22,-10'd22};
ram[38802] = {-9'd19,-10'd19};
ram[38803] = {-9'd16,-10'd16};
ram[38804] = {-9'd13,-10'd13};
ram[38805] = {-9'd10,-10'd10};
ram[38806] = {-9'd7,-10'd7};
ram[38807] = {-9'd4,-10'd4};
ram[38808] = {9'd0,10'd0};
ram[38809] = {9'd3,10'd3};
ram[38810] = {9'd6,10'd6};
ram[38811] = {9'd9,10'd9};
ram[38812] = {9'd12,10'd12};
ram[38813] = {9'd15,10'd15};
ram[38814] = {9'd18,10'd18};
ram[38815] = {9'd21,10'd21};
ram[38816] = {9'd25,10'd25};
ram[38817] = {9'd28,10'd28};
ram[38818] = {9'd31,10'd31};
ram[38819] = {9'd34,10'd34};
ram[38820] = {9'd37,10'd37};
ram[38821] = {9'd40,10'd40};
ram[38822] = {9'd43,10'd43};
ram[38823] = {9'd47,10'd47};
ram[38824] = {9'd50,10'd50};
ram[38825] = {9'd53,10'd53};
ram[38826] = {9'd56,10'd56};
ram[38827] = {9'd59,10'd59};
ram[38828] = {9'd62,10'd62};
ram[38829] = {9'd65,10'd65};
ram[38830] = {9'd69,10'd69};
ram[38831] = {9'd72,10'd72};
ram[38832] = {9'd75,10'd75};
ram[38833] = {9'd78,10'd78};
ram[38834] = {9'd81,10'd81};
ram[38835] = {9'd84,10'd84};
ram[38836] = {9'd87,10'd87};
ram[38837] = {9'd91,10'd91};
ram[38838] = {9'd94,10'd94};
ram[38839] = {9'd97,10'd97};
ram[38840] = {-9'd100,10'd100};
ram[38841] = {-9'd97,10'd103};
ram[38842] = {-9'd94,10'd106};
ram[38843] = {-9'd91,10'd109};
ram[38844] = {-9'd88,10'd113};
ram[38845] = {-9'd85,10'd116};
ram[38846] = {-9'd81,10'd119};
ram[38847] = {-9'd78,10'd122};
ram[38848] = {-9'd75,10'd125};
ram[38849] = {-9'd72,10'd128};
ram[38850] = {-9'd69,10'd131};
ram[38851] = {-9'd66,10'd135};
ram[38852] = {-9'd63,10'd138};
ram[38853] = {-9'd59,10'd141};
ram[38854] = {-9'd56,10'd144};
ram[38855] = {-9'd53,10'd147};
ram[38856] = {-9'd50,10'd150};
ram[38857] = {-9'd47,10'd153};
ram[38858] = {-9'd44,10'd157};
ram[38859] = {-9'd41,10'd160};
ram[38860] = {-9'd37,10'd163};
ram[38861] = {-9'd34,10'd166};
ram[38862] = {-9'd31,10'd169};
ram[38863] = {-9'd28,10'd172};
ram[38864] = {-9'd25,10'd175};
ram[38865] = {-9'd22,10'd179};
ram[38866] = {-9'd19,10'd182};
ram[38867] = {-9'd15,10'd185};
ram[38868] = {-9'd12,10'd188};
ram[38869] = {-9'd9,10'd191};
ram[38870] = {-9'd6,10'd194};
ram[38871] = {-9'd3,10'd197};
ram[38872] = {9'd0,10'd201};
ram[38873] = {9'd3,10'd204};
ram[38874] = {9'd7,10'd207};
ram[38875] = {9'd10,10'd210};
ram[38876] = {9'd13,10'd213};
ram[38877] = {9'd16,10'd216};
ram[38878] = {9'd19,10'd219};
ram[38879] = {9'd22,10'd223};
ram[38880] = {9'd25,10'd226};
ram[38881] = {9'd29,10'd229};
ram[38882] = {9'd32,10'd232};
ram[38883] = {9'd35,10'd235};
ram[38884] = {9'd38,10'd238};
ram[38885] = {9'd41,10'd241};
ram[38886] = {9'd44,10'd245};
ram[38887] = {9'd47,10'd248};
ram[38888] = {9'd51,10'd251};
ram[38889] = {9'd54,10'd254};
ram[38890] = {9'd57,10'd257};
ram[38891] = {9'd60,10'd260};
ram[38892] = {9'd63,10'd263};
ram[38893] = {9'd66,10'd267};
ram[38894] = {9'd69,10'd270};
ram[38895] = {9'd73,10'd273};
ram[38896] = {9'd76,10'd276};
ram[38897] = {9'd79,10'd279};
ram[38898] = {9'd82,10'd282};
ram[38899] = {9'd85,10'd285};
ram[38900] = {9'd88,10'd289};
ram[38901] = {9'd91,10'd292};
ram[38902] = {9'd95,10'd295};
ram[38903] = {9'd98,10'd298};
ram[38904] = {-9'd99,10'd301};
ram[38905] = {-9'd96,10'd304};
ram[38906] = {-9'd93,10'd307};
ram[38907] = {-9'd90,10'd311};
ram[38908] = {-9'd87,10'd314};
ram[38909] = {-9'd84,10'd317};
ram[38910] = {-9'd81,10'd320};
ram[38911] = {-9'd77,10'd323};
ram[38912] = {-9'd77,10'd323};
ram[38913] = {-9'd74,10'd326};
ram[38914] = {-9'd71,10'd329};
ram[38915] = {-9'd68,10'd333};
ram[38916] = {-9'd65,10'd336};
ram[38917] = {-9'd62,10'd339};
ram[38918] = {-9'd59,10'd342};
ram[38919] = {-9'd55,10'd345};
ram[38920] = {-9'd52,10'd348};
ram[38921] = {-9'd49,10'd351};
ram[38922] = {-9'd46,10'd354};
ram[38923] = {-9'd43,10'd358};
ram[38924] = {-9'd40,10'd361};
ram[38925] = {-9'd37,10'd364};
ram[38926] = {-9'd33,10'd367};
ram[38927] = {-9'd30,10'd370};
ram[38928] = {-9'd27,10'd373};
ram[38929] = {-9'd24,10'd376};
ram[38930] = {-9'd21,10'd380};
ram[38931] = {-9'd18,10'd383};
ram[38932] = {-9'd15,10'd386};
ram[38933] = {-9'd11,10'd389};
ram[38934] = {-9'd8,10'd392};
ram[38935] = {-9'd5,10'd395};
ram[38936] = {-9'd2,10'd398};
ram[38937] = {9'd1,-10'd399};
ram[38938] = {9'd4,-10'd396};
ram[38939] = {9'd7,-10'd393};
ram[38940] = {9'd10,-10'd390};
ram[38941] = {9'd14,-10'd387};
ram[38942] = {9'd17,-10'd384};
ram[38943] = {9'd20,-10'd381};
ram[38944] = {9'd23,-10'd377};
ram[38945] = {9'd26,-10'd374};
ram[38946] = {9'd29,-10'd371};
ram[38947] = {9'd32,-10'd368};
ram[38948] = {9'd36,-10'd365};
ram[38949] = {9'd39,-10'd362};
ram[38950] = {9'd42,-10'd359};
ram[38951] = {9'd45,-10'd355};
ram[38952] = {9'd48,-10'd352};
ram[38953] = {9'd51,-10'd349};
ram[38954] = {9'd54,-10'd346};
ram[38955] = {9'd58,-10'd343};
ram[38956] = {9'd61,-10'd340};
ram[38957] = {9'd64,-10'd337};
ram[38958] = {9'd67,-10'd334};
ram[38959] = {9'd70,-10'd330};
ram[38960] = {9'd73,-10'd327};
ram[38961] = {9'd76,-10'd324};
ram[38962] = {9'd80,-10'd321};
ram[38963] = {9'd83,-10'd318};
ram[38964] = {9'd86,-10'd315};
ram[38965] = {9'd89,-10'd312};
ram[38966] = {9'd92,-10'd308};
ram[38967] = {9'd95,-10'd305};
ram[38968] = {9'd98,-10'd302};
ram[38969] = {-9'd99,-10'd299};
ram[38970] = {-9'd96,-10'd296};
ram[38971] = {-9'd92,-10'd293};
ram[38972] = {-9'd89,-10'd290};
ram[38973] = {-9'd86,-10'd286};
ram[38974] = {-9'd83,-10'd283};
ram[38975] = {-9'd80,-10'd280};
ram[38976] = {-9'd77,-10'd277};
ram[38977] = {-9'd74,-10'd274};
ram[38978] = {-9'd70,-10'd271};
ram[38979] = {-9'd67,-10'd268};
ram[38980] = {-9'd64,-10'd264};
ram[38981] = {-9'd61,-10'd261};
ram[38982] = {-9'd58,-10'd258};
ram[38983] = {-9'd55,-10'd255};
ram[38984] = {-9'd52,-10'd252};
ram[38985] = {-9'd48,-10'd249};
ram[38986] = {-9'd45,-10'd246};
ram[38987] = {-9'd42,-10'd242};
ram[38988] = {-9'd39,-10'd239};
ram[38989] = {-9'd36,-10'd236};
ram[38990] = {-9'd33,-10'd233};
ram[38991] = {-9'd30,-10'd230};
ram[38992] = {-9'd26,-10'd227};
ram[38993] = {-9'd23,-10'd224};
ram[38994] = {-9'd20,-10'd220};
ram[38995] = {-9'd17,-10'd217};
ram[38996] = {-9'd14,-10'd214};
ram[38997] = {-9'd11,-10'd211};
ram[38998] = {-9'd8,-10'd208};
ram[38999] = {-9'd4,-10'd205};
ram[39000] = {-9'd1,-10'd202};
ram[39001] = {9'd2,-10'd198};
ram[39002] = {9'd5,-10'd195};
ram[39003] = {9'd8,-10'd192};
ram[39004] = {9'd11,-10'd189};
ram[39005] = {9'd14,-10'd186};
ram[39006] = {9'd18,-10'd183};
ram[39007] = {9'd21,-10'd180};
ram[39008] = {9'd24,-10'd176};
ram[39009] = {9'd27,-10'd173};
ram[39010] = {9'd30,-10'd170};
ram[39011] = {9'd33,-10'd167};
ram[39012] = {9'd36,-10'd164};
ram[39013] = {9'd40,-10'd161};
ram[39014] = {9'd43,-10'd158};
ram[39015] = {9'd46,-10'd154};
ram[39016] = {9'd49,-10'd151};
ram[39017] = {9'd52,-10'd148};
ram[39018] = {9'd55,-10'd145};
ram[39019] = {9'd58,-10'd142};
ram[39020] = {9'd62,-10'd139};
ram[39021] = {9'd65,-10'd136};
ram[39022] = {9'd68,-10'd132};
ram[39023] = {9'd71,-10'd129};
ram[39024] = {9'd74,-10'd126};
ram[39025] = {9'd77,-10'd123};
ram[39026] = {9'd80,-10'd120};
ram[39027] = {9'd84,-10'd117};
ram[39028] = {9'd87,-10'd114};
ram[39029] = {9'd90,-10'd110};
ram[39030] = {9'd93,-10'd107};
ram[39031] = {9'd96,-10'd104};
ram[39032] = {9'd99,-10'd101};
ram[39033] = {-9'd98,-10'd98};
ram[39034] = {-9'd95,-10'd95};
ram[39035] = {-9'd92,-10'd92};
ram[39036] = {-9'd88,-10'd88};
ram[39037] = {-9'd85,-10'd85};
ram[39038] = {-9'd82,-10'd82};
ram[39039] = {-9'd79,-10'd79};
ram[39040] = {-9'd79,-10'd79};
ram[39041] = {-9'd76,-10'd76};
ram[39042] = {-9'd73,-10'd73};
ram[39043] = {-9'd70,-10'd70};
ram[39044] = {-9'd66,-10'd66};
ram[39045] = {-9'd63,-10'd63};
ram[39046] = {-9'd60,-10'd60};
ram[39047] = {-9'd57,-10'd57};
ram[39048] = {-9'd54,-10'd54};
ram[39049] = {-9'd51,-10'd51};
ram[39050] = {-9'd48,-10'd48};
ram[39051] = {-9'd44,-10'd44};
ram[39052] = {-9'd41,-10'd41};
ram[39053] = {-9'd38,-10'd38};
ram[39054] = {-9'd35,-10'd35};
ram[39055] = {-9'd32,-10'd32};
ram[39056] = {-9'd29,-10'd29};
ram[39057] = {-9'd26,-10'd26};
ram[39058] = {-9'd22,-10'd22};
ram[39059] = {-9'd19,-10'd19};
ram[39060] = {-9'd16,-10'd16};
ram[39061] = {-9'd13,-10'd13};
ram[39062] = {-9'd10,-10'd10};
ram[39063] = {-9'd7,-10'd7};
ram[39064] = {-9'd4,-10'd4};
ram[39065] = {9'd0,10'd0};
ram[39066] = {9'd3,10'd3};
ram[39067] = {9'd6,10'd6};
ram[39068] = {9'd9,10'd9};
ram[39069] = {9'd12,10'd12};
ram[39070] = {9'd15,10'd15};
ram[39071] = {9'd18,10'd18};
ram[39072] = {9'd21,10'd21};
ram[39073] = {9'd25,10'd25};
ram[39074] = {9'd28,10'd28};
ram[39075] = {9'd31,10'd31};
ram[39076] = {9'd34,10'd34};
ram[39077] = {9'd37,10'd37};
ram[39078] = {9'd40,10'd40};
ram[39079] = {9'd43,10'd43};
ram[39080] = {9'd47,10'd47};
ram[39081] = {9'd50,10'd50};
ram[39082] = {9'd53,10'd53};
ram[39083] = {9'd56,10'd56};
ram[39084] = {9'd59,10'd59};
ram[39085] = {9'd62,10'd62};
ram[39086] = {9'd65,10'd65};
ram[39087] = {9'd69,10'd69};
ram[39088] = {9'd72,10'd72};
ram[39089] = {9'd75,10'd75};
ram[39090] = {9'd78,10'd78};
ram[39091] = {9'd81,10'd81};
ram[39092] = {9'd84,10'd84};
ram[39093] = {9'd87,10'd87};
ram[39094] = {9'd91,10'd91};
ram[39095] = {9'd94,10'd94};
ram[39096] = {9'd97,10'd97};
ram[39097] = {-9'd100,10'd100};
ram[39098] = {-9'd97,10'd103};
ram[39099] = {-9'd94,10'd106};
ram[39100] = {-9'd91,10'd109};
ram[39101] = {-9'd88,10'd113};
ram[39102] = {-9'd85,10'd116};
ram[39103] = {-9'd81,10'd119};
ram[39104] = {-9'd78,10'd122};
ram[39105] = {-9'd75,10'd125};
ram[39106] = {-9'd72,10'd128};
ram[39107] = {-9'd69,10'd131};
ram[39108] = {-9'd66,10'd135};
ram[39109] = {-9'd63,10'd138};
ram[39110] = {-9'd59,10'd141};
ram[39111] = {-9'd56,10'd144};
ram[39112] = {-9'd53,10'd147};
ram[39113] = {-9'd50,10'd150};
ram[39114] = {-9'd47,10'd153};
ram[39115] = {-9'd44,10'd157};
ram[39116] = {-9'd41,10'd160};
ram[39117] = {-9'd37,10'd163};
ram[39118] = {-9'd34,10'd166};
ram[39119] = {-9'd31,10'd169};
ram[39120] = {-9'd28,10'd172};
ram[39121] = {-9'd25,10'd175};
ram[39122] = {-9'd22,10'd179};
ram[39123] = {-9'd19,10'd182};
ram[39124] = {-9'd15,10'd185};
ram[39125] = {-9'd12,10'd188};
ram[39126] = {-9'd9,10'd191};
ram[39127] = {-9'd6,10'd194};
ram[39128] = {-9'd3,10'd197};
ram[39129] = {9'd0,10'd201};
ram[39130] = {9'd3,10'd204};
ram[39131] = {9'd7,10'd207};
ram[39132] = {9'd10,10'd210};
ram[39133] = {9'd13,10'd213};
ram[39134] = {9'd16,10'd216};
ram[39135] = {9'd19,10'd219};
ram[39136] = {9'd22,10'd223};
ram[39137] = {9'd25,10'd226};
ram[39138] = {9'd29,10'd229};
ram[39139] = {9'd32,10'd232};
ram[39140] = {9'd35,10'd235};
ram[39141] = {9'd38,10'd238};
ram[39142] = {9'd41,10'd241};
ram[39143] = {9'd44,10'd245};
ram[39144] = {9'd47,10'd248};
ram[39145] = {9'd51,10'd251};
ram[39146] = {9'd54,10'd254};
ram[39147] = {9'd57,10'd257};
ram[39148] = {9'd60,10'd260};
ram[39149] = {9'd63,10'd263};
ram[39150] = {9'd66,10'd267};
ram[39151] = {9'd69,10'd270};
ram[39152] = {9'd73,10'd273};
ram[39153] = {9'd76,10'd276};
ram[39154] = {9'd79,10'd279};
ram[39155] = {9'd82,10'd282};
ram[39156] = {9'd85,10'd285};
ram[39157] = {9'd88,10'd289};
ram[39158] = {9'd91,10'd292};
ram[39159] = {9'd95,10'd295};
ram[39160] = {9'd98,10'd298};
ram[39161] = {-9'd99,10'd301};
ram[39162] = {-9'd96,10'd304};
ram[39163] = {-9'd93,10'd307};
ram[39164] = {-9'd90,10'd311};
ram[39165] = {-9'd87,10'd314};
ram[39166] = {-9'd84,10'd317};
ram[39167] = {-9'd81,10'd320};
ram[39168] = {-9'd81,10'd320};
ram[39169] = {-9'd77,10'd323};
ram[39170] = {-9'd74,10'd326};
ram[39171] = {-9'd71,10'd329};
ram[39172] = {-9'd68,10'd333};
ram[39173] = {-9'd65,10'd336};
ram[39174] = {-9'd62,10'd339};
ram[39175] = {-9'd59,10'd342};
ram[39176] = {-9'd55,10'd345};
ram[39177] = {-9'd52,10'd348};
ram[39178] = {-9'd49,10'd351};
ram[39179] = {-9'd46,10'd354};
ram[39180] = {-9'd43,10'd358};
ram[39181] = {-9'd40,10'd361};
ram[39182] = {-9'd37,10'd364};
ram[39183] = {-9'd33,10'd367};
ram[39184] = {-9'd30,10'd370};
ram[39185] = {-9'd27,10'd373};
ram[39186] = {-9'd24,10'd376};
ram[39187] = {-9'd21,10'd380};
ram[39188] = {-9'd18,10'd383};
ram[39189] = {-9'd15,10'd386};
ram[39190] = {-9'd11,10'd389};
ram[39191] = {-9'd8,10'd392};
ram[39192] = {-9'd5,10'd395};
ram[39193] = {-9'd2,10'd398};
ram[39194] = {9'd1,-10'd399};
ram[39195] = {9'd4,-10'd396};
ram[39196] = {9'd7,-10'd393};
ram[39197] = {9'd10,-10'd390};
ram[39198] = {9'd14,-10'd387};
ram[39199] = {9'd17,-10'd384};
ram[39200] = {9'd20,-10'd381};
ram[39201] = {9'd23,-10'd377};
ram[39202] = {9'd26,-10'd374};
ram[39203] = {9'd29,-10'd371};
ram[39204] = {9'd32,-10'd368};
ram[39205] = {9'd36,-10'd365};
ram[39206] = {9'd39,-10'd362};
ram[39207] = {9'd42,-10'd359};
ram[39208] = {9'd45,-10'd355};
ram[39209] = {9'd48,-10'd352};
ram[39210] = {9'd51,-10'd349};
ram[39211] = {9'd54,-10'd346};
ram[39212] = {9'd58,-10'd343};
ram[39213] = {9'd61,-10'd340};
ram[39214] = {9'd64,-10'd337};
ram[39215] = {9'd67,-10'd334};
ram[39216] = {9'd70,-10'd330};
ram[39217] = {9'd73,-10'd327};
ram[39218] = {9'd76,-10'd324};
ram[39219] = {9'd80,-10'd321};
ram[39220] = {9'd83,-10'd318};
ram[39221] = {9'd86,-10'd315};
ram[39222] = {9'd89,-10'd312};
ram[39223] = {9'd92,-10'd308};
ram[39224] = {9'd95,-10'd305};
ram[39225] = {9'd98,-10'd302};
ram[39226] = {-9'd99,-10'd299};
ram[39227] = {-9'd96,-10'd296};
ram[39228] = {-9'd92,-10'd293};
ram[39229] = {-9'd89,-10'd290};
ram[39230] = {-9'd86,-10'd286};
ram[39231] = {-9'd83,-10'd283};
ram[39232] = {-9'd80,-10'd280};
ram[39233] = {-9'd77,-10'd277};
ram[39234] = {-9'd74,-10'd274};
ram[39235] = {-9'd70,-10'd271};
ram[39236] = {-9'd67,-10'd268};
ram[39237] = {-9'd64,-10'd264};
ram[39238] = {-9'd61,-10'd261};
ram[39239] = {-9'd58,-10'd258};
ram[39240] = {-9'd55,-10'd255};
ram[39241] = {-9'd52,-10'd252};
ram[39242] = {-9'd48,-10'd249};
ram[39243] = {-9'd45,-10'd246};
ram[39244] = {-9'd42,-10'd242};
ram[39245] = {-9'd39,-10'd239};
ram[39246] = {-9'd36,-10'd236};
ram[39247] = {-9'd33,-10'd233};
ram[39248] = {-9'd30,-10'd230};
ram[39249] = {-9'd26,-10'd227};
ram[39250] = {-9'd23,-10'd224};
ram[39251] = {-9'd20,-10'd220};
ram[39252] = {-9'd17,-10'd217};
ram[39253] = {-9'd14,-10'd214};
ram[39254] = {-9'd11,-10'd211};
ram[39255] = {-9'd8,-10'd208};
ram[39256] = {-9'd4,-10'd205};
ram[39257] = {-9'd1,-10'd202};
ram[39258] = {9'd2,-10'd198};
ram[39259] = {9'd5,-10'd195};
ram[39260] = {9'd8,-10'd192};
ram[39261] = {9'd11,-10'd189};
ram[39262] = {9'd14,-10'd186};
ram[39263] = {9'd18,-10'd183};
ram[39264] = {9'd21,-10'd180};
ram[39265] = {9'd24,-10'd176};
ram[39266] = {9'd27,-10'd173};
ram[39267] = {9'd30,-10'd170};
ram[39268] = {9'd33,-10'd167};
ram[39269] = {9'd36,-10'd164};
ram[39270] = {9'd40,-10'd161};
ram[39271] = {9'd43,-10'd158};
ram[39272] = {9'd46,-10'd154};
ram[39273] = {9'd49,-10'd151};
ram[39274] = {9'd52,-10'd148};
ram[39275] = {9'd55,-10'd145};
ram[39276] = {9'd58,-10'd142};
ram[39277] = {9'd62,-10'd139};
ram[39278] = {9'd65,-10'd136};
ram[39279] = {9'd68,-10'd132};
ram[39280] = {9'd71,-10'd129};
ram[39281] = {9'd74,-10'd126};
ram[39282] = {9'd77,-10'd123};
ram[39283] = {9'd80,-10'd120};
ram[39284] = {9'd84,-10'd117};
ram[39285] = {9'd87,-10'd114};
ram[39286] = {9'd90,-10'd110};
ram[39287] = {9'd93,-10'd107};
ram[39288] = {9'd96,-10'd104};
ram[39289] = {9'd99,-10'd101};
ram[39290] = {-9'd98,-10'd98};
ram[39291] = {-9'd95,-10'd95};
ram[39292] = {-9'd92,-10'd92};
ram[39293] = {-9'd88,-10'd88};
ram[39294] = {-9'd85,-10'd85};
ram[39295] = {-9'd82,-10'd82};
ram[39296] = {-9'd82,-10'd82};
ram[39297] = {-9'd79,-10'd79};
ram[39298] = {-9'd76,-10'd76};
ram[39299] = {-9'd73,-10'd73};
ram[39300] = {-9'd70,-10'd70};
ram[39301] = {-9'd66,-10'd66};
ram[39302] = {-9'd63,-10'd63};
ram[39303] = {-9'd60,-10'd60};
ram[39304] = {-9'd57,-10'd57};
ram[39305] = {-9'd54,-10'd54};
ram[39306] = {-9'd51,-10'd51};
ram[39307] = {-9'd48,-10'd48};
ram[39308] = {-9'd44,-10'd44};
ram[39309] = {-9'd41,-10'd41};
ram[39310] = {-9'd38,-10'd38};
ram[39311] = {-9'd35,-10'd35};
ram[39312] = {-9'd32,-10'd32};
ram[39313] = {-9'd29,-10'd29};
ram[39314] = {-9'd26,-10'd26};
ram[39315] = {-9'd22,-10'd22};
ram[39316] = {-9'd19,-10'd19};
ram[39317] = {-9'd16,-10'd16};
ram[39318] = {-9'd13,-10'd13};
ram[39319] = {-9'd10,-10'd10};
ram[39320] = {-9'd7,-10'd7};
ram[39321] = {-9'd4,-10'd4};
ram[39322] = {9'd0,10'd0};
ram[39323] = {9'd3,10'd3};
ram[39324] = {9'd6,10'd6};
ram[39325] = {9'd9,10'd9};
ram[39326] = {9'd12,10'd12};
ram[39327] = {9'd15,10'd15};
ram[39328] = {9'd18,10'd18};
ram[39329] = {9'd21,10'd21};
ram[39330] = {9'd25,10'd25};
ram[39331] = {9'd28,10'd28};
ram[39332] = {9'd31,10'd31};
ram[39333] = {9'd34,10'd34};
ram[39334] = {9'd37,10'd37};
ram[39335] = {9'd40,10'd40};
ram[39336] = {9'd43,10'd43};
ram[39337] = {9'd47,10'd47};
ram[39338] = {9'd50,10'd50};
ram[39339] = {9'd53,10'd53};
ram[39340] = {9'd56,10'd56};
ram[39341] = {9'd59,10'd59};
ram[39342] = {9'd62,10'd62};
ram[39343] = {9'd65,10'd65};
ram[39344] = {9'd69,10'd69};
ram[39345] = {9'd72,10'd72};
ram[39346] = {9'd75,10'd75};
ram[39347] = {9'd78,10'd78};
ram[39348] = {9'd81,10'd81};
ram[39349] = {9'd84,10'd84};
ram[39350] = {9'd87,10'd87};
ram[39351] = {9'd91,10'd91};
ram[39352] = {9'd94,10'd94};
ram[39353] = {9'd97,10'd97};
ram[39354] = {-9'd100,10'd100};
ram[39355] = {-9'd97,10'd103};
ram[39356] = {-9'd94,10'd106};
ram[39357] = {-9'd91,10'd109};
ram[39358] = {-9'd88,10'd113};
ram[39359] = {-9'd85,10'd116};
ram[39360] = {-9'd81,10'd119};
ram[39361] = {-9'd78,10'd122};
ram[39362] = {-9'd75,10'd125};
ram[39363] = {-9'd72,10'd128};
ram[39364] = {-9'd69,10'd131};
ram[39365] = {-9'd66,10'd135};
ram[39366] = {-9'd63,10'd138};
ram[39367] = {-9'd59,10'd141};
ram[39368] = {-9'd56,10'd144};
ram[39369] = {-9'd53,10'd147};
ram[39370] = {-9'd50,10'd150};
ram[39371] = {-9'd47,10'd153};
ram[39372] = {-9'd44,10'd157};
ram[39373] = {-9'd41,10'd160};
ram[39374] = {-9'd37,10'd163};
ram[39375] = {-9'd34,10'd166};
ram[39376] = {-9'd31,10'd169};
ram[39377] = {-9'd28,10'd172};
ram[39378] = {-9'd25,10'd175};
ram[39379] = {-9'd22,10'd179};
ram[39380] = {-9'd19,10'd182};
ram[39381] = {-9'd15,10'd185};
ram[39382] = {-9'd12,10'd188};
ram[39383] = {-9'd9,10'd191};
ram[39384] = {-9'd6,10'd194};
ram[39385] = {-9'd3,10'd197};
ram[39386] = {9'd0,10'd201};
ram[39387] = {9'd3,10'd204};
ram[39388] = {9'd7,10'd207};
ram[39389] = {9'd10,10'd210};
ram[39390] = {9'd13,10'd213};
ram[39391] = {9'd16,10'd216};
ram[39392] = {9'd19,10'd219};
ram[39393] = {9'd22,10'd223};
ram[39394] = {9'd25,10'd226};
ram[39395] = {9'd29,10'd229};
ram[39396] = {9'd32,10'd232};
ram[39397] = {9'd35,10'd235};
ram[39398] = {9'd38,10'd238};
ram[39399] = {9'd41,10'd241};
ram[39400] = {9'd44,10'd245};
ram[39401] = {9'd47,10'd248};
ram[39402] = {9'd51,10'd251};
ram[39403] = {9'd54,10'd254};
ram[39404] = {9'd57,10'd257};
ram[39405] = {9'd60,10'd260};
ram[39406] = {9'd63,10'd263};
ram[39407] = {9'd66,10'd267};
ram[39408] = {9'd69,10'd270};
ram[39409] = {9'd73,10'd273};
ram[39410] = {9'd76,10'd276};
ram[39411] = {9'd79,10'd279};
ram[39412] = {9'd82,10'd282};
ram[39413] = {9'd85,10'd285};
ram[39414] = {9'd88,10'd289};
ram[39415] = {9'd91,10'd292};
ram[39416] = {9'd95,10'd295};
ram[39417] = {9'd98,10'd298};
ram[39418] = {-9'd99,10'd301};
ram[39419] = {-9'd96,10'd304};
ram[39420] = {-9'd93,10'd307};
ram[39421] = {-9'd90,10'd311};
ram[39422] = {-9'd87,10'd314};
ram[39423] = {-9'd84,10'd317};
ram[39424] = {-9'd84,10'd317};
ram[39425] = {-9'd81,10'd320};
ram[39426] = {-9'd77,10'd323};
ram[39427] = {-9'd74,10'd326};
ram[39428] = {-9'd71,10'd329};
ram[39429] = {-9'd68,10'd333};
ram[39430] = {-9'd65,10'd336};
ram[39431] = {-9'd62,10'd339};
ram[39432] = {-9'd59,10'd342};
ram[39433] = {-9'd55,10'd345};
ram[39434] = {-9'd52,10'd348};
ram[39435] = {-9'd49,10'd351};
ram[39436] = {-9'd46,10'd354};
ram[39437] = {-9'd43,10'd358};
ram[39438] = {-9'd40,10'd361};
ram[39439] = {-9'd37,10'd364};
ram[39440] = {-9'd33,10'd367};
ram[39441] = {-9'd30,10'd370};
ram[39442] = {-9'd27,10'd373};
ram[39443] = {-9'd24,10'd376};
ram[39444] = {-9'd21,10'd380};
ram[39445] = {-9'd18,10'd383};
ram[39446] = {-9'd15,10'd386};
ram[39447] = {-9'd11,10'd389};
ram[39448] = {-9'd8,10'd392};
ram[39449] = {-9'd5,10'd395};
ram[39450] = {-9'd2,10'd398};
ram[39451] = {9'd1,-10'd399};
ram[39452] = {9'd4,-10'd396};
ram[39453] = {9'd7,-10'd393};
ram[39454] = {9'd10,-10'd390};
ram[39455] = {9'd14,-10'd387};
ram[39456] = {9'd17,-10'd384};
ram[39457] = {9'd20,-10'd381};
ram[39458] = {9'd23,-10'd377};
ram[39459] = {9'd26,-10'd374};
ram[39460] = {9'd29,-10'd371};
ram[39461] = {9'd32,-10'd368};
ram[39462] = {9'd36,-10'd365};
ram[39463] = {9'd39,-10'd362};
ram[39464] = {9'd42,-10'd359};
ram[39465] = {9'd45,-10'd355};
ram[39466] = {9'd48,-10'd352};
ram[39467] = {9'd51,-10'd349};
ram[39468] = {9'd54,-10'd346};
ram[39469] = {9'd58,-10'd343};
ram[39470] = {9'd61,-10'd340};
ram[39471] = {9'd64,-10'd337};
ram[39472] = {9'd67,-10'd334};
ram[39473] = {9'd70,-10'd330};
ram[39474] = {9'd73,-10'd327};
ram[39475] = {9'd76,-10'd324};
ram[39476] = {9'd80,-10'd321};
ram[39477] = {9'd83,-10'd318};
ram[39478] = {9'd86,-10'd315};
ram[39479] = {9'd89,-10'd312};
ram[39480] = {9'd92,-10'd308};
ram[39481] = {9'd95,-10'd305};
ram[39482] = {9'd98,-10'd302};
ram[39483] = {-9'd99,-10'd299};
ram[39484] = {-9'd96,-10'd296};
ram[39485] = {-9'd92,-10'd293};
ram[39486] = {-9'd89,-10'd290};
ram[39487] = {-9'd86,-10'd286};
ram[39488] = {-9'd83,-10'd283};
ram[39489] = {-9'd80,-10'd280};
ram[39490] = {-9'd77,-10'd277};
ram[39491] = {-9'd74,-10'd274};
ram[39492] = {-9'd70,-10'd271};
ram[39493] = {-9'd67,-10'd268};
ram[39494] = {-9'd64,-10'd264};
ram[39495] = {-9'd61,-10'd261};
ram[39496] = {-9'd58,-10'd258};
ram[39497] = {-9'd55,-10'd255};
ram[39498] = {-9'd52,-10'd252};
ram[39499] = {-9'd48,-10'd249};
ram[39500] = {-9'd45,-10'd246};
ram[39501] = {-9'd42,-10'd242};
ram[39502] = {-9'd39,-10'd239};
ram[39503] = {-9'd36,-10'd236};
ram[39504] = {-9'd33,-10'd233};
ram[39505] = {-9'd30,-10'd230};
ram[39506] = {-9'd26,-10'd227};
ram[39507] = {-9'd23,-10'd224};
ram[39508] = {-9'd20,-10'd220};
ram[39509] = {-9'd17,-10'd217};
ram[39510] = {-9'd14,-10'd214};
ram[39511] = {-9'd11,-10'd211};
ram[39512] = {-9'd8,-10'd208};
ram[39513] = {-9'd4,-10'd205};
ram[39514] = {-9'd1,-10'd202};
ram[39515] = {9'd2,-10'd198};
ram[39516] = {9'd5,-10'd195};
ram[39517] = {9'd8,-10'd192};
ram[39518] = {9'd11,-10'd189};
ram[39519] = {9'd14,-10'd186};
ram[39520] = {9'd18,-10'd183};
ram[39521] = {9'd21,-10'd180};
ram[39522] = {9'd24,-10'd176};
ram[39523] = {9'd27,-10'd173};
ram[39524] = {9'd30,-10'd170};
ram[39525] = {9'd33,-10'd167};
ram[39526] = {9'd36,-10'd164};
ram[39527] = {9'd40,-10'd161};
ram[39528] = {9'd43,-10'd158};
ram[39529] = {9'd46,-10'd154};
ram[39530] = {9'd49,-10'd151};
ram[39531] = {9'd52,-10'd148};
ram[39532] = {9'd55,-10'd145};
ram[39533] = {9'd58,-10'd142};
ram[39534] = {9'd62,-10'd139};
ram[39535] = {9'd65,-10'd136};
ram[39536] = {9'd68,-10'd132};
ram[39537] = {9'd71,-10'd129};
ram[39538] = {9'd74,-10'd126};
ram[39539] = {9'd77,-10'd123};
ram[39540] = {9'd80,-10'd120};
ram[39541] = {9'd84,-10'd117};
ram[39542] = {9'd87,-10'd114};
ram[39543] = {9'd90,-10'd110};
ram[39544] = {9'd93,-10'd107};
ram[39545] = {9'd96,-10'd104};
ram[39546] = {9'd99,-10'd101};
ram[39547] = {-9'd98,-10'd98};
ram[39548] = {-9'd95,-10'd95};
ram[39549] = {-9'd92,-10'd92};
ram[39550] = {-9'd88,-10'd88};
ram[39551] = {-9'd85,-10'd85};
ram[39552] = {-9'd85,-10'd85};
ram[39553] = {-9'd82,-10'd82};
ram[39554] = {-9'd79,-10'd79};
ram[39555] = {-9'd76,-10'd76};
ram[39556] = {-9'd73,-10'd73};
ram[39557] = {-9'd70,-10'd70};
ram[39558] = {-9'd66,-10'd66};
ram[39559] = {-9'd63,-10'd63};
ram[39560] = {-9'd60,-10'd60};
ram[39561] = {-9'd57,-10'd57};
ram[39562] = {-9'd54,-10'd54};
ram[39563] = {-9'd51,-10'd51};
ram[39564] = {-9'd48,-10'd48};
ram[39565] = {-9'd44,-10'd44};
ram[39566] = {-9'd41,-10'd41};
ram[39567] = {-9'd38,-10'd38};
ram[39568] = {-9'd35,-10'd35};
ram[39569] = {-9'd32,-10'd32};
ram[39570] = {-9'd29,-10'd29};
ram[39571] = {-9'd26,-10'd26};
ram[39572] = {-9'd22,-10'd22};
ram[39573] = {-9'd19,-10'd19};
ram[39574] = {-9'd16,-10'd16};
ram[39575] = {-9'd13,-10'd13};
ram[39576] = {-9'd10,-10'd10};
ram[39577] = {-9'd7,-10'd7};
ram[39578] = {-9'd4,-10'd4};
ram[39579] = {9'd0,10'd0};
ram[39580] = {9'd3,10'd3};
ram[39581] = {9'd6,10'd6};
ram[39582] = {9'd9,10'd9};
ram[39583] = {9'd12,10'd12};
ram[39584] = {9'd15,10'd15};
ram[39585] = {9'd18,10'd18};
ram[39586] = {9'd21,10'd21};
ram[39587] = {9'd25,10'd25};
ram[39588] = {9'd28,10'd28};
ram[39589] = {9'd31,10'd31};
ram[39590] = {9'd34,10'd34};
ram[39591] = {9'd37,10'd37};
ram[39592] = {9'd40,10'd40};
ram[39593] = {9'd43,10'd43};
ram[39594] = {9'd47,10'd47};
ram[39595] = {9'd50,10'd50};
ram[39596] = {9'd53,10'd53};
ram[39597] = {9'd56,10'd56};
ram[39598] = {9'd59,10'd59};
ram[39599] = {9'd62,10'd62};
ram[39600] = {9'd65,10'd65};
ram[39601] = {9'd69,10'd69};
ram[39602] = {9'd72,10'd72};
ram[39603] = {9'd75,10'd75};
ram[39604] = {9'd78,10'd78};
ram[39605] = {9'd81,10'd81};
ram[39606] = {9'd84,10'd84};
ram[39607] = {9'd87,10'd87};
ram[39608] = {9'd91,10'd91};
ram[39609] = {9'd94,10'd94};
ram[39610] = {9'd97,10'd97};
ram[39611] = {-9'd100,10'd100};
ram[39612] = {-9'd97,10'd103};
ram[39613] = {-9'd94,10'd106};
ram[39614] = {-9'd91,10'd109};
ram[39615] = {-9'd88,10'd113};
ram[39616] = {-9'd85,10'd116};
ram[39617] = {-9'd81,10'd119};
ram[39618] = {-9'd78,10'd122};
ram[39619] = {-9'd75,10'd125};
ram[39620] = {-9'd72,10'd128};
ram[39621] = {-9'd69,10'd131};
ram[39622] = {-9'd66,10'd135};
ram[39623] = {-9'd63,10'd138};
ram[39624] = {-9'd59,10'd141};
ram[39625] = {-9'd56,10'd144};
ram[39626] = {-9'd53,10'd147};
ram[39627] = {-9'd50,10'd150};
ram[39628] = {-9'd47,10'd153};
ram[39629] = {-9'd44,10'd157};
ram[39630] = {-9'd41,10'd160};
ram[39631] = {-9'd37,10'd163};
ram[39632] = {-9'd34,10'd166};
ram[39633] = {-9'd31,10'd169};
ram[39634] = {-9'd28,10'd172};
ram[39635] = {-9'd25,10'd175};
ram[39636] = {-9'd22,10'd179};
ram[39637] = {-9'd19,10'd182};
ram[39638] = {-9'd15,10'd185};
ram[39639] = {-9'd12,10'd188};
ram[39640] = {-9'd9,10'd191};
ram[39641] = {-9'd6,10'd194};
ram[39642] = {-9'd3,10'd197};
ram[39643] = {9'd0,10'd201};
ram[39644] = {9'd3,10'd204};
ram[39645] = {9'd7,10'd207};
ram[39646] = {9'd10,10'd210};
ram[39647] = {9'd13,10'd213};
ram[39648] = {9'd16,10'd216};
ram[39649] = {9'd19,10'd219};
ram[39650] = {9'd22,10'd223};
ram[39651] = {9'd25,10'd226};
ram[39652] = {9'd29,10'd229};
ram[39653] = {9'd32,10'd232};
ram[39654] = {9'd35,10'd235};
ram[39655] = {9'd38,10'd238};
ram[39656] = {9'd41,10'd241};
ram[39657] = {9'd44,10'd245};
ram[39658] = {9'd47,10'd248};
ram[39659] = {9'd51,10'd251};
ram[39660] = {9'd54,10'd254};
ram[39661] = {9'd57,10'd257};
ram[39662] = {9'd60,10'd260};
ram[39663] = {9'd63,10'd263};
ram[39664] = {9'd66,10'd267};
ram[39665] = {9'd69,10'd270};
ram[39666] = {9'd73,10'd273};
ram[39667] = {9'd76,10'd276};
ram[39668] = {9'd79,10'd279};
ram[39669] = {9'd82,10'd282};
ram[39670] = {9'd85,10'd285};
ram[39671] = {9'd88,10'd289};
ram[39672] = {9'd91,10'd292};
ram[39673] = {9'd95,10'd295};
ram[39674] = {9'd98,10'd298};
ram[39675] = {-9'd99,10'd301};
ram[39676] = {-9'd96,10'd304};
ram[39677] = {-9'd93,10'd307};
ram[39678] = {-9'd90,10'd311};
ram[39679] = {-9'd87,10'd314};
ram[39680] = {-9'd87,10'd314};
ram[39681] = {-9'd84,10'd317};
ram[39682] = {-9'd81,10'd320};
ram[39683] = {-9'd77,10'd323};
ram[39684] = {-9'd74,10'd326};
ram[39685] = {-9'd71,10'd329};
ram[39686] = {-9'd68,10'd333};
ram[39687] = {-9'd65,10'd336};
ram[39688] = {-9'd62,10'd339};
ram[39689] = {-9'd59,10'd342};
ram[39690] = {-9'd55,10'd345};
ram[39691] = {-9'd52,10'd348};
ram[39692] = {-9'd49,10'd351};
ram[39693] = {-9'd46,10'd354};
ram[39694] = {-9'd43,10'd358};
ram[39695] = {-9'd40,10'd361};
ram[39696] = {-9'd37,10'd364};
ram[39697] = {-9'd33,10'd367};
ram[39698] = {-9'd30,10'd370};
ram[39699] = {-9'd27,10'd373};
ram[39700] = {-9'd24,10'd376};
ram[39701] = {-9'd21,10'd380};
ram[39702] = {-9'd18,10'd383};
ram[39703] = {-9'd15,10'd386};
ram[39704] = {-9'd11,10'd389};
ram[39705] = {-9'd8,10'd392};
ram[39706] = {-9'd5,10'd395};
ram[39707] = {-9'd2,10'd398};
ram[39708] = {9'd1,-10'd399};
ram[39709] = {9'd4,-10'd396};
ram[39710] = {9'd7,-10'd393};
ram[39711] = {9'd10,-10'd390};
ram[39712] = {9'd14,-10'd387};
ram[39713] = {9'd17,-10'd384};
ram[39714] = {9'd20,-10'd381};
ram[39715] = {9'd23,-10'd377};
ram[39716] = {9'd26,-10'd374};
ram[39717] = {9'd29,-10'd371};
ram[39718] = {9'd32,-10'd368};
ram[39719] = {9'd36,-10'd365};
ram[39720] = {9'd39,-10'd362};
ram[39721] = {9'd42,-10'd359};
ram[39722] = {9'd45,-10'd355};
ram[39723] = {9'd48,-10'd352};
ram[39724] = {9'd51,-10'd349};
ram[39725] = {9'd54,-10'd346};
ram[39726] = {9'd58,-10'd343};
ram[39727] = {9'd61,-10'd340};
ram[39728] = {9'd64,-10'd337};
ram[39729] = {9'd67,-10'd334};
ram[39730] = {9'd70,-10'd330};
ram[39731] = {9'd73,-10'd327};
ram[39732] = {9'd76,-10'd324};
ram[39733] = {9'd80,-10'd321};
ram[39734] = {9'd83,-10'd318};
ram[39735] = {9'd86,-10'd315};
ram[39736] = {9'd89,-10'd312};
ram[39737] = {9'd92,-10'd308};
ram[39738] = {9'd95,-10'd305};
ram[39739] = {9'd98,-10'd302};
ram[39740] = {-9'd99,-10'd299};
ram[39741] = {-9'd96,-10'd296};
ram[39742] = {-9'd92,-10'd293};
ram[39743] = {-9'd89,-10'd290};
ram[39744] = {-9'd86,-10'd286};
ram[39745] = {-9'd83,-10'd283};
ram[39746] = {-9'd80,-10'd280};
ram[39747] = {-9'd77,-10'd277};
ram[39748] = {-9'd74,-10'd274};
ram[39749] = {-9'd70,-10'd271};
ram[39750] = {-9'd67,-10'd268};
ram[39751] = {-9'd64,-10'd264};
ram[39752] = {-9'd61,-10'd261};
ram[39753] = {-9'd58,-10'd258};
ram[39754] = {-9'd55,-10'd255};
ram[39755] = {-9'd52,-10'd252};
ram[39756] = {-9'd48,-10'd249};
ram[39757] = {-9'd45,-10'd246};
ram[39758] = {-9'd42,-10'd242};
ram[39759] = {-9'd39,-10'd239};
ram[39760] = {-9'd36,-10'd236};
ram[39761] = {-9'd33,-10'd233};
ram[39762] = {-9'd30,-10'd230};
ram[39763] = {-9'd26,-10'd227};
ram[39764] = {-9'd23,-10'd224};
ram[39765] = {-9'd20,-10'd220};
ram[39766] = {-9'd17,-10'd217};
ram[39767] = {-9'd14,-10'd214};
ram[39768] = {-9'd11,-10'd211};
ram[39769] = {-9'd8,-10'd208};
ram[39770] = {-9'd4,-10'd205};
ram[39771] = {-9'd1,-10'd202};
ram[39772] = {9'd2,-10'd198};
ram[39773] = {9'd5,-10'd195};
ram[39774] = {9'd8,-10'd192};
ram[39775] = {9'd11,-10'd189};
ram[39776] = {9'd14,-10'd186};
ram[39777] = {9'd18,-10'd183};
ram[39778] = {9'd21,-10'd180};
ram[39779] = {9'd24,-10'd176};
ram[39780] = {9'd27,-10'd173};
ram[39781] = {9'd30,-10'd170};
ram[39782] = {9'd33,-10'd167};
ram[39783] = {9'd36,-10'd164};
ram[39784] = {9'd40,-10'd161};
ram[39785] = {9'd43,-10'd158};
ram[39786] = {9'd46,-10'd154};
ram[39787] = {9'd49,-10'd151};
ram[39788] = {9'd52,-10'd148};
ram[39789] = {9'd55,-10'd145};
ram[39790] = {9'd58,-10'd142};
ram[39791] = {9'd62,-10'd139};
ram[39792] = {9'd65,-10'd136};
ram[39793] = {9'd68,-10'd132};
ram[39794] = {9'd71,-10'd129};
ram[39795] = {9'd74,-10'd126};
ram[39796] = {9'd77,-10'd123};
ram[39797] = {9'd80,-10'd120};
ram[39798] = {9'd84,-10'd117};
ram[39799] = {9'd87,-10'd114};
ram[39800] = {9'd90,-10'd110};
ram[39801] = {9'd93,-10'd107};
ram[39802] = {9'd96,-10'd104};
ram[39803] = {9'd99,-10'd101};
ram[39804] = {-9'd98,-10'd98};
ram[39805] = {-9'd95,-10'd95};
ram[39806] = {-9'd92,-10'd92};
ram[39807] = {-9'd88,-10'd88};
ram[39808] = {-9'd88,-10'd88};
ram[39809] = {-9'd85,-10'd85};
ram[39810] = {-9'd82,-10'd82};
ram[39811] = {-9'd79,-10'd79};
ram[39812] = {-9'd76,-10'd76};
ram[39813] = {-9'd73,-10'd73};
ram[39814] = {-9'd70,-10'd70};
ram[39815] = {-9'd66,-10'd66};
ram[39816] = {-9'd63,-10'd63};
ram[39817] = {-9'd60,-10'd60};
ram[39818] = {-9'd57,-10'd57};
ram[39819] = {-9'd54,-10'd54};
ram[39820] = {-9'd51,-10'd51};
ram[39821] = {-9'd48,-10'd48};
ram[39822] = {-9'd44,-10'd44};
ram[39823] = {-9'd41,-10'd41};
ram[39824] = {-9'd38,-10'd38};
ram[39825] = {-9'd35,-10'd35};
ram[39826] = {-9'd32,-10'd32};
ram[39827] = {-9'd29,-10'd29};
ram[39828] = {-9'd26,-10'd26};
ram[39829] = {-9'd22,-10'd22};
ram[39830] = {-9'd19,-10'd19};
ram[39831] = {-9'd16,-10'd16};
ram[39832] = {-9'd13,-10'd13};
ram[39833] = {-9'd10,-10'd10};
ram[39834] = {-9'd7,-10'd7};
ram[39835] = {-9'd4,-10'd4};
ram[39836] = {9'd0,10'd0};
ram[39837] = {9'd3,10'd3};
ram[39838] = {9'd6,10'd6};
ram[39839] = {9'd9,10'd9};
ram[39840] = {9'd12,10'd12};
ram[39841] = {9'd15,10'd15};
ram[39842] = {9'd18,10'd18};
ram[39843] = {9'd21,10'd21};
ram[39844] = {9'd25,10'd25};
ram[39845] = {9'd28,10'd28};
ram[39846] = {9'd31,10'd31};
ram[39847] = {9'd34,10'd34};
ram[39848] = {9'd37,10'd37};
ram[39849] = {9'd40,10'd40};
ram[39850] = {9'd43,10'd43};
ram[39851] = {9'd47,10'd47};
ram[39852] = {9'd50,10'd50};
ram[39853] = {9'd53,10'd53};
ram[39854] = {9'd56,10'd56};
ram[39855] = {9'd59,10'd59};
ram[39856] = {9'd62,10'd62};
ram[39857] = {9'd65,10'd65};
ram[39858] = {9'd69,10'd69};
ram[39859] = {9'd72,10'd72};
ram[39860] = {9'd75,10'd75};
ram[39861] = {9'd78,10'd78};
ram[39862] = {9'd81,10'd81};
ram[39863] = {9'd84,10'd84};
ram[39864] = {9'd87,10'd87};
ram[39865] = {9'd91,10'd91};
ram[39866] = {9'd94,10'd94};
ram[39867] = {9'd97,10'd97};
ram[39868] = {-9'd100,10'd100};
ram[39869] = {-9'd97,10'd103};
ram[39870] = {-9'd94,10'd106};
ram[39871] = {-9'd91,10'd109};
ram[39872] = {-9'd88,10'd113};
ram[39873] = {-9'd85,10'd116};
ram[39874] = {-9'd81,10'd119};
ram[39875] = {-9'd78,10'd122};
ram[39876] = {-9'd75,10'd125};
ram[39877] = {-9'd72,10'd128};
ram[39878] = {-9'd69,10'd131};
ram[39879] = {-9'd66,10'd135};
ram[39880] = {-9'd63,10'd138};
ram[39881] = {-9'd59,10'd141};
ram[39882] = {-9'd56,10'd144};
ram[39883] = {-9'd53,10'd147};
ram[39884] = {-9'd50,10'd150};
ram[39885] = {-9'd47,10'd153};
ram[39886] = {-9'd44,10'd157};
ram[39887] = {-9'd41,10'd160};
ram[39888] = {-9'd37,10'd163};
ram[39889] = {-9'd34,10'd166};
ram[39890] = {-9'd31,10'd169};
ram[39891] = {-9'd28,10'd172};
ram[39892] = {-9'd25,10'd175};
ram[39893] = {-9'd22,10'd179};
ram[39894] = {-9'd19,10'd182};
ram[39895] = {-9'd15,10'd185};
ram[39896] = {-9'd12,10'd188};
ram[39897] = {-9'd9,10'd191};
ram[39898] = {-9'd6,10'd194};
ram[39899] = {-9'd3,10'd197};
ram[39900] = {9'd0,10'd201};
ram[39901] = {9'd3,10'd204};
ram[39902] = {9'd7,10'd207};
ram[39903] = {9'd10,10'd210};
ram[39904] = {9'd13,10'd213};
ram[39905] = {9'd16,10'd216};
ram[39906] = {9'd19,10'd219};
ram[39907] = {9'd22,10'd223};
ram[39908] = {9'd25,10'd226};
ram[39909] = {9'd29,10'd229};
ram[39910] = {9'd32,10'd232};
ram[39911] = {9'd35,10'd235};
ram[39912] = {9'd38,10'd238};
ram[39913] = {9'd41,10'd241};
ram[39914] = {9'd44,10'd245};
ram[39915] = {9'd47,10'd248};
ram[39916] = {9'd51,10'd251};
ram[39917] = {9'd54,10'd254};
ram[39918] = {9'd57,10'd257};
ram[39919] = {9'd60,10'd260};
ram[39920] = {9'd63,10'd263};
ram[39921] = {9'd66,10'd267};
ram[39922] = {9'd69,10'd270};
ram[39923] = {9'd73,10'd273};
ram[39924] = {9'd76,10'd276};
ram[39925] = {9'd79,10'd279};
ram[39926] = {9'd82,10'd282};
ram[39927] = {9'd85,10'd285};
ram[39928] = {9'd88,10'd289};
ram[39929] = {9'd91,10'd292};
ram[39930] = {9'd95,10'd295};
ram[39931] = {9'd98,10'd298};
ram[39932] = {-9'd99,10'd301};
ram[39933] = {-9'd96,10'd304};
ram[39934] = {-9'd93,10'd307};
ram[39935] = {-9'd90,10'd311};
ram[39936] = {-9'd90,10'd311};
ram[39937] = {-9'd87,10'd314};
ram[39938] = {-9'd84,10'd317};
ram[39939] = {-9'd81,10'd320};
ram[39940] = {-9'd77,10'd323};
ram[39941] = {-9'd74,10'd326};
ram[39942] = {-9'd71,10'd329};
ram[39943] = {-9'd68,10'd333};
ram[39944] = {-9'd65,10'd336};
ram[39945] = {-9'd62,10'd339};
ram[39946] = {-9'd59,10'd342};
ram[39947] = {-9'd55,10'd345};
ram[39948] = {-9'd52,10'd348};
ram[39949] = {-9'd49,10'd351};
ram[39950] = {-9'd46,10'd354};
ram[39951] = {-9'd43,10'd358};
ram[39952] = {-9'd40,10'd361};
ram[39953] = {-9'd37,10'd364};
ram[39954] = {-9'd33,10'd367};
ram[39955] = {-9'd30,10'd370};
ram[39956] = {-9'd27,10'd373};
ram[39957] = {-9'd24,10'd376};
ram[39958] = {-9'd21,10'd380};
ram[39959] = {-9'd18,10'd383};
ram[39960] = {-9'd15,10'd386};
ram[39961] = {-9'd11,10'd389};
ram[39962] = {-9'd8,10'd392};
ram[39963] = {-9'd5,10'd395};
ram[39964] = {-9'd2,10'd398};
ram[39965] = {9'd1,-10'd399};
ram[39966] = {9'd4,-10'd396};
ram[39967] = {9'd7,-10'd393};
ram[39968] = {9'd10,-10'd390};
ram[39969] = {9'd14,-10'd387};
ram[39970] = {9'd17,-10'd384};
ram[39971] = {9'd20,-10'd381};
ram[39972] = {9'd23,-10'd377};
ram[39973] = {9'd26,-10'd374};
ram[39974] = {9'd29,-10'd371};
ram[39975] = {9'd32,-10'd368};
ram[39976] = {9'd36,-10'd365};
ram[39977] = {9'd39,-10'd362};
ram[39978] = {9'd42,-10'd359};
ram[39979] = {9'd45,-10'd355};
ram[39980] = {9'd48,-10'd352};
ram[39981] = {9'd51,-10'd349};
ram[39982] = {9'd54,-10'd346};
ram[39983] = {9'd58,-10'd343};
ram[39984] = {9'd61,-10'd340};
ram[39985] = {9'd64,-10'd337};
ram[39986] = {9'd67,-10'd334};
ram[39987] = {9'd70,-10'd330};
ram[39988] = {9'd73,-10'd327};
ram[39989] = {9'd76,-10'd324};
ram[39990] = {9'd80,-10'd321};
ram[39991] = {9'd83,-10'd318};
ram[39992] = {9'd86,-10'd315};
ram[39993] = {9'd89,-10'd312};
ram[39994] = {9'd92,-10'd308};
ram[39995] = {9'd95,-10'd305};
ram[39996] = {9'd98,-10'd302};
ram[39997] = {-9'd99,-10'd299};
ram[39998] = {-9'd96,-10'd296};
ram[39999] = {-9'd92,-10'd293};
ram[40000] = {-9'd89,-10'd290};
ram[40001] = {-9'd86,-10'd286};
ram[40002] = {-9'd83,-10'd283};
ram[40003] = {-9'd80,-10'd280};
ram[40004] = {-9'd77,-10'd277};
ram[40005] = {-9'd74,-10'd274};
ram[40006] = {-9'd70,-10'd271};
ram[40007] = {-9'd67,-10'd268};
ram[40008] = {-9'd64,-10'd264};
ram[40009] = {-9'd61,-10'd261};
ram[40010] = {-9'd58,-10'd258};
ram[40011] = {-9'd55,-10'd255};
ram[40012] = {-9'd52,-10'd252};
ram[40013] = {-9'd48,-10'd249};
ram[40014] = {-9'd45,-10'd246};
ram[40015] = {-9'd42,-10'd242};
ram[40016] = {-9'd39,-10'd239};
ram[40017] = {-9'd36,-10'd236};
ram[40018] = {-9'd33,-10'd233};
ram[40019] = {-9'd30,-10'd230};
ram[40020] = {-9'd26,-10'd227};
ram[40021] = {-9'd23,-10'd224};
ram[40022] = {-9'd20,-10'd220};
ram[40023] = {-9'd17,-10'd217};
ram[40024] = {-9'd14,-10'd214};
ram[40025] = {-9'd11,-10'd211};
ram[40026] = {-9'd8,-10'd208};
ram[40027] = {-9'd4,-10'd205};
ram[40028] = {-9'd1,-10'd202};
ram[40029] = {9'd2,-10'd198};
ram[40030] = {9'd5,-10'd195};
ram[40031] = {9'd8,-10'd192};
ram[40032] = {9'd11,-10'd189};
ram[40033] = {9'd14,-10'd186};
ram[40034] = {9'd18,-10'd183};
ram[40035] = {9'd21,-10'd180};
ram[40036] = {9'd24,-10'd176};
ram[40037] = {9'd27,-10'd173};
ram[40038] = {9'd30,-10'd170};
ram[40039] = {9'd33,-10'd167};
ram[40040] = {9'd36,-10'd164};
ram[40041] = {9'd40,-10'd161};
ram[40042] = {9'd43,-10'd158};
ram[40043] = {9'd46,-10'd154};
ram[40044] = {9'd49,-10'd151};
ram[40045] = {9'd52,-10'd148};
ram[40046] = {9'd55,-10'd145};
ram[40047] = {9'd58,-10'd142};
ram[40048] = {9'd62,-10'd139};
ram[40049] = {9'd65,-10'd136};
ram[40050] = {9'd68,-10'd132};
ram[40051] = {9'd71,-10'd129};
ram[40052] = {9'd74,-10'd126};
ram[40053] = {9'd77,-10'd123};
ram[40054] = {9'd80,-10'd120};
ram[40055] = {9'd84,-10'd117};
ram[40056] = {9'd87,-10'd114};
ram[40057] = {9'd90,-10'd110};
ram[40058] = {9'd93,-10'd107};
ram[40059] = {9'd96,-10'd104};
ram[40060] = {9'd99,-10'd101};
ram[40061] = {-9'd98,-10'd98};
ram[40062] = {-9'd95,-10'd95};
ram[40063] = {-9'd92,-10'd92};
ram[40064] = {-9'd92,-10'd92};
ram[40065] = {-9'd88,-10'd88};
ram[40066] = {-9'd85,-10'd85};
ram[40067] = {-9'd82,-10'd82};
ram[40068] = {-9'd79,-10'd79};
ram[40069] = {-9'd76,-10'd76};
ram[40070] = {-9'd73,-10'd73};
ram[40071] = {-9'd70,-10'd70};
ram[40072] = {-9'd66,-10'd66};
ram[40073] = {-9'd63,-10'd63};
ram[40074] = {-9'd60,-10'd60};
ram[40075] = {-9'd57,-10'd57};
ram[40076] = {-9'd54,-10'd54};
ram[40077] = {-9'd51,-10'd51};
ram[40078] = {-9'd48,-10'd48};
ram[40079] = {-9'd44,-10'd44};
ram[40080] = {-9'd41,-10'd41};
ram[40081] = {-9'd38,-10'd38};
ram[40082] = {-9'd35,-10'd35};
ram[40083] = {-9'd32,-10'd32};
ram[40084] = {-9'd29,-10'd29};
ram[40085] = {-9'd26,-10'd26};
ram[40086] = {-9'd22,-10'd22};
ram[40087] = {-9'd19,-10'd19};
ram[40088] = {-9'd16,-10'd16};
ram[40089] = {-9'd13,-10'd13};
ram[40090] = {-9'd10,-10'd10};
ram[40091] = {-9'd7,-10'd7};
ram[40092] = {-9'd4,-10'd4};
ram[40093] = {9'd0,10'd0};
ram[40094] = {9'd3,10'd3};
ram[40095] = {9'd6,10'd6};
ram[40096] = {9'd9,10'd9};
ram[40097] = {9'd12,10'd12};
ram[40098] = {9'd15,10'd15};
ram[40099] = {9'd18,10'd18};
ram[40100] = {9'd21,10'd21};
ram[40101] = {9'd25,10'd25};
ram[40102] = {9'd28,10'd28};
ram[40103] = {9'd31,10'd31};
ram[40104] = {9'd34,10'd34};
ram[40105] = {9'd37,10'd37};
ram[40106] = {9'd40,10'd40};
ram[40107] = {9'd43,10'd43};
ram[40108] = {9'd47,10'd47};
ram[40109] = {9'd50,10'd50};
ram[40110] = {9'd53,10'd53};
ram[40111] = {9'd56,10'd56};
ram[40112] = {9'd59,10'd59};
ram[40113] = {9'd62,10'd62};
ram[40114] = {9'd65,10'd65};
ram[40115] = {9'd69,10'd69};
ram[40116] = {9'd72,10'd72};
ram[40117] = {9'd75,10'd75};
ram[40118] = {9'd78,10'd78};
ram[40119] = {9'd81,10'd81};
ram[40120] = {9'd84,10'd84};
ram[40121] = {9'd87,10'd87};
ram[40122] = {9'd91,10'd91};
ram[40123] = {9'd94,10'd94};
ram[40124] = {9'd97,10'd97};
ram[40125] = {-9'd100,10'd100};
ram[40126] = {-9'd97,10'd103};
ram[40127] = {-9'd94,10'd106};
ram[40128] = {-9'd91,10'd109};
ram[40129] = {-9'd88,10'd113};
ram[40130] = {-9'd85,10'd116};
ram[40131] = {-9'd81,10'd119};
ram[40132] = {-9'd78,10'd122};
ram[40133] = {-9'd75,10'd125};
ram[40134] = {-9'd72,10'd128};
ram[40135] = {-9'd69,10'd131};
ram[40136] = {-9'd66,10'd135};
ram[40137] = {-9'd63,10'd138};
ram[40138] = {-9'd59,10'd141};
ram[40139] = {-9'd56,10'd144};
ram[40140] = {-9'd53,10'd147};
ram[40141] = {-9'd50,10'd150};
ram[40142] = {-9'd47,10'd153};
ram[40143] = {-9'd44,10'd157};
ram[40144] = {-9'd41,10'd160};
ram[40145] = {-9'd37,10'd163};
ram[40146] = {-9'd34,10'd166};
ram[40147] = {-9'd31,10'd169};
ram[40148] = {-9'd28,10'd172};
ram[40149] = {-9'd25,10'd175};
ram[40150] = {-9'd22,10'd179};
ram[40151] = {-9'd19,10'd182};
ram[40152] = {-9'd15,10'd185};
ram[40153] = {-9'd12,10'd188};
ram[40154] = {-9'd9,10'd191};
ram[40155] = {-9'd6,10'd194};
ram[40156] = {-9'd3,10'd197};
ram[40157] = {9'd0,10'd201};
ram[40158] = {9'd3,10'd204};
ram[40159] = {9'd7,10'd207};
ram[40160] = {9'd10,10'd210};
ram[40161] = {9'd13,10'd213};
ram[40162] = {9'd16,10'd216};
ram[40163] = {9'd19,10'd219};
ram[40164] = {9'd22,10'd223};
ram[40165] = {9'd25,10'd226};
ram[40166] = {9'd29,10'd229};
ram[40167] = {9'd32,10'd232};
ram[40168] = {9'd35,10'd235};
ram[40169] = {9'd38,10'd238};
ram[40170] = {9'd41,10'd241};
ram[40171] = {9'd44,10'd245};
ram[40172] = {9'd47,10'd248};
ram[40173] = {9'd51,10'd251};
ram[40174] = {9'd54,10'd254};
ram[40175] = {9'd57,10'd257};
ram[40176] = {9'd60,10'd260};
ram[40177] = {9'd63,10'd263};
ram[40178] = {9'd66,10'd267};
ram[40179] = {9'd69,10'd270};
ram[40180] = {9'd73,10'd273};
ram[40181] = {9'd76,10'd276};
ram[40182] = {9'd79,10'd279};
ram[40183] = {9'd82,10'd282};
ram[40184] = {9'd85,10'd285};
ram[40185] = {9'd88,10'd289};
ram[40186] = {9'd91,10'd292};
ram[40187] = {9'd95,10'd295};
ram[40188] = {9'd98,10'd298};
ram[40189] = {-9'd99,10'd301};
ram[40190] = {-9'd96,10'd304};
ram[40191] = {-9'd93,10'd307};
ram[40192] = {-9'd93,10'd307};
ram[40193] = {-9'd90,10'd311};
ram[40194] = {-9'd87,10'd314};
ram[40195] = {-9'd84,10'd317};
ram[40196] = {-9'd81,10'd320};
ram[40197] = {-9'd77,10'd323};
ram[40198] = {-9'd74,10'd326};
ram[40199] = {-9'd71,10'd329};
ram[40200] = {-9'd68,10'd333};
ram[40201] = {-9'd65,10'd336};
ram[40202] = {-9'd62,10'd339};
ram[40203] = {-9'd59,10'd342};
ram[40204] = {-9'd55,10'd345};
ram[40205] = {-9'd52,10'd348};
ram[40206] = {-9'd49,10'd351};
ram[40207] = {-9'd46,10'd354};
ram[40208] = {-9'd43,10'd358};
ram[40209] = {-9'd40,10'd361};
ram[40210] = {-9'd37,10'd364};
ram[40211] = {-9'd33,10'd367};
ram[40212] = {-9'd30,10'd370};
ram[40213] = {-9'd27,10'd373};
ram[40214] = {-9'd24,10'd376};
ram[40215] = {-9'd21,10'd380};
ram[40216] = {-9'd18,10'd383};
ram[40217] = {-9'd15,10'd386};
ram[40218] = {-9'd11,10'd389};
ram[40219] = {-9'd8,10'd392};
ram[40220] = {-9'd5,10'd395};
ram[40221] = {-9'd2,10'd398};
ram[40222] = {9'd1,-10'd399};
ram[40223] = {9'd4,-10'd396};
ram[40224] = {9'd7,-10'd393};
ram[40225] = {9'd10,-10'd390};
ram[40226] = {9'd14,-10'd387};
ram[40227] = {9'd17,-10'd384};
ram[40228] = {9'd20,-10'd381};
ram[40229] = {9'd23,-10'd377};
ram[40230] = {9'd26,-10'd374};
ram[40231] = {9'd29,-10'd371};
ram[40232] = {9'd32,-10'd368};
ram[40233] = {9'd36,-10'd365};
ram[40234] = {9'd39,-10'd362};
ram[40235] = {9'd42,-10'd359};
ram[40236] = {9'd45,-10'd355};
ram[40237] = {9'd48,-10'd352};
ram[40238] = {9'd51,-10'd349};
ram[40239] = {9'd54,-10'd346};
ram[40240] = {9'd58,-10'd343};
ram[40241] = {9'd61,-10'd340};
ram[40242] = {9'd64,-10'd337};
ram[40243] = {9'd67,-10'd334};
ram[40244] = {9'd70,-10'd330};
ram[40245] = {9'd73,-10'd327};
ram[40246] = {9'd76,-10'd324};
ram[40247] = {9'd80,-10'd321};
ram[40248] = {9'd83,-10'd318};
ram[40249] = {9'd86,-10'd315};
ram[40250] = {9'd89,-10'd312};
ram[40251] = {9'd92,-10'd308};
ram[40252] = {9'd95,-10'd305};
ram[40253] = {9'd98,-10'd302};
ram[40254] = {-9'd99,-10'd299};
ram[40255] = {-9'd96,-10'd296};
ram[40256] = {-9'd92,-10'd293};
ram[40257] = {-9'd89,-10'd290};
ram[40258] = {-9'd86,-10'd286};
ram[40259] = {-9'd83,-10'd283};
ram[40260] = {-9'd80,-10'd280};
ram[40261] = {-9'd77,-10'd277};
ram[40262] = {-9'd74,-10'd274};
ram[40263] = {-9'd70,-10'd271};
ram[40264] = {-9'd67,-10'd268};
ram[40265] = {-9'd64,-10'd264};
ram[40266] = {-9'd61,-10'd261};
ram[40267] = {-9'd58,-10'd258};
ram[40268] = {-9'd55,-10'd255};
ram[40269] = {-9'd52,-10'd252};
ram[40270] = {-9'd48,-10'd249};
ram[40271] = {-9'd45,-10'd246};
ram[40272] = {-9'd42,-10'd242};
ram[40273] = {-9'd39,-10'd239};
ram[40274] = {-9'd36,-10'd236};
ram[40275] = {-9'd33,-10'd233};
ram[40276] = {-9'd30,-10'd230};
ram[40277] = {-9'd26,-10'd227};
ram[40278] = {-9'd23,-10'd224};
ram[40279] = {-9'd20,-10'd220};
ram[40280] = {-9'd17,-10'd217};
ram[40281] = {-9'd14,-10'd214};
ram[40282] = {-9'd11,-10'd211};
ram[40283] = {-9'd8,-10'd208};
ram[40284] = {-9'd4,-10'd205};
ram[40285] = {-9'd1,-10'd202};
ram[40286] = {9'd2,-10'd198};
ram[40287] = {9'd5,-10'd195};
ram[40288] = {9'd8,-10'd192};
ram[40289] = {9'd11,-10'd189};
ram[40290] = {9'd14,-10'd186};
ram[40291] = {9'd18,-10'd183};
ram[40292] = {9'd21,-10'd180};
ram[40293] = {9'd24,-10'd176};
ram[40294] = {9'd27,-10'd173};
ram[40295] = {9'd30,-10'd170};
ram[40296] = {9'd33,-10'd167};
ram[40297] = {9'd36,-10'd164};
ram[40298] = {9'd40,-10'd161};
ram[40299] = {9'd43,-10'd158};
ram[40300] = {9'd46,-10'd154};
ram[40301] = {9'd49,-10'd151};
ram[40302] = {9'd52,-10'd148};
ram[40303] = {9'd55,-10'd145};
ram[40304] = {9'd58,-10'd142};
ram[40305] = {9'd62,-10'd139};
ram[40306] = {9'd65,-10'd136};
ram[40307] = {9'd68,-10'd132};
ram[40308] = {9'd71,-10'd129};
ram[40309] = {9'd74,-10'd126};
ram[40310] = {9'd77,-10'd123};
ram[40311] = {9'd80,-10'd120};
ram[40312] = {9'd84,-10'd117};
ram[40313] = {9'd87,-10'd114};
ram[40314] = {9'd90,-10'd110};
ram[40315] = {9'd93,-10'd107};
ram[40316] = {9'd96,-10'd104};
ram[40317] = {9'd99,-10'd101};
ram[40318] = {-9'd98,-10'd98};
ram[40319] = {-9'd95,-10'd95};
ram[40320] = {-9'd95,-10'd95};
ram[40321] = {-9'd92,-10'd92};
ram[40322] = {-9'd88,-10'd88};
ram[40323] = {-9'd85,-10'd85};
ram[40324] = {-9'd82,-10'd82};
ram[40325] = {-9'd79,-10'd79};
ram[40326] = {-9'd76,-10'd76};
ram[40327] = {-9'd73,-10'd73};
ram[40328] = {-9'd70,-10'd70};
ram[40329] = {-9'd66,-10'd66};
ram[40330] = {-9'd63,-10'd63};
ram[40331] = {-9'd60,-10'd60};
ram[40332] = {-9'd57,-10'd57};
ram[40333] = {-9'd54,-10'd54};
ram[40334] = {-9'd51,-10'd51};
ram[40335] = {-9'd48,-10'd48};
ram[40336] = {-9'd44,-10'd44};
ram[40337] = {-9'd41,-10'd41};
ram[40338] = {-9'd38,-10'd38};
ram[40339] = {-9'd35,-10'd35};
ram[40340] = {-9'd32,-10'd32};
ram[40341] = {-9'd29,-10'd29};
ram[40342] = {-9'd26,-10'd26};
ram[40343] = {-9'd22,-10'd22};
ram[40344] = {-9'd19,-10'd19};
ram[40345] = {-9'd16,-10'd16};
ram[40346] = {-9'd13,-10'd13};
ram[40347] = {-9'd10,-10'd10};
ram[40348] = {-9'd7,-10'd7};
ram[40349] = {-9'd4,-10'd4};
ram[40350] = {9'd0,10'd0};
ram[40351] = {9'd3,10'd3};
ram[40352] = {9'd6,10'd6};
ram[40353] = {9'd9,10'd9};
ram[40354] = {9'd12,10'd12};
ram[40355] = {9'd15,10'd15};
ram[40356] = {9'd18,10'd18};
ram[40357] = {9'd21,10'd21};
ram[40358] = {9'd25,10'd25};
ram[40359] = {9'd28,10'd28};
ram[40360] = {9'd31,10'd31};
ram[40361] = {9'd34,10'd34};
ram[40362] = {9'd37,10'd37};
ram[40363] = {9'd40,10'd40};
ram[40364] = {9'd43,10'd43};
ram[40365] = {9'd47,10'd47};
ram[40366] = {9'd50,10'd50};
ram[40367] = {9'd53,10'd53};
ram[40368] = {9'd56,10'd56};
ram[40369] = {9'd59,10'd59};
ram[40370] = {9'd62,10'd62};
ram[40371] = {9'd65,10'd65};
ram[40372] = {9'd69,10'd69};
ram[40373] = {9'd72,10'd72};
ram[40374] = {9'd75,10'd75};
ram[40375] = {9'd78,10'd78};
ram[40376] = {9'd81,10'd81};
ram[40377] = {9'd84,10'd84};
ram[40378] = {9'd87,10'd87};
ram[40379] = {9'd91,10'd91};
ram[40380] = {9'd94,10'd94};
ram[40381] = {9'd97,10'd97};
ram[40382] = {-9'd100,10'd100};
ram[40383] = {-9'd97,10'd103};
ram[40384] = {-9'd94,10'd106};
ram[40385] = {-9'd91,10'd109};
ram[40386] = {-9'd88,10'd113};
ram[40387] = {-9'd85,10'd116};
ram[40388] = {-9'd81,10'd119};
ram[40389] = {-9'd78,10'd122};
ram[40390] = {-9'd75,10'd125};
ram[40391] = {-9'd72,10'd128};
ram[40392] = {-9'd69,10'd131};
ram[40393] = {-9'd66,10'd135};
ram[40394] = {-9'd63,10'd138};
ram[40395] = {-9'd59,10'd141};
ram[40396] = {-9'd56,10'd144};
ram[40397] = {-9'd53,10'd147};
ram[40398] = {-9'd50,10'd150};
ram[40399] = {-9'd47,10'd153};
ram[40400] = {-9'd44,10'd157};
ram[40401] = {-9'd41,10'd160};
ram[40402] = {-9'd37,10'd163};
ram[40403] = {-9'd34,10'd166};
ram[40404] = {-9'd31,10'd169};
ram[40405] = {-9'd28,10'd172};
ram[40406] = {-9'd25,10'd175};
ram[40407] = {-9'd22,10'd179};
ram[40408] = {-9'd19,10'd182};
ram[40409] = {-9'd15,10'd185};
ram[40410] = {-9'd12,10'd188};
ram[40411] = {-9'd9,10'd191};
ram[40412] = {-9'd6,10'd194};
ram[40413] = {-9'd3,10'd197};
ram[40414] = {9'd0,10'd201};
ram[40415] = {9'd3,10'd204};
ram[40416] = {9'd7,10'd207};
ram[40417] = {9'd10,10'd210};
ram[40418] = {9'd13,10'd213};
ram[40419] = {9'd16,10'd216};
ram[40420] = {9'd19,10'd219};
ram[40421] = {9'd22,10'd223};
ram[40422] = {9'd25,10'd226};
ram[40423] = {9'd29,10'd229};
ram[40424] = {9'd32,10'd232};
ram[40425] = {9'd35,10'd235};
ram[40426] = {9'd38,10'd238};
ram[40427] = {9'd41,10'd241};
ram[40428] = {9'd44,10'd245};
ram[40429] = {9'd47,10'd248};
ram[40430] = {9'd51,10'd251};
ram[40431] = {9'd54,10'd254};
ram[40432] = {9'd57,10'd257};
ram[40433] = {9'd60,10'd260};
ram[40434] = {9'd63,10'd263};
ram[40435] = {9'd66,10'd267};
ram[40436] = {9'd69,10'd270};
ram[40437] = {9'd73,10'd273};
ram[40438] = {9'd76,10'd276};
ram[40439] = {9'd79,10'd279};
ram[40440] = {9'd82,10'd282};
ram[40441] = {9'd85,10'd285};
ram[40442] = {9'd88,10'd289};
ram[40443] = {9'd91,10'd292};
ram[40444] = {9'd95,10'd295};
ram[40445] = {9'd98,10'd298};
ram[40446] = {-9'd99,10'd301};
ram[40447] = {-9'd96,10'd304};
ram[40448] = {-9'd96,10'd304};
ram[40449] = {-9'd93,10'd307};
ram[40450] = {-9'd90,10'd311};
ram[40451] = {-9'd87,10'd314};
ram[40452] = {-9'd84,10'd317};
ram[40453] = {-9'd81,10'd320};
ram[40454] = {-9'd77,10'd323};
ram[40455] = {-9'd74,10'd326};
ram[40456] = {-9'd71,10'd329};
ram[40457] = {-9'd68,10'd333};
ram[40458] = {-9'd65,10'd336};
ram[40459] = {-9'd62,10'd339};
ram[40460] = {-9'd59,10'd342};
ram[40461] = {-9'd55,10'd345};
ram[40462] = {-9'd52,10'd348};
ram[40463] = {-9'd49,10'd351};
ram[40464] = {-9'd46,10'd354};
ram[40465] = {-9'd43,10'd358};
ram[40466] = {-9'd40,10'd361};
ram[40467] = {-9'd37,10'd364};
ram[40468] = {-9'd33,10'd367};
ram[40469] = {-9'd30,10'd370};
ram[40470] = {-9'd27,10'd373};
ram[40471] = {-9'd24,10'd376};
ram[40472] = {-9'd21,10'd380};
ram[40473] = {-9'd18,10'd383};
ram[40474] = {-9'd15,10'd386};
ram[40475] = {-9'd11,10'd389};
ram[40476] = {-9'd8,10'd392};
ram[40477] = {-9'd5,10'd395};
ram[40478] = {-9'd2,10'd398};
ram[40479] = {9'd1,-10'd399};
ram[40480] = {9'd4,-10'd396};
ram[40481] = {9'd7,-10'd393};
ram[40482] = {9'd10,-10'd390};
ram[40483] = {9'd14,-10'd387};
ram[40484] = {9'd17,-10'd384};
ram[40485] = {9'd20,-10'd381};
ram[40486] = {9'd23,-10'd377};
ram[40487] = {9'd26,-10'd374};
ram[40488] = {9'd29,-10'd371};
ram[40489] = {9'd32,-10'd368};
ram[40490] = {9'd36,-10'd365};
ram[40491] = {9'd39,-10'd362};
ram[40492] = {9'd42,-10'd359};
ram[40493] = {9'd45,-10'd355};
ram[40494] = {9'd48,-10'd352};
ram[40495] = {9'd51,-10'd349};
ram[40496] = {9'd54,-10'd346};
ram[40497] = {9'd58,-10'd343};
ram[40498] = {9'd61,-10'd340};
ram[40499] = {9'd64,-10'd337};
ram[40500] = {9'd67,-10'd334};
ram[40501] = {9'd70,-10'd330};
ram[40502] = {9'd73,-10'd327};
ram[40503] = {9'd76,-10'd324};
ram[40504] = {9'd80,-10'd321};
ram[40505] = {9'd83,-10'd318};
ram[40506] = {9'd86,-10'd315};
ram[40507] = {9'd89,-10'd312};
ram[40508] = {9'd92,-10'd308};
ram[40509] = {9'd95,-10'd305};
ram[40510] = {9'd98,-10'd302};
ram[40511] = {-9'd99,-10'd299};
ram[40512] = {-9'd96,-10'd296};
ram[40513] = {-9'd92,-10'd293};
ram[40514] = {-9'd89,-10'd290};
ram[40515] = {-9'd86,-10'd286};
ram[40516] = {-9'd83,-10'd283};
ram[40517] = {-9'd80,-10'd280};
ram[40518] = {-9'd77,-10'd277};
ram[40519] = {-9'd74,-10'd274};
ram[40520] = {-9'd70,-10'd271};
ram[40521] = {-9'd67,-10'd268};
ram[40522] = {-9'd64,-10'd264};
ram[40523] = {-9'd61,-10'd261};
ram[40524] = {-9'd58,-10'd258};
ram[40525] = {-9'd55,-10'd255};
ram[40526] = {-9'd52,-10'd252};
ram[40527] = {-9'd48,-10'd249};
ram[40528] = {-9'd45,-10'd246};
ram[40529] = {-9'd42,-10'd242};
ram[40530] = {-9'd39,-10'd239};
ram[40531] = {-9'd36,-10'd236};
ram[40532] = {-9'd33,-10'd233};
ram[40533] = {-9'd30,-10'd230};
ram[40534] = {-9'd26,-10'd227};
ram[40535] = {-9'd23,-10'd224};
ram[40536] = {-9'd20,-10'd220};
ram[40537] = {-9'd17,-10'd217};
ram[40538] = {-9'd14,-10'd214};
ram[40539] = {-9'd11,-10'd211};
ram[40540] = {-9'd8,-10'd208};
ram[40541] = {-9'd4,-10'd205};
ram[40542] = {-9'd1,-10'd202};
ram[40543] = {9'd2,-10'd198};
ram[40544] = {9'd5,-10'd195};
ram[40545] = {9'd8,-10'd192};
ram[40546] = {9'd11,-10'd189};
ram[40547] = {9'd14,-10'd186};
ram[40548] = {9'd18,-10'd183};
ram[40549] = {9'd21,-10'd180};
ram[40550] = {9'd24,-10'd176};
ram[40551] = {9'd27,-10'd173};
ram[40552] = {9'd30,-10'd170};
ram[40553] = {9'd33,-10'd167};
ram[40554] = {9'd36,-10'd164};
ram[40555] = {9'd40,-10'd161};
ram[40556] = {9'd43,-10'd158};
ram[40557] = {9'd46,-10'd154};
ram[40558] = {9'd49,-10'd151};
ram[40559] = {9'd52,-10'd148};
ram[40560] = {9'd55,-10'd145};
ram[40561] = {9'd58,-10'd142};
ram[40562] = {9'd62,-10'd139};
ram[40563] = {9'd65,-10'd136};
ram[40564] = {9'd68,-10'd132};
ram[40565] = {9'd71,-10'd129};
ram[40566] = {9'd74,-10'd126};
ram[40567] = {9'd77,-10'd123};
ram[40568] = {9'd80,-10'd120};
ram[40569] = {9'd84,-10'd117};
ram[40570] = {9'd87,-10'd114};
ram[40571] = {9'd90,-10'd110};
ram[40572] = {9'd93,-10'd107};
ram[40573] = {9'd96,-10'd104};
ram[40574] = {9'd99,-10'd101};
ram[40575] = {-9'd98,-10'd98};
ram[40576] = {-9'd98,-10'd98};
ram[40577] = {-9'd95,-10'd95};
ram[40578] = {-9'd92,-10'd92};
ram[40579] = {-9'd88,-10'd88};
ram[40580] = {-9'd85,-10'd85};
ram[40581] = {-9'd82,-10'd82};
ram[40582] = {-9'd79,-10'd79};
ram[40583] = {-9'd76,-10'd76};
ram[40584] = {-9'd73,-10'd73};
ram[40585] = {-9'd70,-10'd70};
ram[40586] = {-9'd66,-10'd66};
ram[40587] = {-9'd63,-10'd63};
ram[40588] = {-9'd60,-10'd60};
ram[40589] = {-9'd57,-10'd57};
ram[40590] = {-9'd54,-10'd54};
ram[40591] = {-9'd51,-10'd51};
ram[40592] = {-9'd48,-10'd48};
ram[40593] = {-9'd44,-10'd44};
ram[40594] = {-9'd41,-10'd41};
ram[40595] = {-9'd38,-10'd38};
ram[40596] = {-9'd35,-10'd35};
ram[40597] = {-9'd32,-10'd32};
ram[40598] = {-9'd29,-10'd29};
ram[40599] = {-9'd26,-10'd26};
ram[40600] = {-9'd22,-10'd22};
ram[40601] = {-9'd19,-10'd19};
ram[40602] = {-9'd16,-10'd16};
ram[40603] = {-9'd13,-10'd13};
ram[40604] = {-9'd10,-10'd10};
ram[40605] = {-9'd7,-10'd7};
ram[40606] = {-9'd4,-10'd4};
ram[40607] = {9'd0,10'd0};
ram[40608] = {9'd3,10'd3};
ram[40609] = {9'd6,10'd6};
ram[40610] = {9'd9,10'd9};
ram[40611] = {9'd12,10'd12};
ram[40612] = {9'd15,10'd15};
ram[40613] = {9'd18,10'd18};
ram[40614] = {9'd21,10'd21};
ram[40615] = {9'd25,10'd25};
ram[40616] = {9'd28,10'd28};
ram[40617] = {9'd31,10'd31};
ram[40618] = {9'd34,10'd34};
ram[40619] = {9'd37,10'd37};
ram[40620] = {9'd40,10'd40};
ram[40621] = {9'd43,10'd43};
ram[40622] = {9'd47,10'd47};
ram[40623] = {9'd50,10'd50};
ram[40624] = {9'd53,10'd53};
ram[40625] = {9'd56,10'd56};
ram[40626] = {9'd59,10'd59};
ram[40627] = {9'd62,10'd62};
ram[40628] = {9'd65,10'd65};
ram[40629] = {9'd69,10'd69};
ram[40630] = {9'd72,10'd72};
ram[40631] = {9'd75,10'd75};
ram[40632] = {9'd78,10'd78};
ram[40633] = {9'd81,10'd81};
ram[40634] = {9'd84,10'd84};
ram[40635] = {9'd87,10'd87};
ram[40636] = {9'd91,10'd91};
ram[40637] = {9'd94,10'd94};
ram[40638] = {9'd97,10'd97};
ram[40639] = {-9'd100,10'd100};
ram[40640] = {-9'd97,10'd103};
ram[40641] = {-9'd94,10'd106};
ram[40642] = {-9'd91,10'd109};
ram[40643] = {-9'd88,10'd113};
ram[40644] = {-9'd85,10'd116};
ram[40645] = {-9'd81,10'd119};
ram[40646] = {-9'd78,10'd122};
ram[40647] = {-9'd75,10'd125};
ram[40648] = {-9'd72,10'd128};
ram[40649] = {-9'd69,10'd131};
ram[40650] = {-9'd66,10'd135};
ram[40651] = {-9'd63,10'd138};
ram[40652] = {-9'd59,10'd141};
ram[40653] = {-9'd56,10'd144};
ram[40654] = {-9'd53,10'd147};
ram[40655] = {-9'd50,10'd150};
ram[40656] = {-9'd47,10'd153};
ram[40657] = {-9'd44,10'd157};
ram[40658] = {-9'd41,10'd160};
ram[40659] = {-9'd37,10'd163};
ram[40660] = {-9'd34,10'd166};
ram[40661] = {-9'd31,10'd169};
ram[40662] = {-9'd28,10'd172};
ram[40663] = {-9'd25,10'd175};
ram[40664] = {-9'd22,10'd179};
ram[40665] = {-9'd19,10'd182};
ram[40666] = {-9'd15,10'd185};
ram[40667] = {-9'd12,10'd188};
ram[40668] = {-9'd9,10'd191};
ram[40669] = {-9'd6,10'd194};
ram[40670] = {-9'd3,10'd197};
ram[40671] = {9'd0,10'd201};
ram[40672] = {9'd3,10'd204};
ram[40673] = {9'd7,10'd207};
ram[40674] = {9'd10,10'd210};
ram[40675] = {9'd13,10'd213};
ram[40676] = {9'd16,10'd216};
ram[40677] = {9'd19,10'd219};
ram[40678] = {9'd22,10'd223};
ram[40679] = {9'd25,10'd226};
ram[40680] = {9'd29,10'd229};
ram[40681] = {9'd32,10'd232};
ram[40682] = {9'd35,10'd235};
ram[40683] = {9'd38,10'd238};
ram[40684] = {9'd41,10'd241};
ram[40685] = {9'd44,10'd245};
ram[40686] = {9'd47,10'd248};
ram[40687] = {9'd51,10'd251};
ram[40688] = {9'd54,10'd254};
ram[40689] = {9'd57,10'd257};
ram[40690] = {9'd60,10'd260};
ram[40691] = {9'd63,10'd263};
ram[40692] = {9'd66,10'd267};
ram[40693] = {9'd69,10'd270};
ram[40694] = {9'd73,10'd273};
ram[40695] = {9'd76,10'd276};
ram[40696] = {9'd79,10'd279};
ram[40697] = {9'd82,10'd282};
ram[40698] = {9'd85,10'd285};
ram[40699] = {9'd88,10'd289};
ram[40700] = {9'd91,10'd292};
ram[40701] = {9'd95,10'd295};
ram[40702] = {9'd98,10'd298};
ram[40703] = {-9'd99,10'd301};
ram[40704] = {-9'd99,10'd301};
ram[40705] = {-9'd96,10'd304};
ram[40706] = {-9'd93,10'd307};
ram[40707] = {-9'd90,10'd311};
ram[40708] = {-9'd87,10'd314};
ram[40709] = {-9'd84,10'd317};
ram[40710] = {-9'd81,10'd320};
ram[40711] = {-9'd77,10'd323};
ram[40712] = {-9'd74,10'd326};
ram[40713] = {-9'd71,10'd329};
ram[40714] = {-9'd68,10'd333};
ram[40715] = {-9'd65,10'd336};
ram[40716] = {-9'd62,10'd339};
ram[40717] = {-9'd59,10'd342};
ram[40718] = {-9'd55,10'd345};
ram[40719] = {-9'd52,10'd348};
ram[40720] = {-9'd49,10'd351};
ram[40721] = {-9'd46,10'd354};
ram[40722] = {-9'd43,10'd358};
ram[40723] = {-9'd40,10'd361};
ram[40724] = {-9'd37,10'd364};
ram[40725] = {-9'd33,10'd367};
ram[40726] = {-9'd30,10'd370};
ram[40727] = {-9'd27,10'd373};
ram[40728] = {-9'd24,10'd376};
ram[40729] = {-9'd21,10'd380};
ram[40730] = {-9'd18,10'd383};
ram[40731] = {-9'd15,10'd386};
ram[40732] = {-9'd11,10'd389};
ram[40733] = {-9'd8,10'd392};
ram[40734] = {-9'd5,10'd395};
ram[40735] = {-9'd2,10'd398};
ram[40736] = {9'd1,-10'd399};
ram[40737] = {9'd4,-10'd396};
ram[40738] = {9'd7,-10'd393};
ram[40739] = {9'd10,-10'd390};
ram[40740] = {9'd14,-10'd387};
ram[40741] = {9'd17,-10'd384};
ram[40742] = {9'd20,-10'd381};
ram[40743] = {9'd23,-10'd377};
ram[40744] = {9'd26,-10'd374};
ram[40745] = {9'd29,-10'd371};
ram[40746] = {9'd32,-10'd368};
ram[40747] = {9'd36,-10'd365};
ram[40748] = {9'd39,-10'd362};
ram[40749] = {9'd42,-10'd359};
ram[40750] = {9'd45,-10'd355};
ram[40751] = {9'd48,-10'd352};
ram[40752] = {9'd51,-10'd349};
ram[40753] = {9'd54,-10'd346};
ram[40754] = {9'd58,-10'd343};
ram[40755] = {9'd61,-10'd340};
ram[40756] = {9'd64,-10'd337};
ram[40757] = {9'd67,-10'd334};
ram[40758] = {9'd70,-10'd330};
ram[40759] = {9'd73,-10'd327};
ram[40760] = {9'd76,-10'd324};
ram[40761] = {9'd80,-10'd321};
ram[40762] = {9'd83,-10'd318};
ram[40763] = {9'd86,-10'd315};
ram[40764] = {9'd89,-10'd312};
ram[40765] = {9'd92,-10'd308};
ram[40766] = {9'd95,-10'd305};
ram[40767] = {9'd98,-10'd302};
ram[40768] = {-9'd99,-10'd299};
ram[40769] = {-9'd96,-10'd296};
ram[40770] = {-9'd92,-10'd293};
ram[40771] = {-9'd89,-10'd290};
ram[40772] = {-9'd86,-10'd286};
ram[40773] = {-9'd83,-10'd283};
ram[40774] = {-9'd80,-10'd280};
ram[40775] = {-9'd77,-10'd277};
ram[40776] = {-9'd74,-10'd274};
ram[40777] = {-9'd70,-10'd271};
ram[40778] = {-9'd67,-10'd268};
ram[40779] = {-9'd64,-10'd264};
ram[40780] = {-9'd61,-10'd261};
ram[40781] = {-9'd58,-10'd258};
ram[40782] = {-9'd55,-10'd255};
ram[40783] = {-9'd52,-10'd252};
ram[40784] = {-9'd48,-10'd249};
ram[40785] = {-9'd45,-10'd246};
ram[40786] = {-9'd42,-10'd242};
ram[40787] = {-9'd39,-10'd239};
ram[40788] = {-9'd36,-10'd236};
ram[40789] = {-9'd33,-10'd233};
ram[40790] = {-9'd30,-10'd230};
ram[40791] = {-9'd26,-10'd227};
ram[40792] = {-9'd23,-10'd224};
ram[40793] = {-9'd20,-10'd220};
ram[40794] = {-9'd17,-10'd217};
ram[40795] = {-9'd14,-10'd214};
ram[40796] = {-9'd11,-10'd211};
ram[40797] = {-9'd8,-10'd208};
ram[40798] = {-9'd4,-10'd205};
ram[40799] = {-9'd1,-10'd202};
ram[40800] = {9'd2,-10'd198};
ram[40801] = {9'd5,-10'd195};
ram[40802] = {9'd8,-10'd192};
ram[40803] = {9'd11,-10'd189};
ram[40804] = {9'd14,-10'd186};
ram[40805] = {9'd18,-10'd183};
ram[40806] = {9'd21,-10'd180};
ram[40807] = {9'd24,-10'd176};
ram[40808] = {9'd27,-10'd173};
ram[40809] = {9'd30,-10'd170};
ram[40810] = {9'd33,-10'd167};
ram[40811] = {9'd36,-10'd164};
ram[40812] = {9'd40,-10'd161};
ram[40813] = {9'd43,-10'd158};
ram[40814] = {9'd46,-10'd154};
ram[40815] = {9'd49,-10'd151};
ram[40816] = {9'd52,-10'd148};
ram[40817] = {9'd55,-10'd145};
ram[40818] = {9'd58,-10'd142};
ram[40819] = {9'd62,-10'd139};
ram[40820] = {9'd65,-10'd136};
ram[40821] = {9'd68,-10'd132};
ram[40822] = {9'd71,-10'd129};
ram[40823] = {9'd74,-10'd126};
ram[40824] = {9'd77,-10'd123};
ram[40825] = {9'd80,-10'd120};
ram[40826] = {9'd84,-10'd117};
ram[40827] = {9'd87,-10'd114};
ram[40828] = {9'd90,-10'd110};
ram[40829] = {9'd93,-10'd107};
ram[40830] = {9'd96,-10'd104};
ram[40831] = {9'd99,-10'd101};
ram[40832] = {9'd99,-10'd101};
ram[40833] = {-9'd98,-10'd98};
ram[40834] = {-9'd95,-10'd95};
ram[40835] = {-9'd92,-10'd92};
ram[40836] = {-9'd88,-10'd88};
ram[40837] = {-9'd85,-10'd85};
ram[40838] = {-9'd82,-10'd82};
ram[40839] = {-9'd79,-10'd79};
ram[40840] = {-9'd76,-10'd76};
ram[40841] = {-9'd73,-10'd73};
ram[40842] = {-9'd70,-10'd70};
ram[40843] = {-9'd66,-10'd66};
ram[40844] = {-9'd63,-10'd63};
ram[40845] = {-9'd60,-10'd60};
ram[40846] = {-9'd57,-10'd57};
ram[40847] = {-9'd54,-10'd54};
ram[40848] = {-9'd51,-10'd51};
ram[40849] = {-9'd48,-10'd48};
ram[40850] = {-9'd44,-10'd44};
ram[40851] = {-9'd41,-10'd41};
ram[40852] = {-9'd38,-10'd38};
ram[40853] = {-9'd35,-10'd35};
ram[40854] = {-9'd32,-10'd32};
ram[40855] = {-9'd29,-10'd29};
ram[40856] = {-9'd26,-10'd26};
ram[40857] = {-9'd22,-10'd22};
ram[40858] = {-9'd19,-10'd19};
ram[40859] = {-9'd16,-10'd16};
ram[40860] = {-9'd13,-10'd13};
ram[40861] = {-9'd10,-10'd10};
ram[40862] = {-9'd7,-10'd7};
ram[40863] = {-9'd4,-10'd4};
ram[40864] = {9'd0,10'd0};
ram[40865] = {9'd3,10'd3};
ram[40866] = {9'd6,10'd6};
ram[40867] = {9'd9,10'd9};
ram[40868] = {9'd12,10'd12};
ram[40869] = {9'd15,10'd15};
ram[40870] = {9'd18,10'd18};
ram[40871] = {9'd21,10'd21};
ram[40872] = {9'd25,10'd25};
ram[40873] = {9'd28,10'd28};
ram[40874] = {9'd31,10'd31};
ram[40875] = {9'd34,10'd34};
ram[40876] = {9'd37,10'd37};
ram[40877] = {9'd40,10'd40};
ram[40878] = {9'd43,10'd43};
ram[40879] = {9'd47,10'd47};
ram[40880] = {9'd50,10'd50};
ram[40881] = {9'd53,10'd53};
ram[40882] = {9'd56,10'd56};
ram[40883] = {9'd59,10'd59};
ram[40884] = {9'd62,10'd62};
ram[40885] = {9'd65,10'd65};
ram[40886] = {9'd69,10'd69};
ram[40887] = {9'd72,10'd72};
ram[40888] = {9'd75,10'd75};
ram[40889] = {9'd78,10'd78};
ram[40890] = {9'd81,10'd81};
ram[40891] = {9'd84,10'd84};
ram[40892] = {9'd87,10'd87};
ram[40893] = {9'd91,10'd91};
ram[40894] = {9'd94,10'd94};
ram[40895] = {9'd97,10'd97};
ram[40896] = {-9'd100,10'd100};
ram[40897] = {-9'd97,10'd103};
ram[40898] = {-9'd94,10'd106};
ram[40899] = {-9'd91,10'd109};
ram[40900] = {-9'd88,10'd113};
ram[40901] = {-9'd85,10'd116};
ram[40902] = {-9'd81,10'd119};
ram[40903] = {-9'd78,10'd122};
ram[40904] = {-9'd75,10'd125};
ram[40905] = {-9'd72,10'd128};
ram[40906] = {-9'd69,10'd131};
ram[40907] = {-9'd66,10'd135};
ram[40908] = {-9'd63,10'd138};
ram[40909] = {-9'd59,10'd141};
ram[40910] = {-9'd56,10'd144};
ram[40911] = {-9'd53,10'd147};
ram[40912] = {-9'd50,10'd150};
ram[40913] = {-9'd47,10'd153};
ram[40914] = {-9'd44,10'd157};
ram[40915] = {-9'd41,10'd160};
ram[40916] = {-9'd37,10'd163};
ram[40917] = {-9'd34,10'd166};
ram[40918] = {-9'd31,10'd169};
ram[40919] = {-9'd28,10'd172};
ram[40920] = {-9'd25,10'd175};
ram[40921] = {-9'd22,10'd179};
ram[40922] = {-9'd19,10'd182};
ram[40923] = {-9'd15,10'd185};
ram[40924] = {-9'd12,10'd188};
ram[40925] = {-9'd9,10'd191};
ram[40926] = {-9'd6,10'd194};
ram[40927] = {-9'd3,10'd197};
ram[40928] = {9'd0,10'd201};
ram[40929] = {9'd3,10'd204};
ram[40930] = {9'd7,10'd207};
ram[40931] = {9'd10,10'd210};
ram[40932] = {9'd13,10'd213};
ram[40933] = {9'd16,10'd216};
ram[40934] = {9'd19,10'd219};
ram[40935] = {9'd22,10'd223};
ram[40936] = {9'd25,10'd226};
ram[40937] = {9'd29,10'd229};
ram[40938] = {9'd32,10'd232};
ram[40939] = {9'd35,10'd235};
ram[40940] = {9'd38,10'd238};
ram[40941] = {9'd41,10'd241};
ram[40942] = {9'd44,10'd245};
ram[40943] = {9'd47,10'd248};
ram[40944] = {9'd51,10'd251};
ram[40945] = {9'd54,10'd254};
ram[40946] = {9'd57,10'd257};
ram[40947] = {9'd60,10'd260};
ram[40948] = {9'd63,10'd263};
ram[40949] = {9'd66,10'd267};
ram[40950] = {9'd69,10'd270};
ram[40951] = {9'd73,10'd273};
ram[40952] = {9'd76,10'd276};
ram[40953] = {9'd79,10'd279};
ram[40954] = {9'd82,10'd282};
ram[40955] = {9'd85,10'd285};
ram[40956] = {9'd88,10'd289};
ram[40957] = {9'd91,10'd292};
ram[40958] = {9'd95,10'd295};
ram[40959] = {9'd98,10'd298};
ram[40960] = {9'd98,10'd298};
ram[40961] = {-9'd99,10'd301};
ram[40962] = {-9'd96,10'd304};
ram[40963] = {-9'd93,10'd307};
ram[40964] = {-9'd90,10'd311};
ram[40965] = {-9'd87,10'd314};
ram[40966] = {-9'd84,10'd317};
ram[40967] = {-9'd81,10'd320};
ram[40968] = {-9'd77,10'd323};
ram[40969] = {-9'd74,10'd326};
ram[40970] = {-9'd71,10'd329};
ram[40971] = {-9'd68,10'd333};
ram[40972] = {-9'd65,10'd336};
ram[40973] = {-9'd62,10'd339};
ram[40974] = {-9'd59,10'd342};
ram[40975] = {-9'd55,10'd345};
ram[40976] = {-9'd52,10'd348};
ram[40977] = {-9'd49,10'd351};
ram[40978] = {-9'd46,10'd354};
ram[40979] = {-9'd43,10'd358};
ram[40980] = {-9'd40,10'd361};
ram[40981] = {-9'd37,10'd364};
ram[40982] = {-9'd33,10'd367};
ram[40983] = {-9'd30,10'd370};
ram[40984] = {-9'd27,10'd373};
ram[40985] = {-9'd24,10'd376};
ram[40986] = {-9'd21,10'd380};
ram[40987] = {-9'd18,10'd383};
ram[40988] = {-9'd15,10'd386};
ram[40989] = {-9'd11,10'd389};
ram[40990] = {-9'd8,10'd392};
ram[40991] = {-9'd5,10'd395};
ram[40992] = {-9'd2,10'd398};
ram[40993] = {9'd1,-10'd399};
ram[40994] = {9'd4,-10'd396};
ram[40995] = {9'd7,-10'd393};
ram[40996] = {9'd10,-10'd390};
ram[40997] = {9'd14,-10'd387};
ram[40998] = {9'd17,-10'd384};
ram[40999] = {9'd20,-10'd381};
ram[41000] = {9'd23,-10'd377};
ram[41001] = {9'd26,-10'd374};
ram[41002] = {9'd29,-10'd371};
ram[41003] = {9'd32,-10'd368};
ram[41004] = {9'd36,-10'd365};
ram[41005] = {9'd39,-10'd362};
ram[41006] = {9'd42,-10'd359};
ram[41007] = {9'd45,-10'd355};
ram[41008] = {9'd48,-10'd352};
ram[41009] = {9'd51,-10'd349};
ram[41010] = {9'd54,-10'd346};
ram[41011] = {9'd58,-10'd343};
ram[41012] = {9'd61,-10'd340};
ram[41013] = {9'd64,-10'd337};
ram[41014] = {9'd67,-10'd334};
ram[41015] = {9'd70,-10'd330};
ram[41016] = {9'd73,-10'd327};
ram[41017] = {9'd76,-10'd324};
ram[41018] = {9'd80,-10'd321};
ram[41019] = {9'd83,-10'd318};
ram[41020] = {9'd86,-10'd315};
ram[41021] = {9'd89,-10'd312};
ram[41022] = {9'd92,-10'd308};
ram[41023] = {9'd95,-10'd305};
ram[41024] = {9'd98,-10'd302};
ram[41025] = {-9'd99,-10'd299};
ram[41026] = {-9'd96,-10'd296};
ram[41027] = {-9'd92,-10'd293};
ram[41028] = {-9'd89,-10'd290};
ram[41029] = {-9'd86,-10'd286};
ram[41030] = {-9'd83,-10'd283};
ram[41031] = {-9'd80,-10'd280};
ram[41032] = {-9'd77,-10'd277};
ram[41033] = {-9'd74,-10'd274};
ram[41034] = {-9'd70,-10'd271};
ram[41035] = {-9'd67,-10'd268};
ram[41036] = {-9'd64,-10'd264};
ram[41037] = {-9'd61,-10'd261};
ram[41038] = {-9'd58,-10'd258};
ram[41039] = {-9'd55,-10'd255};
ram[41040] = {-9'd52,-10'd252};
ram[41041] = {-9'd48,-10'd249};
ram[41042] = {-9'd45,-10'd246};
ram[41043] = {-9'd42,-10'd242};
ram[41044] = {-9'd39,-10'd239};
ram[41045] = {-9'd36,-10'd236};
ram[41046] = {-9'd33,-10'd233};
ram[41047] = {-9'd30,-10'd230};
ram[41048] = {-9'd26,-10'd227};
ram[41049] = {-9'd23,-10'd224};
ram[41050] = {-9'd20,-10'd220};
ram[41051] = {-9'd17,-10'd217};
ram[41052] = {-9'd14,-10'd214};
ram[41053] = {-9'd11,-10'd211};
ram[41054] = {-9'd8,-10'd208};
ram[41055] = {-9'd4,-10'd205};
ram[41056] = {-9'd1,-10'd202};
ram[41057] = {9'd2,-10'd198};
ram[41058] = {9'd5,-10'd195};
ram[41059] = {9'd8,-10'd192};
ram[41060] = {9'd11,-10'd189};
ram[41061] = {9'd14,-10'd186};
ram[41062] = {9'd18,-10'd183};
ram[41063] = {9'd21,-10'd180};
ram[41064] = {9'd24,-10'd176};
ram[41065] = {9'd27,-10'd173};
ram[41066] = {9'd30,-10'd170};
ram[41067] = {9'd33,-10'd167};
ram[41068] = {9'd36,-10'd164};
ram[41069] = {9'd40,-10'd161};
ram[41070] = {9'd43,-10'd158};
ram[41071] = {9'd46,-10'd154};
ram[41072] = {9'd49,-10'd151};
ram[41073] = {9'd52,-10'd148};
ram[41074] = {9'd55,-10'd145};
ram[41075] = {9'd58,-10'd142};
ram[41076] = {9'd62,-10'd139};
ram[41077] = {9'd65,-10'd136};
ram[41078] = {9'd68,-10'd132};
ram[41079] = {9'd71,-10'd129};
ram[41080] = {9'd74,-10'd126};
ram[41081] = {9'd77,-10'd123};
ram[41082] = {9'd80,-10'd120};
ram[41083] = {9'd84,-10'd117};
ram[41084] = {9'd87,-10'd114};
ram[41085] = {9'd90,-10'd110};
ram[41086] = {9'd93,-10'd107};
ram[41087] = {9'd96,-10'd104};
ram[41088] = {9'd96,-10'd104};
ram[41089] = {9'd99,-10'd101};
ram[41090] = {-9'd98,-10'd98};
ram[41091] = {-9'd95,-10'd95};
ram[41092] = {-9'd92,-10'd92};
ram[41093] = {-9'd88,-10'd88};
ram[41094] = {-9'd85,-10'd85};
ram[41095] = {-9'd82,-10'd82};
ram[41096] = {-9'd79,-10'd79};
ram[41097] = {-9'd76,-10'd76};
ram[41098] = {-9'd73,-10'd73};
ram[41099] = {-9'd70,-10'd70};
ram[41100] = {-9'd66,-10'd66};
ram[41101] = {-9'd63,-10'd63};
ram[41102] = {-9'd60,-10'd60};
ram[41103] = {-9'd57,-10'd57};
ram[41104] = {-9'd54,-10'd54};
ram[41105] = {-9'd51,-10'd51};
ram[41106] = {-9'd48,-10'd48};
ram[41107] = {-9'd44,-10'd44};
ram[41108] = {-9'd41,-10'd41};
ram[41109] = {-9'd38,-10'd38};
ram[41110] = {-9'd35,-10'd35};
ram[41111] = {-9'd32,-10'd32};
ram[41112] = {-9'd29,-10'd29};
ram[41113] = {-9'd26,-10'd26};
ram[41114] = {-9'd22,-10'd22};
ram[41115] = {-9'd19,-10'd19};
ram[41116] = {-9'd16,-10'd16};
ram[41117] = {-9'd13,-10'd13};
ram[41118] = {-9'd10,-10'd10};
ram[41119] = {-9'd7,-10'd7};
ram[41120] = {-9'd4,-10'd4};
ram[41121] = {9'd0,10'd0};
ram[41122] = {9'd3,10'd3};
ram[41123] = {9'd6,10'd6};
ram[41124] = {9'd9,10'd9};
ram[41125] = {9'd12,10'd12};
ram[41126] = {9'd15,10'd15};
ram[41127] = {9'd18,10'd18};
ram[41128] = {9'd21,10'd21};
ram[41129] = {9'd25,10'd25};
ram[41130] = {9'd28,10'd28};
ram[41131] = {9'd31,10'd31};
ram[41132] = {9'd34,10'd34};
ram[41133] = {9'd37,10'd37};
ram[41134] = {9'd40,10'd40};
ram[41135] = {9'd43,10'd43};
ram[41136] = {9'd47,10'd47};
ram[41137] = {9'd50,10'd50};
ram[41138] = {9'd53,10'd53};
ram[41139] = {9'd56,10'd56};
ram[41140] = {9'd59,10'd59};
ram[41141] = {9'd62,10'd62};
ram[41142] = {9'd65,10'd65};
ram[41143] = {9'd69,10'd69};
ram[41144] = {9'd72,10'd72};
ram[41145] = {9'd75,10'd75};
ram[41146] = {9'd78,10'd78};
ram[41147] = {9'd81,10'd81};
ram[41148] = {9'd84,10'd84};
ram[41149] = {9'd87,10'd87};
ram[41150] = {9'd91,10'd91};
ram[41151] = {9'd94,10'd94};
ram[41152] = {9'd97,10'd97};
ram[41153] = {-9'd100,10'd100};
ram[41154] = {-9'd97,10'd103};
ram[41155] = {-9'd94,10'd106};
ram[41156] = {-9'd91,10'd109};
ram[41157] = {-9'd88,10'd113};
ram[41158] = {-9'd85,10'd116};
ram[41159] = {-9'd81,10'd119};
ram[41160] = {-9'd78,10'd122};
ram[41161] = {-9'd75,10'd125};
ram[41162] = {-9'd72,10'd128};
ram[41163] = {-9'd69,10'd131};
ram[41164] = {-9'd66,10'd135};
ram[41165] = {-9'd63,10'd138};
ram[41166] = {-9'd59,10'd141};
ram[41167] = {-9'd56,10'd144};
ram[41168] = {-9'd53,10'd147};
ram[41169] = {-9'd50,10'd150};
ram[41170] = {-9'd47,10'd153};
ram[41171] = {-9'd44,10'd157};
ram[41172] = {-9'd41,10'd160};
ram[41173] = {-9'd37,10'd163};
ram[41174] = {-9'd34,10'd166};
ram[41175] = {-9'd31,10'd169};
ram[41176] = {-9'd28,10'd172};
ram[41177] = {-9'd25,10'd175};
ram[41178] = {-9'd22,10'd179};
ram[41179] = {-9'd19,10'd182};
ram[41180] = {-9'd15,10'd185};
ram[41181] = {-9'd12,10'd188};
ram[41182] = {-9'd9,10'd191};
ram[41183] = {-9'd6,10'd194};
ram[41184] = {-9'd3,10'd197};
ram[41185] = {9'd0,10'd201};
ram[41186] = {9'd3,10'd204};
ram[41187] = {9'd7,10'd207};
ram[41188] = {9'd10,10'd210};
ram[41189] = {9'd13,10'd213};
ram[41190] = {9'd16,10'd216};
ram[41191] = {9'd19,10'd219};
ram[41192] = {9'd22,10'd223};
ram[41193] = {9'd25,10'd226};
ram[41194] = {9'd29,10'd229};
ram[41195] = {9'd32,10'd232};
ram[41196] = {9'd35,10'd235};
ram[41197] = {9'd38,10'd238};
ram[41198] = {9'd41,10'd241};
ram[41199] = {9'd44,10'd245};
ram[41200] = {9'd47,10'd248};
ram[41201] = {9'd51,10'd251};
ram[41202] = {9'd54,10'd254};
ram[41203] = {9'd57,10'd257};
ram[41204] = {9'd60,10'd260};
ram[41205] = {9'd63,10'd263};
ram[41206] = {9'd66,10'd267};
ram[41207] = {9'd69,10'd270};
ram[41208] = {9'd73,10'd273};
ram[41209] = {9'd76,10'd276};
ram[41210] = {9'd79,10'd279};
ram[41211] = {9'd82,10'd282};
ram[41212] = {9'd85,10'd285};
ram[41213] = {9'd88,10'd289};
ram[41214] = {9'd91,10'd292};
ram[41215] = {9'd95,10'd295};
ram[41216] = {9'd95,10'd295};
ram[41217] = {9'd98,10'd298};
ram[41218] = {-9'd99,10'd301};
ram[41219] = {-9'd96,10'd304};
ram[41220] = {-9'd93,10'd307};
ram[41221] = {-9'd90,10'd311};
ram[41222] = {-9'd87,10'd314};
ram[41223] = {-9'd84,10'd317};
ram[41224] = {-9'd81,10'd320};
ram[41225] = {-9'd77,10'd323};
ram[41226] = {-9'd74,10'd326};
ram[41227] = {-9'd71,10'd329};
ram[41228] = {-9'd68,10'd333};
ram[41229] = {-9'd65,10'd336};
ram[41230] = {-9'd62,10'd339};
ram[41231] = {-9'd59,10'd342};
ram[41232] = {-9'd55,10'd345};
ram[41233] = {-9'd52,10'd348};
ram[41234] = {-9'd49,10'd351};
ram[41235] = {-9'd46,10'd354};
ram[41236] = {-9'd43,10'd358};
ram[41237] = {-9'd40,10'd361};
ram[41238] = {-9'd37,10'd364};
ram[41239] = {-9'd33,10'd367};
ram[41240] = {-9'd30,10'd370};
ram[41241] = {-9'd27,10'd373};
ram[41242] = {-9'd24,10'd376};
ram[41243] = {-9'd21,10'd380};
ram[41244] = {-9'd18,10'd383};
ram[41245] = {-9'd15,10'd386};
ram[41246] = {-9'd11,10'd389};
ram[41247] = {-9'd8,10'd392};
ram[41248] = {-9'd5,10'd395};
ram[41249] = {-9'd2,10'd398};
ram[41250] = {9'd1,-10'd399};
ram[41251] = {9'd4,-10'd396};
ram[41252] = {9'd7,-10'd393};
ram[41253] = {9'd10,-10'd390};
ram[41254] = {9'd14,-10'd387};
ram[41255] = {9'd17,-10'd384};
ram[41256] = {9'd20,-10'd381};
ram[41257] = {9'd23,-10'd377};
ram[41258] = {9'd26,-10'd374};
ram[41259] = {9'd29,-10'd371};
ram[41260] = {9'd32,-10'd368};
ram[41261] = {9'd36,-10'd365};
ram[41262] = {9'd39,-10'd362};
ram[41263] = {9'd42,-10'd359};
ram[41264] = {9'd45,-10'd355};
ram[41265] = {9'd48,-10'd352};
ram[41266] = {9'd51,-10'd349};
ram[41267] = {9'd54,-10'd346};
ram[41268] = {9'd58,-10'd343};
ram[41269] = {9'd61,-10'd340};
ram[41270] = {9'd64,-10'd337};
ram[41271] = {9'd67,-10'd334};
ram[41272] = {9'd70,-10'd330};
ram[41273] = {9'd73,-10'd327};
ram[41274] = {9'd76,-10'd324};
ram[41275] = {9'd80,-10'd321};
ram[41276] = {9'd83,-10'd318};
ram[41277] = {9'd86,-10'd315};
ram[41278] = {9'd89,-10'd312};
ram[41279] = {9'd92,-10'd308};
ram[41280] = {9'd95,-10'd305};
ram[41281] = {9'd98,-10'd302};
ram[41282] = {-9'd99,-10'd299};
ram[41283] = {-9'd96,-10'd296};
ram[41284] = {-9'd92,-10'd293};
ram[41285] = {-9'd89,-10'd290};
ram[41286] = {-9'd86,-10'd286};
ram[41287] = {-9'd83,-10'd283};
ram[41288] = {-9'd80,-10'd280};
ram[41289] = {-9'd77,-10'd277};
ram[41290] = {-9'd74,-10'd274};
ram[41291] = {-9'd70,-10'd271};
ram[41292] = {-9'd67,-10'd268};
ram[41293] = {-9'd64,-10'd264};
ram[41294] = {-9'd61,-10'd261};
ram[41295] = {-9'd58,-10'd258};
ram[41296] = {-9'd55,-10'd255};
ram[41297] = {-9'd52,-10'd252};
ram[41298] = {-9'd48,-10'd249};
ram[41299] = {-9'd45,-10'd246};
ram[41300] = {-9'd42,-10'd242};
ram[41301] = {-9'd39,-10'd239};
ram[41302] = {-9'd36,-10'd236};
ram[41303] = {-9'd33,-10'd233};
ram[41304] = {-9'd30,-10'd230};
ram[41305] = {-9'd26,-10'd227};
ram[41306] = {-9'd23,-10'd224};
ram[41307] = {-9'd20,-10'd220};
ram[41308] = {-9'd17,-10'd217};
ram[41309] = {-9'd14,-10'd214};
ram[41310] = {-9'd11,-10'd211};
ram[41311] = {-9'd8,-10'd208};
ram[41312] = {-9'd4,-10'd205};
ram[41313] = {-9'd1,-10'd202};
ram[41314] = {9'd2,-10'd198};
ram[41315] = {9'd5,-10'd195};
ram[41316] = {9'd8,-10'd192};
ram[41317] = {9'd11,-10'd189};
ram[41318] = {9'd14,-10'd186};
ram[41319] = {9'd18,-10'd183};
ram[41320] = {9'd21,-10'd180};
ram[41321] = {9'd24,-10'd176};
ram[41322] = {9'd27,-10'd173};
ram[41323] = {9'd30,-10'd170};
ram[41324] = {9'd33,-10'd167};
ram[41325] = {9'd36,-10'd164};
ram[41326] = {9'd40,-10'd161};
ram[41327] = {9'd43,-10'd158};
ram[41328] = {9'd46,-10'd154};
ram[41329] = {9'd49,-10'd151};
ram[41330] = {9'd52,-10'd148};
ram[41331] = {9'd55,-10'd145};
ram[41332] = {9'd58,-10'd142};
ram[41333] = {9'd62,-10'd139};
ram[41334] = {9'd65,-10'd136};
ram[41335] = {9'd68,-10'd132};
ram[41336] = {9'd71,-10'd129};
ram[41337] = {9'd74,-10'd126};
ram[41338] = {9'd77,-10'd123};
ram[41339] = {9'd80,-10'd120};
ram[41340] = {9'd84,-10'd117};
ram[41341] = {9'd87,-10'd114};
ram[41342] = {9'd90,-10'd110};
ram[41343] = {9'd93,-10'd107};
ram[41344] = {9'd93,-10'd107};
ram[41345] = {9'd96,-10'd104};
ram[41346] = {9'd99,-10'd101};
ram[41347] = {-9'd98,-10'd98};
ram[41348] = {-9'd95,-10'd95};
ram[41349] = {-9'd92,-10'd92};
ram[41350] = {-9'd88,-10'd88};
ram[41351] = {-9'd85,-10'd85};
ram[41352] = {-9'd82,-10'd82};
ram[41353] = {-9'd79,-10'd79};
ram[41354] = {-9'd76,-10'd76};
ram[41355] = {-9'd73,-10'd73};
ram[41356] = {-9'd70,-10'd70};
ram[41357] = {-9'd66,-10'd66};
ram[41358] = {-9'd63,-10'd63};
ram[41359] = {-9'd60,-10'd60};
ram[41360] = {-9'd57,-10'd57};
ram[41361] = {-9'd54,-10'd54};
ram[41362] = {-9'd51,-10'd51};
ram[41363] = {-9'd48,-10'd48};
ram[41364] = {-9'd44,-10'd44};
ram[41365] = {-9'd41,-10'd41};
ram[41366] = {-9'd38,-10'd38};
ram[41367] = {-9'd35,-10'd35};
ram[41368] = {-9'd32,-10'd32};
ram[41369] = {-9'd29,-10'd29};
ram[41370] = {-9'd26,-10'd26};
ram[41371] = {-9'd22,-10'd22};
ram[41372] = {-9'd19,-10'd19};
ram[41373] = {-9'd16,-10'd16};
ram[41374] = {-9'd13,-10'd13};
ram[41375] = {-9'd10,-10'd10};
ram[41376] = {-9'd7,-10'd7};
ram[41377] = {-9'd4,-10'd4};
ram[41378] = {9'd0,10'd0};
ram[41379] = {9'd3,10'd3};
ram[41380] = {9'd6,10'd6};
ram[41381] = {9'd9,10'd9};
ram[41382] = {9'd12,10'd12};
ram[41383] = {9'd15,10'd15};
ram[41384] = {9'd18,10'd18};
ram[41385] = {9'd21,10'd21};
ram[41386] = {9'd25,10'd25};
ram[41387] = {9'd28,10'd28};
ram[41388] = {9'd31,10'd31};
ram[41389] = {9'd34,10'd34};
ram[41390] = {9'd37,10'd37};
ram[41391] = {9'd40,10'd40};
ram[41392] = {9'd43,10'd43};
ram[41393] = {9'd47,10'd47};
ram[41394] = {9'd50,10'd50};
ram[41395] = {9'd53,10'd53};
ram[41396] = {9'd56,10'd56};
ram[41397] = {9'd59,10'd59};
ram[41398] = {9'd62,10'd62};
ram[41399] = {9'd65,10'd65};
ram[41400] = {9'd69,10'd69};
ram[41401] = {9'd72,10'd72};
ram[41402] = {9'd75,10'd75};
ram[41403] = {9'd78,10'd78};
ram[41404] = {9'd81,10'd81};
ram[41405] = {9'd84,10'd84};
ram[41406] = {9'd87,10'd87};
ram[41407] = {9'd91,10'd91};
ram[41408] = {9'd94,10'd94};
ram[41409] = {9'd97,10'd97};
ram[41410] = {-9'd100,10'd100};
ram[41411] = {-9'd97,10'd103};
ram[41412] = {-9'd94,10'd106};
ram[41413] = {-9'd91,10'd109};
ram[41414] = {-9'd88,10'd113};
ram[41415] = {-9'd85,10'd116};
ram[41416] = {-9'd81,10'd119};
ram[41417] = {-9'd78,10'd122};
ram[41418] = {-9'd75,10'd125};
ram[41419] = {-9'd72,10'd128};
ram[41420] = {-9'd69,10'd131};
ram[41421] = {-9'd66,10'd135};
ram[41422] = {-9'd63,10'd138};
ram[41423] = {-9'd59,10'd141};
ram[41424] = {-9'd56,10'd144};
ram[41425] = {-9'd53,10'd147};
ram[41426] = {-9'd50,10'd150};
ram[41427] = {-9'd47,10'd153};
ram[41428] = {-9'd44,10'd157};
ram[41429] = {-9'd41,10'd160};
ram[41430] = {-9'd37,10'd163};
ram[41431] = {-9'd34,10'd166};
ram[41432] = {-9'd31,10'd169};
ram[41433] = {-9'd28,10'd172};
ram[41434] = {-9'd25,10'd175};
ram[41435] = {-9'd22,10'd179};
ram[41436] = {-9'd19,10'd182};
ram[41437] = {-9'd15,10'd185};
ram[41438] = {-9'd12,10'd188};
ram[41439] = {-9'd9,10'd191};
ram[41440] = {-9'd6,10'd194};
ram[41441] = {-9'd3,10'd197};
ram[41442] = {9'd0,10'd201};
ram[41443] = {9'd3,10'd204};
ram[41444] = {9'd7,10'd207};
ram[41445] = {9'd10,10'd210};
ram[41446] = {9'd13,10'd213};
ram[41447] = {9'd16,10'd216};
ram[41448] = {9'd19,10'd219};
ram[41449] = {9'd22,10'd223};
ram[41450] = {9'd25,10'd226};
ram[41451] = {9'd29,10'd229};
ram[41452] = {9'd32,10'd232};
ram[41453] = {9'd35,10'd235};
ram[41454] = {9'd38,10'd238};
ram[41455] = {9'd41,10'd241};
ram[41456] = {9'd44,10'd245};
ram[41457] = {9'd47,10'd248};
ram[41458] = {9'd51,10'd251};
ram[41459] = {9'd54,10'd254};
ram[41460] = {9'd57,10'd257};
ram[41461] = {9'd60,10'd260};
ram[41462] = {9'd63,10'd263};
ram[41463] = {9'd66,10'd267};
ram[41464] = {9'd69,10'd270};
ram[41465] = {9'd73,10'd273};
ram[41466] = {9'd76,10'd276};
ram[41467] = {9'd79,10'd279};
ram[41468] = {9'd82,10'd282};
ram[41469] = {9'd85,10'd285};
ram[41470] = {9'd88,10'd289};
ram[41471] = {9'd91,10'd292};
ram[41472] = {9'd91,10'd292};
ram[41473] = {9'd95,10'd295};
ram[41474] = {9'd98,10'd298};
ram[41475] = {-9'd99,10'd301};
ram[41476] = {-9'd96,10'd304};
ram[41477] = {-9'd93,10'd307};
ram[41478] = {-9'd90,10'd311};
ram[41479] = {-9'd87,10'd314};
ram[41480] = {-9'd84,10'd317};
ram[41481] = {-9'd81,10'd320};
ram[41482] = {-9'd77,10'd323};
ram[41483] = {-9'd74,10'd326};
ram[41484] = {-9'd71,10'd329};
ram[41485] = {-9'd68,10'd333};
ram[41486] = {-9'd65,10'd336};
ram[41487] = {-9'd62,10'd339};
ram[41488] = {-9'd59,10'd342};
ram[41489] = {-9'd55,10'd345};
ram[41490] = {-9'd52,10'd348};
ram[41491] = {-9'd49,10'd351};
ram[41492] = {-9'd46,10'd354};
ram[41493] = {-9'd43,10'd358};
ram[41494] = {-9'd40,10'd361};
ram[41495] = {-9'd37,10'd364};
ram[41496] = {-9'd33,10'd367};
ram[41497] = {-9'd30,10'd370};
ram[41498] = {-9'd27,10'd373};
ram[41499] = {-9'd24,10'd376};
ram[41500] = {-9'd21,10'd380};
ram[41501] = {-9'd18,10'd383};
ram[41502] = {-9'd15,10'd386};
ram[41503] = {-9'd11,10'd389};
ram[41504] = {-9'd8,10'd392};
ram[41505] = {-9'd5,10'd395};
ram[41506] = {-9'd2,10'd398};
ram[41507] = {9'd1,-10'd399};
ram[41508] = {9'd4,-10'd396};
ram[41509] = {9'd7,-10'd393};
ram[41510] = {9'd10,-10'd390};
ram[41511] = {9'd14,-10'd387};
ram[41512] = {9'd17,-10'd384};
ram[41513] = {9'd20,-10'd381};
ram[41514] = {9'd23,-10'd377};
ram[41515] = {9'd26,-10'd374};
ram[41516] = {9'd29,-10'd371};
ram[41517] = {9'd32,-10'd368};
ram[41518] = {9'd36,-10'd365};
ram[41519] = {9'd39,-10'd362};
ram[41520] = {9'd42,-10'd359};
ram[41521] = {9'd45,-10'd355};
ram[41522] = {9'd48,-10'd352};
ram[41523] = {9'd51,-10'd349};
ram[41524] = {9'd54,-10'd346};
ram[41525] = {9'd58,-10'd343};
ram[41526] = {9'd61,-10'd340};
ram[41527] = {9'd64,-10'd337};
ram[41528] = {9'd67,-10'd334};
ram[41529] = {9'd70,-10'd330};
ram[41530] = {9'd73,-10'd327};
ram[41531] = {9'd76,-10'd324};
ram[41532] = {9'd80,-10'd321};
ram[41533] = {9'd83,-10'd318};
ram[41534] = {9'd86,-10'd315};
ram[41535] = {9'd89,-10'd312};
ram[41536] = {9'd92,-10'd308};
ram[41537] = {9'd95,-10'd305};
ram[41538] = {9'd98,-10'd302};
ram[41539] = {-9'd99,-10'd299};
ram[41540] = {-9'd96,-10'd296};
ram[41541] = {-9'd92,-10'd293};
ram[41542] = {-9'd89,-10'd290};
ram[41543] = {-9'd86,-10'd286};
ram[41544] = {-9'd83,-10'd283};
ram[41545] = {-9'd80,-10'd280};
ram[41546] = {-9'd77,-10'd277};
ram[41547] = {-9'd74,-10'd274};
ram[41548] = {-9'd70,-10'd271};
ram[41549] = {-9'd67,-10'd268};
ram[41550] = {-9'd64,-10'd264};
ram[41551] = {-9'd61,-10'd261};
ram[41552] = {-9'd58,-10'd258};
ram[41553] = {-9'd55,-10'd255};
ram[41554] = {-9'd52,-10'd252};
ram[41555] = {-9'd48,-10'd249};
ram[41556] = {-9'd45,-10'd246};
ram[41557] = {-9'd42,-10'd242};
ram[41558] = {-9'd39,-10'd239};
ram[41559] = {-9'd36,-10'd236};
ram[41560] = {-9'd33,-10'd233};
ram[41561] = {-9'd30,-10'd230};
ram[41562] = {-9'd26,-10'd227};
ram[41563] = {-9'd23,-10'd224};
ram[41564] = {-9'd20,-10'd220};
ram[41565] = {-9'd17,-10'd217};
ram[41566] = {-9'd14,-10'd214};
ram[41567] = {-9'd11,-10'd211};
ram[41568] = {-9'd8,-10'd208};
ram[41569] = {-9'd4,-10'd205};
ram[41570] = {-9'd1,-10'd202};
ram[41571] = {9'd2,-10'd198};
ram[41572] = {9'd5,-10'd195};
ram[41573] = {9'd8,-10'd192};
ram[41574] = {9'd11,-10'd189};
ram[41575] = {9'd14,-10'd186};
ram[41576] = {9'd18,-10'd183};
ram[41577] = {9'd21,-10'd180};
ram[41578] = {9'd24,-10'd176};
ram[41579] = {9'd27,-10'd173};
ram[41580] = {9'd30,-10'd170};
ram[41581] = {9'd33,-10'd167};
ram[41582] = {9'd36,-10'd164};
ram[41583] = {9'd40,-10'd161};
ram[41584] = {9'd43,-10'd158};
ram[41585] = {9'd46,-10'd154};
ram[41586] = {9'd49,-10'd151};
ram[41587] = {9'd52,-10'd148};
ram[41588] = {9'd55,-10'd145};
ram[41589] = {9'd58,-10'd142};
ram[41590] = {9'd62,-10'd139};
ram[41591] = {9'd65,-10'd136};
ram[41592] = {9'd68,-10'd132};
ram[41593] = {9'd71,-10'd129};
ram[41594] = {9'd74,-10'd126};
ram[41595] = {9'd77,-10'd123};
ram[41596] = {9'd80,-10'd120};
ram[41597] = {9'd84,-10'd117};
ram[41598] = {9'd87,-10'd114};
ram[41599] = {9'd90,-10'd110};
ram[41600] = {9'd90,-10'd110};
ram[41601] = {9'd93,-10'd107};
ram[41602] = {9'd96,-10'd104};
ram[41603] = {9'd99,-10'd101};
ram[41604] = {-9'd98,-10'd98};
ram[41605] = {-9'd95,-10'd95};
ram[41606] = {-9'd92,-10'd92};
ram[41607] = {-9'd88,-10'd88};
ram[41608] = {-9'd85,-10'd85};
ram[41609] = {-9'd82,-10'd82};
ram[41610] = {-9'd79,-10'd79};
ram[41611] = {-9'd76,-10'd76};
ram[41612] = {-9'd73,-10'd73};
ram[41613] = {-9'd70,-10'd70};
ram[41614] = {-9'd66,-10'd66};
ram[41615] = {-9'd63,-10'd63};
ram[41616] = {-9'd60,-10'd60};
ram[41617] = {-9'd57,-10'd57};
ram[41618] = {-9'd54,-10'd54};
ram[41619] = {-9'd51,-10'd51};
ram[41620] = {-9'd48,-10'd48};
ram[41621] = {-9'd44,-10'd44};
ram[41622] = {-9'd41,-10'd41};
ram[41623] = {-9'd38,-10'd38};
ram[41624] = {-9'd35,-10'd35};
ram[41625] = {-9'd32,-10'd32};
ram[41626] = {-9'd29,-10'd29};
ram[41627] = {-9'd26,-10'd26};
ram[41628] = {-9'd22,-10'd22};
ram[41629] = {-9'd19,-10'd19};
ram[41630] = {-9'd16,-10'd16};
ram[41631] = {-9'd13,-10'd13};
ram[41632] = {-9'd10,-10'd10};
ram[41633] = {-9'd7,-10'd7};
ram[41634] = {-9'd4,-10'd4};
ram[41635] = {9'd0,10'd0};
ram[41636] = {9'd3,10'd3};
ram[41637] = {9'd6,10'd6};
ram[41638] = {9'd9,10'd9};
ram[41639] = {9'd12,10'd12};
ram[41640] = {9'd15,10'd15};
ram[41641] = {9'd18,10'd18};
ram[41642] = {9'd21,10'd21};
ram[41643] = {9'd25,10'd25};
ram[41644] = {9'd28,10'd28};
ram[41645] = {9'd31,10'd31};
ram[41646] = {9'd34,10'd34};
ram[41647] = {9'd37,10'd37};
ram[41648] = {9'd40,10'd40};
ram[41649] = {9'd43,10'd43};
ram[41650] = {9'd47,10'd47};
ram[41651] = {9'd50,10'd50};
ram[41652] = {9'd53,10'd53};
ram[41653] = {9'd56,10'd56};
ram[41654] = {9'd59,10'd59};
ram[41655] = {9'd62,10'd62};
ram[41656] = {9'd65,10'd65};
ram[41657] = {9'd69,10'd69};
ram[41658] = {9'd72,10'd72};
ram[41659] = {9'd75,10'd75};
ram[41660] = {9'd78,10'd78};
ram[41661] = {9'd81,10'd81};
ram[41662] = {9'd84,10'd84};
ram[41663] = {9'd87,10'd87};
ram[41664] = {9'd91,10'd91};
ram[41665] = {9'd94,10'd94};
ram[41666] = {9'd97,10'd97};
ram[41667] = {-9'd100,10'd100};
ram[41668] = {-9'd97,10'd103};
ram[41669] = {-9'd94,10'd106};
ram[41670] = {-9'd91,10'd109};
ram[41671] = {-9'd88,10'd113};
ram[41672] = {-9'd85,10'd116};
ram[41673] = {-9'd81,10'd119};
ram[41674] = {-9'd78,10'd122};
ram[41675] = {-9'd75,10'd125};
ram[41676] = {-9'd72,10'd128};
ram[41677] = {-9'd69,10'd131};
ram[41678] = {-9'd66,10'd135};
ram[41679] = {-9'd63,10'd138};
ram[41680] = {-9'd59,10'd141};
ram[41681] = {-9'd56,10'd144};
ram[41682] = {-9'd53,10'd147};
ram[41683] = {-9'd50,10'd150};
ram[41684] = {-9'd47,10'd153};
ram[41685] = {-9'd44,10'd157};
ram[41686] = {-9'd41,10'd160};
ram[41687] = {-9'd37,10'd163};
ram[41688] = {-9'd34,10'd166};
ram[41689] = {-9'd31,10'd169};
ram[41690] = {-9'd28,10'd172};
ram[41691] = {-9'd25,10'd175};
ram[41692] = {-9'd22,10'd179};
ram[41693] = {-9'd19,10'd182};
ram[41694] = {-9'd15,10'd185};
ram[41695] = {-9'd12,10'd188};
ram[41696] = {-9'd9,10'd191};
ram[41697] = {-9'd6,10'd194};
ram[41698] = {-9'd3,10'd197};
ram[41699] = {9'd0,10'd201};
ram[41700] = {9'd3,10'd204};
ram[41701] = {9'd7,10'd207};
ram[41702] = {9'd10,10'd210};
ram[41703] = {9'd13,10'd213};
ram[41704] = {9'd16,10'd216};
ram[41705] = {9'd19,10'd219};
ram[41706] = {9'd22,10'd223};
ram[41707] = {9'd25,10'd226};
ram[41708] = {9'd29,10'd229};
ram[41709] = {9'd32,10'd232};
ram[41710] = {9'd35,10'd235};
ram[41711] = {9'd38,10'd238};
ram[41712] = {9'd41,10'd241};
ram[41713] = {9'd44,10'd245};
ram[41714] = {9'd47,10'd248};
ram[41715] = {9'd51,10'd251};
ram[41716] = {9'd54,10'd254};
ram[41717] = {9'd57,10'd257};
ram[41718] = {9'd60,10'd260};
ram[41719] = {9'd63,10'd263};
ram[41720] = {9'd66,10'd267};
ram[41721] = {9'd69,10'd270};
ram[41722] = {9'd73,10'd273};
ram[41723] = {9'd76,10'd276};
ram[41724] = {9'd79,10'd279};
ram[41725] = {9'd82,10'd282};
ram[41726] = {9'd85,10'd285};
ram[41727] = {9'd88,10'd289};
ram[41728] = {9'd88,10'd289};
ram[41729] = {9'd91,10'd292};
ram[41730] = {9'd95,10'd295};
ram[41731] = {9'd98,10'd298};
ram[41732] = {-9'd99,10'd301};
ram[41733] = {-9'd96,10'd304};
ram[41734] = {-9'd93,10'd307};
ram[41735] = {-9'd90,10'd311};
ram[41736] = {-9'd87,10'd314};
ram[41737] = {-9'd84,10'd317};
ram[41738] = {-9'd81,10'd320};
ram[41739] = {-9'd77,10'd323};
ram[41740] = {-9'd74,10'd326};
ram[41741] = {-9'd71,10'd329};
ram[41742] = {-9'd68,10'd333};
ram[41743] = {-9'd65,10'd336};
ram[41744] = {-9'd62,10'd339};
ram[41745] = {-9'd59,10'd342};
ram[41746] = {-9'd55,10'd345};
ram[41747] = {-9'd52,10'd348};
ram[41748] = {-9'd49,10'd351};
ram[41749] = {-9'd46,10'd354};
ram[41750] = {-9'd43,10'd358};
ram[41751] = {-9'd40,10'd361};
ram[41752] = {-9'd37,10'd364};
ram[41753] = {-9'd33,10'd367};
ram[41754] = {-9'd30,10'd370};
ram[41755] = {-9'd27,10'd373};
ram[41756] = {-9'd24,10'd376};
ram[41757] = {-9'd21,10'd380};
ram[41758] = {-9'd18,10'd383};
ram[41759] = {-9'd15,10'd386};
ram[41760] = {-9'd11,10'd389};
ram[41761] = {-9'd8,10'd392};
ram[41762] = {-9'd5,10'd395};
ram[41763] = {-9'd2,10'd398};
ram[41764] = {9'd1,-10'd399};
ram[41765] = {9'd4,-10'd396};
ram[41766] = {9'd7,-10'd393};
ram[41767] = {9'd10,-10'd390};
ram[41768] = {9'd14,-10'd387};
ram[41769] = {9'd17,-10'd384};
ram[41770] = {9'd20,-10'd381};
ram[41771] = {9'd23,-10'd377};
ram[41772] = {9'd26,-10'd374};
ram[41773] = {9'd29,-10'd371};
ram[41774] = {9'd32,-10'd368};
ram[41775] = {9'd36,-10'd365};
ram[41776] = {9'd39,-10'd362};
ram[41777] = {9'd42,-10'd359};
ram[41778] = {9'd45,-10'd355};
ram[41779] = {9'd48,-10'd352};
ram[41780] = {9'd51,-10'd349};
ram[41781] = {9'd54,-10'd346};
ram[41782] = {9'd58,-10'd343};
ram[41783] = {9'd61,-10'd340};
ram[41784] = {9'd64,-10'd337};
ram[41785] = {9'd67,-10'd334};
ram[41786] = {9'd70,-10'd330};
ram[41787] = {9'd73,-10'd327};
ram[41788] = {9'd76,-10'd324};
ram[41789] = {9'd80,-10'd321};
ram[41790] = {9'd83,-10'd318};
ram[41791] = {9'd86,-10'd315};
ram[41792] = {9'd89,-10'd312};
ram[41793] = {9'd92,-10'd308};
ram[41794] = {9'd95,-10'd305};
ram[41795] = {9'd98,-10'd302};
ram[41796] = {-9'd99,-10'd299};
ram[41797] = {-9'd96,-10'd296};
ram[41798] = {-9'd92,-10'd293};
ram[41799] = {-9'd89,-10'd290};
ram[41800] = {-9'd86,-10'd286};
ram[41801] = {-9'd83,-10'd283};
ram[41802] = {-9'd80,-10'd280};
ram[41803] = {-9'd77,-10'd277};
ram[41804] = {-9'd74,-10'd274};
ram[41805] = {-9'd70,-10'd271};
ram[41806] = {-9'd67,-10'd268};
ram[41807] = {-9'd64,-10'd264};
ram[41808] = {-9'd61,-10'd261};
ram[41809] = {-9'd58,-10'd258};
ram[41810] = {-9'd55,-10'd255};
ram[41811] = {-9'd52,-10'd252};
ram[41812] = {-9'd48,-10'd249};
ram[41813] = {-9'd45,-10'd246};
ram[41814] = {-9'd42,-10'd242};
ram[41815] = {-9'd39,-10'd239};
ram[41816] = {-9'd36,-10'd236};
ram[41817] = {-9'd33,-10'd233};
ram[41818] = {-9'd30,-10'd230};
ram[41819] = {-9'd26,-10'd227};
ram[41820] = {-9'd23,-10'd224};
ram[41821] = {-9'd20,-10'd220};
ram[41822] = {-9'd17,-10'd217};
ram[41823] = {-9'd14,-10'd214};
ram[41824] = {-9'd11,-10'd211};
ram[41825] = {-9'd8,-10'd208};
ram[41826] = {-9'd4,-10'd205};
ram[41827] = {-9'd1,-10'd202};
ram[41828] = {9'd2,-10'd198};
ram[41829] = {9'd5,-10'd195};
ram[41830] = {9'd8,-10'd192};
ram[41831] = {9'd11,-10'd189};
ram[41832] = {9'd14,-10'd186};
ram[41833] = {9'd18,-10'd183};
ram[41834] = {9'd21,-10'd180};
ram[41835] = {9'd24,-10'd176};
ram[41836] = {9'd27,-10'd173};
ram[41837] = {9'd30,-10'd170};
ram[41838] = {9'd33,-10'd167};
ram[41839] = {9'd36,-10'd164};
ram[41840] = {9'd40,-10'd161};
ram[41841] = {9'd43,-10'd158};
ram[41842] = {9'd46,-10'd154};
ram[41843] = {9'd49,-10'd151};
ram[41844] = {9'd52,-10'd148};
ram[41845] = {9'd55,-10'd145};
ram[41846] = {9'd58,-10'd142};
ram[41847] = {9'd62,-10'd139};
ram[41848] = {9'd65,-10'd136};
ram[41849] = {9'd68,-10'd132};
ram[41850] = {9'd71,-10'd129};
ram[41851] = {9'd74,-10'd126};
ram[41852] = {9'd77,-10'd123};
ram[41853] = {9'd80,-10'd120};
ram[41854] = {9'd84,-10'd117};
ram[41855] = {9'd87,-10'd114};
ram[41856] = {9'd87,-10'd114};
ram[41857] = {9'd90,-10'd110};
ram[41858] = {9'd93,-10'd107};
ram[41859] = {9'd96,-10'd104};
ram[41860] = {9'd99,-10'd101};
ram[41861] = {-9'd98,-10'd98};
ram[41862] = {-9'd95,-10'd95};
ram[41863] = {-9'd92,-10'd92};
ram[41864] = {-9'd88,-10'd88};
ram[41865] = {-9'd85,-10'd85};
ram[41866] = {-9'd82,-10'd82};
ram[41867] = {-9'd79,-10'd79};
ram[41868] = {-9'd76,-10'd76};
ram[41869] = {-9'd73,-10'd73};
ram[41870] = {-9'd70,-10'd70};
ram[41871] = {-9'd66,-10'd66};
ram[41872] = {-9'd63,-10'd63};
ram[41873] = {-9'd60,-10'd60};
ram[41874] = {-9'd57,-10'd57};
ram[41875] = {-9'd54,-10'd54};
ram[41876] = {-9'd51,-10'd51};
ram[41877] = {-9'd48,-10'd48};
ram[41878] = {-9'd44,-10'd44};
ram[41879] = {-9'd41,-10'd41};
ram[41880] = {-9'd38,-10'd38};
ram[41881] = {-9'd35,-10'd35};
ram[41882] = {-9'd32,-10'd32};
ram[41883] = {-9'd29,-10'd29};
ram[41884] = {-9'd26,-10'd26};
ram[41885] = {-9'd22,-10'd22};
ram[41886] = {-9'd19,-10'd19};
ram[41887] = {-9'd16,-10'd16};
ram[41888] = {-9'd13,-10'd13};
ram[41889] = {-9'd10,-10'd10};
ram[41890] = {-9'd7,-10'd7};
ram[41891] = {-9'd4,-10'd4};
ram[41892] = {9'd0,10'd0};
ram[41893] = {9'd3,10'd3};
ram[41894] = {9'd6,10'd6};
ram[41895] = {9'd9,10'd9};
ram[41896] = {9'd12,10'd12};
ram[41897] = {9'd15,10'd15};
ram[41898] = {9'd18,10'd18};
ram[41899] = {9'd21,10'd21};
ram[41900] = {9'd25,10'd25};
ram[41901] = {9'd28,10'd28};
ram[41902] = {9'd31,10'd31};
ram[41903] = {9'd34,10'd34};
ram[41904] = {9'd37,10'd37};
ram[41905] = {9'd40,10'd40};
ram[41906] = {9'd43,10'd43};
ram[41907] = {9'd47,10'd47};
ram[41908] = {9'd50,10'd50};
ram[41909] = {9'd53,10'd53};
ram[41910] = {9'd56,10'd56};
ram[41911] = {9'd59,10'd59};
ram[41912] = {9'd62,10'd62};
ram[41913] = {9'd65,10'd65};
ram[41914] = {9'd69,10'd69};
ram[41915] = {9'd72,10'd72};
ram[41916] = {9'd75,10'd75};
ram[41917] = {9'd78,10'd78};
ram[41918] = {9'd81,10'd81};
ram[41919] = {9'd84,10'd84};
ram[41920] = {9'd87,10'd87};
ram[41921] = {9'd91,10'd91};
ram[41922] = {9'd94,10'd94};
ram[41923] = {9'd97,10'd97};
ram[41924] = {-9'd100,10'd100};
ram[41925] = {-9'd97,10'd103};
ram[41926] = {-9'd94,10'd106};
ram[41927] = {-9'd91,10'd109};
ram[41928] = {-9'd88,10'd113};
ram[41929] = {-9'd85,10'd116};
ram[41930] = {-9'd81,10'd119};
ram[41931] = {-9'd78,10'd122};
ram[41932] = {-9'd75,10'd125};
ram[41933] = {-9'd72,10'd128};
ram[41934] = {-9'd69,10'd131};
ram[41935] = {-9'd66,10'd135};
ram[41936] = {-9'd63,10'd138};
ram[41937] = {-9'd59,10'd141};
ram[41938] = {-9'd56,10'd144};
ram[41939] = {-9'd53,10'd147};
ram[41940] = {-9'd50,10'd150};
ram[41941] = {-9'd47,10'd153};
ram[41942] = {-9'd44,10'd157};
ram[41943] = {-9'd41,10'd160};
ram[41944] = {-9'd37,10'd163};
ram[41945] = {-9'd34,10'd166};
ram[41946] = {-9'd31,10'd169};
ram[41947] = {-9'd28,10'd172};
ram[41948] = {-9'd25,10'd175};
ram[41949] = {-9'd22,10'd179};
ram[41950] = {-9'd19,10'd182};
ram[41951] = {-9'd15,10'd185};
ram[41952] = {-9'd12,10'd188};
ram[41953] = {-9'd9,10'd191};
ram[41954] = {-9'd6,10'd194};
ram[41955] = {-9'd3,10'd197};
ram[41956] = {9'd0,10'd201};
ram[41957] = {9'd3,10'd204};
ram[41958] = {9'd7,10'd207};
ram[41959] = {9'd10,10'd210};
ram[41960] = {9'd13,10'd213};
ram[41961] = {9'd16,10'd216};
ram[41962] = {9'd19,10'd219};
ram[41963] = {9'd22,10'd223};
ram[41964] = {9'd25,10'd226};
ram[41965] = {9'd29,10'd229};
ram[41966] = {9'd32,10'd232};
ram[41967] = {9'd35,10'd235};
ram[41968] = {9'd38,10'd238};
ram[41969] = {9'd41,10'd241};
ram[41970] = {9'd44,10'd245};
ram[41971] = {9'd47,10'd248};
ram[41972] = {9'd51,10'd251};
ram[41973] = {9'd54,10'd254};
ram[41974] = {9'd57,10'd257};
ram[41975] = {9'd60,10'd260};
ram[41976] = {9'd63,10'd263};
ram[41977] = {9'd66,10'd267};
ram[41978] = {9'd69,10'd270};
ram[41979] = {9'd73,10'd273};
ram[41980] = {9'd76,10'd276};
ram[41981] = {9'd79,10'd279};
ram[41982] = {9'd82,10'd282};
ram[41983] = {9'd85,10'd285};
ram[41984] = {9'd85,10'd285};
ram[41985] = {9'd88,10'd289};
ram[41986] = {9'd91,10'd292};
ram[41987] = {9'd95,10'd295};
ram[41988] = {9'd98,10'd298};
ram[41989] = {-9'd99,10'd301};
ram[41990] = {-9'd96,10'd304};
ram[41991] = {-9'd93,10'd307};
ram[41992] = {-9'd90,10'd311};
ram[41993] = {-9'd87,10'd314};
ram[41994] = {-9'd84,10'd317};
ram[41995] = {-9'd81,10'd320};
ram[41996] = {-9'd77,10'd323};
ram[41997] = {-9'd74,10'd326};
ram[41998] = {-9'd71,10'd329};
ram[41999] = {-9'd68,10'd333};
ram[42000] = {-9'd65,10'd336};
ram[42001] = {-9'd62,10'd339};
ram[42002] = {-9'd59,10'd342};
ram[42003] = {-9'd55,10'd345};
ram[42004] = {-9'd52,10'd348};
ram[42005] = {-9'd49,10'd351};
ram[42006] = {-9'd46,10'd354};
ram[42007] = {-9'd43,10'd358};
ram[42008] = {-9'd40,10'd361};
ram[42009] = {-9'd37,10'd364};
ram[42010] = {-9'd33,10'd367};
ram[42011] = {-9'd30,10'd370};
ram[42012] = {-9'd27,10'd373};
ram[42013] = {-9'd24,10'd376};
ram[42014] = {-9'd21,10'd380};
ram[42015] = {-9'd18,10'd383};
ram[42016] = {-9'd15,10'd386};
ram[42017] = {-9'd11,10'd389};
ram[42018] = {-9'd8,10'd392};
ram[42019] = {-9'd5,10'd395};
ram[42020] = {-9'd2,10'd398};
ram[42021] = {9'd1,-10'd399};
ram[42022] = {9'd4,-10'd396};
ram[42023] = {9'd7,-10'd393};
ram[42024] = {9'd10,-10'd390};
ram[42025] = {9'd14,-10'd387};
ram[42026] = {9'd17,-10'd384};
ram[42027] = {9'd20,-10'd381};
ram[42028] = {9'd23,-10'd377};
ram[42029] = {9'd26,-10'd374};
ram[42030] = {9'd29,-10'd371};
ram[42031] = {9'd32,-10'd368};
ram[42032] = {9'd36,-10'd365};
ram[42033] = {9'd39,-10'd362};
ram[42034] = {9'd42,-10'd359};
ram[42035] = {9'd45,-10'd355};
ram[42036] = {9'd48,-10'd352};
ram[42037] = {9'd51,-10'd349};
ram[42038] = {9'd54,-10'd346};
ram[42039] = {9'd58,-10'd343};
ram[42040] = {9'd61,-10'd340};
ram[42041] = {9'd64,-10'd337};
ram[42042] = {9'd67,-10'd334};
ram[42043] = {9'd70,-10'd330};
ram[42044] = {9'd73,-10'd327};
ram[42045] = {9'd76,-10'd324};
ram[42046] = {9'd80,-10'd321};
ram[42047] = {9'd83,-10'd318};
ram[42048] = {9'd86,-10'd315};
ram[42049] = {9'd89,-10'd312};
ram[42050] = {9'd92,-10'd308};
ram[42051] = {9'd95,-10'd305};
ram[42052] = {9'd98,-10'd302};
ram[42053] = {-9'd99,-10'd299};
ram[42054] = {-9'd96,-10'd296};
ram[42055] = {-9'd92,-10'd293};
ram[42056] = {-9'd89,-10'd290};
ram[42057] = {-9'd86,-10'd286};
ram[42058] = {-9'd83,-10'd283};
ram[42059] = {-9'd80,-10'd280};
ram[42060] = {-9'd77,-10'd277};
ram[42061] = {-9'd74,-10'd274};
ram[42062] = {-9'd70,-10'd271};
ram[42063] = {-9'd67,-10'd268};
ram[42064] = {-9'd64,-10'd264};
ram[42065] = {-9'd61,-10'd261};
ram[42066] = {-9'd58,-10'd258};
ram[42067] = {-9'd55,-10'd255};
ram[42068] = {-9'd52,-10'd252};
ram[42069] = {-9'd48,-10'd249};
ram[42070] = {-9'd45,-10'd246};
ram[42071] = {-9'd42,-10'd242};
ram[42072] = {-9'd39,-10'd239};
ram[42073] = {-9'd36,-10'd236};
ram[42074] = {-9'd33,-10'd233};
ram[42075] = {-9'd30,-10'd230};
ram[42076] = {-9'd26,-10'd227};
ram[42077] = {-9'd23,-10'd224};
ram[42078] = {-9'd20,-10'd220};
ram[42079] = {-9'd17,-10'd217};
ram[42080] = {-9'd14,-10'd214};
ram[42081] = {-9'd11,-10'd211};
ram[42082] = {-9'd8,-10'd208};
ram[42083] = {-9'd4,-10'd205};
ram[42084] = {-9'd1,-10'd202};
ram[42085] = {9'd2,-10'd198};
ram[42086] = {9'd5,-10'd195};
ram[42087] = {9'd8,-10'd192};
ram[42088] = {9'd11,-10'd189};
ram[42089] = {9'd14,-10'd186};
ram[42090] = {9'd18,-10'd183};
ram[42091] = {9'd21,-10'd180};
ram[42092] = {9'd24,-10'd176};
ram[42093] = {9'd27,-10'd173};
ram[42094] = {9'd30,-10'd170};
ram[42095] = {9'd33,-10'd167};
ram[42096] = {9'd36,-10'd164};
ram[42097] = {9'd40,-10'd161};
ram[42098] = {9'd43,-10'd158};
ram[42099] = {9'd46,-10'd154};
ram[42100] = {9'd49,-10'd151};
ram[42101] = {9'd52,-10'd148};
ram[42102] = {9'd55,-10'd145};
ram[42103] = {9'd58,-10'd142};
ram[42104] = {9'd62,-10'd139};
ram[42105] = {9'd65,-10'd136};
ram[42106] = {9'd68,-10'd132};
ram[42107] = {9'd71,-10'd129};
ram[42108] = {9'd74,-10'd126};
ram[42109] = {9'd77,-10'd123};
ram[42110] = {9'd80,-10'd120};
ram[42111] = {9'd84,-10'd117};
ram[42112] = {9'd84,-10'd117};
ram[42113] = {9'd87,-10'd114};
ram[42114] = {9'd90,-10'd110};
ram[42115] = {9'd93,-10'd107};
ram[42116] = {9'd96,-10'd104};
ram[42117] = {9'd99,-10'd101};
ram[42118] = {-9'd98,-10'd98};
ram[42119] = {-9'd95,-10'd95};
ram[42120] = {-9'd92,-10'd92};
ram[42121] = {-9'd88,-10'd88};
ram[42122] = {-9'd85,-10'd85};
ram[42123] = {-9'd82,-10'd82};
ram[42124] = {-9'd79,-10'd79};
ram[42125] = {-9'd76,-10'd76};
ram[42126] = {-9'd73,-10'd73};
ram[42127] = {-9'd70,-10'd70};
ram[42128] = {-9'd66,-10'd66};
ram[42129] = {-9'd63,-10'd63};
ram[42130] = {-9'd60,-10'd60};
ram[42131] = {-9'd57,-10'd57};
ram[42132] = {-9'd54,-10'd54};
ram[42133] = {-9'd51,-10'd51};
ram[42134] = {-9'd48,-10'd48};
ram[42135] = {-9'd44,-10'd44};
ram[42136] = {-9'd41,-10'd41};
ram[42137] = {-9'd38,-10'd38};
ram[42138] = {-9'd35,-10'd35};
ram[42139] = {-9'd32,-10'd32};
ram[42140] = {-9'd29,-10'd29};
ram[42141] = {-9'd26,-10'd26};
ram[42142] = {-9'd22,-10'd22};
ram[42143] = {-9'd19,-10'd19};
ram[42144] = {-9'd16,-10'd16};
ram[42145] = {-9'd13,-10'd13};
ram[42146] = {-9'd10,-10'd10};
ram[42147] = {-9'd7,-10'd7};
ram[42148] = {-9'd4,-10'd4};
ram[42149] = {9'd0,10'd0};
ram[42150] = {9'd3,10'd3};
ram[42151] = {9'd6,10'd6};
ram[42152] = {9'd9,10'd9};
ram[42153] = {9'd12,10'd12};
ram[42154] = {9'd15,10'd15};
ram[42155] = {9'd18,10'd18};
ram[42156] = {9'd21,10'd21};
ram[42157] = {9'd25,10'd25};
ram[42158] = {9'd28,10'd28};
ram[42159] = {9'd31,10'd31};
ram[42160] = {9'd34,10'd34};
ram[42161] = {9'd37,10'd37};
ram[42162] = {9'd40,10'd40};
ram[42163] = {9'd43,10'd43};
ram[42164] = {9'd47,10'd47};
ram[42165] = {9'd50,10'd50};
ram[42166] = {9'd53,10'd53};
ram[42167] = {9'd56,10'd56};
ram[42168] = {9'd59,10'd59};
ram[42169] = {9'd62,10'd62};
ram[42170] = {9'd65,10'd65};
ram[42171] = {9'd69,10'd69};
ram[42172] = {9'd72,10'd72};
ram[42173] = {9'd75,10'd75};
ram[42174] = {9'd78,10'd78};
ram[42175] = {9'd81,10'd81};
ram[42176] = {9'd84,10'd84};
ram[42177] = {9'd87,10'd87};
ram[42178] = {9'd91,10'd91};
ram[42179] = {9'd94,10'd94};
ram[42180] = {9'd97,10'd97};
ram[42181] = {-9'd100,10'd100};
ram[42182] = {-9'd97,10'd103};
ram[42183] = {-9'd94,10'd106};
ram[42184] = {-9'd91,10'd109};
ram[42185] = {-9'd88,10'd113};
ram[42186] = {-9'd85,10'd116};
ram[42187] = {-9'd81,10'd119};
ram[42188] = {-9'd78,10'd122};
ram[42189] = {-9'd75,10'd125};
ram[42190] = {-9'd72,10'd128};
ram[42191] = {-9'd69,10'd131};
ram[42192] = {-9'd66,10'd135};
ram[42193] = {-9'd63,10'd138};
ram[42194] = {-9'd59,10'd141};
ram[42195] = {-9'd56,10'd144};
ram[42196] = {-9'd53,10'd147};
ram[42197] = {-9'd50,10'd150};
ram[42198] = {-9'd47,10'd153};
ram[42199] = {-9'd44,10'd157};
ram[42200] = {-9'd41,10'd160};
ram[42201] = {-9'd37,10'd163};
ram[42202] = {-9'd34,10'd166};
ram[42203] = {-9'd31,10'd169};
ram[42204] = {-9'd28,10'd172};
ram[42205] = {-9'd25,10'd175};
ram[42206] = {-9'd22,10'd179};
ram[42207] = {-9'd19,10'd182};
ram[42208] = {-9'd15,10'd185};
ram[42209] = {-9'd12,10'd188};
ram[42210] = {-9'd9,10'd191};
ram[42211] = {-9'd6,10'd194};
ram[42212] = {-9'd3,10'd197};
ram[42213] = {9'd0,10'd201};
ram[42214] = {9'd3,10'd204};
ram[42215] = {9'd7,10'd207};
ram[42216] = {9'd10,10'd210};
ram[42217] = {9'd13,10'd213};
ram[42218] = {9'd16,10'd216};
ram[42219] = {9'd19,10'd219};
ram[42220] = {9'd22,10'd223};
ram[42221] = {9'd25,10'd226};
ram[42222] = {9'd29,10'd229};
ram[42223] = {9'd32,10'd232};
ram[42224] = {9'd35,10'd235};
ram[42225] = {9'd38,10'd238};
ram[42226] = {9'd41,10'd241};
ram[42227] = {9'd44,10'd245};
ram[42228] = {9'd47,10'd248};
ram[42229] = {9'd51,10'd251};
ram[42230] = {9'd54,10'd254};
ram[42231] = {9'd57,10'd257};
ram[42232] = {9'd60,10'd260};
ram[42233] = {9'd63,10'd263};
ram[42234] = {9'd66,10'd267};
ram[42235] = {9'd69,10'd270};
ram[42236] = {9'd73,10'd273};
ram[42237] = {9'd76,10'd276};
ram[42238] = {9'd79,10'd279};
ram[42239] = {9'd82,10'd282};
ram[42240] = {9'd82,10'd282};
ram[42241] = {9'd85,10'd285};
ram[42242] = {9'd88,10'd289};
ram[42243] = {9'd91,10'd292};
ram[42244] = {9'd95,10'd295};
ram[42245] = {9'd98,10'd298};
ram[42246] = {-9'd99,10'd301};
ram[42247] = {-9'd96,10'd304};
ram[42248] = {-9'd93,10'd307};
ram[42249] = {-9'd90,10'd311};
ram[42250] = {-9'd87,10'd314};
ram[42251] = {-9'd84,10'd317};
ram[42252] = {-9'd81,10'd320};
ram[42253] = {-9'd77,10'd323};
ram[42254] = {-9'd74,10'd326};
ram[42255] = {-9'd71,10'd329};
ram[42256] = {-9'd68,10'd333};
ram[42257] = {-9'd65,10'd336};
ram[42258] = {-9'd62,10'd339};
ram[42259] = {-9'd59,10'd342};
ram[42260] = {-9'd55,10'd345};
ram[42261] = {-9'd52,10'd348};
ram[42262] = {-9'd49,10'd351};
ram[42263] = {-9'd46,10'd354};
ram[42264] = {-9'd43,10'd358};
ram[42265] = {-9'd40,10'd361};
ram[42266] = {-9'd37,10'd364};
ram[42267] = {-9'd33,10'd367};
ram[42268] = {-9'd30,10'd370};
ram[42269] = {-9'd27,10'd373};
ram[42270] = {-9'd24,10'd376};
ram[42271] = {-9'd21,10'd380};
ram[42272] = {-9'd18,10'd383};
ram[42273] = {-9'd15,10'd386};
ram[42274] = {-9'd11,10'd389};
ram[42275] = {-9'd8,10'd392};
ram[42276] = {-9'd5,10'd395};
ram[42277] = {-9'd2,10'd398};
ram[42278] = {9'd1,-10'd399};
ram[42279] = {9'd4,-10'd396};
ram[42280] = {9'd7,-10'd393};
ram[42281] = {9'd10,-10'd390};
ram[42282] = {9'd14,-10'd387};
ram[42283] = {9'd17,-10'd384};
ram[42284] = {9'd20,-10'd381};
ram[42285] = {9'd23,-10'd377};
ram[42286] = {9'd26,-10'd374};
ram[42287] = {9'd29,-10'd371};
ram[42288] = {9'd32,-10'd368};
ram[42289] = {9'd36,-10'd365};
ram[42290] = {9'd39,-10'd362};
ram[42291] = {9'd42,-10'd359};
ram[42292] = {9'd45,-10'd355};
ram[42293] = {9'd48,-10'd352};
ram[42294] = {9'd51,-10'd349};
ram[42295] = {9'd54,-10'd346};
ram[42296] = {9'd58,-10'd343};
ram[42297] = {9'd61,-10'd340};
ram[42298] = {9'd64,-10'd337};
ram[42299] = {9'd67,-10'd334};
ram[42300] = {9'd70,-10'd330};
ram[42301] = {9'd73,-10'd327};
ram[42302] = {9'd76,-10'd324};
ram[42303] = {9'd80,-10'd321};
ram[42304] = {9'd83,-10'd318};
ram[42305] = {9'd86,-10'd315};
ram[42306] = {9'd89,-10'd312};
ram[42307] = {9'd92,-10'd308};
ram[42308] = {9'd95,-10'd305};
ram[42309] = {9'd98,-10'd302};
ram[42310] = {-9'd99,-10'd299};
ram[42311] = {-9'd96,-10'd296};
ram[42312] = {-9'd92,-10'd293};
ram[42313] = {-9'd89,-10'd290};
ram[42314] = {-9'd86,-10'd286};
ram[42315] = {-9'd83,-10'd283};
ram[42316] = {-9'd80,-10'd280};
ram[42317] = {-9'd77,-10'd277};
ram[42318] = {-9'd74,-10'd274};
ram[42319] = {-9'd70,-10'd271};
ram[42320] = {-9'd67,-10'd268};
ram[42321] = {-9'd64,-10'd264};
ram[42322] = {-9'd61,-10'd261};
ram[42323] = {-9'd58,-10'd258};
ram[42324] = {-9'd55,-10'd255};
ram[42325] = {-9'd52,-10'd252};
ram[42326] = {-9'd48,-10'd249};
ram[42327] = {-9'd45,-10'd246};
ram[42328] = {-9'd42,-10'd242};
ram[42329] = {-9'd39,-10'd239};
ram[42330] = {-9'd36,-10'd236};
ram[42331] = {-9'd33,-10'd233};
ram[42332] = {-9'd30,-10'd230};
ram[42333] = {-9'd26,-10'd227};
ram[42334] = {-9'd23,-10'd224};
ram[42335] = {-9'd20,-10'd220};
ram[42336] = {-9'd17,-10'd217};
ram[42337] = {-9'd14,-10'd214};
ram[42338] = {-9'd11,-10'd211};
ram[42339] = {-9'd8,-10'd208};
ram[42340] = {-9'd4,-10'd205};
ram[42341] = {-9'd1,-10'd202};
ram[42342] = {9'd2,-10'd198};
ram[42343] = {9'd5,-10'd195};
ram[42344] = {9'd8,-10'd192};
ram[42345] = {9'd11,-10'd189};
ram[42346] = {9'd14,-10'd186};
ram[42347] = {9'd18,-10'd183};
ram[42348] = {9'd21,-10'd180};
ram[42349] = {9'd24,-10'd176};
ram[42350] = {9'd27,-10'd173};
ram[42351] = {9'd30,-10'd170};
ram[42352] = {9'd33,-10'd167};
ram[42353] = {9'd36,-10'd164};
ram[42354] = {9'd40,-10'd161};
ram[42355] = {9'd43,-10'd158};
ram[42356] = {9'd46,-10'd154};
ram[42357] = {9'd49,-10'd151};
ram[42358] = {9'd52,-10'd148};
ram[42359] = {9'd55,-10'd145};
ram[42360] = {9'd58,-10'd142};
ram[42361] = {9'd62,-10'd139};
ram[42362] = {9'd65,-10'd136};
ram[42363] = {9'd68,-10'd132};
ram[42364] = {9'd71,-10'd129};
ram[42365] = {9'd74,-10'd126};
ram[42366] = {9'd77,-10'd123};
ram[42367] = {9'd80,-10'd120};
ram[42368] = {9'd80,-10'd120};
ram[42369] = {9'd84,-10'd117};
ram[42370] = {9'd87,-10'd114};
ram[42371] = {9'd90,-10'd110};
ram[42372] = {9'd93,-10'd107};
ram[42373] = {9'd96,-10'd104};
ram[42374] = {9'd99,-10'd101};
ram[42375] = {-9'd98,-10'd98};
ram[42376] = {-9'd95,-10'd95};
ram[42377] = {-9'd92,-10'd92};
ram[42378] = {-9'd88,-10'd88};
ram[42379] = {-9'd85,-10'd85};
ram[42380] = {-9'd82,-10'd82};
ram[42381] = {-9'd79,-10'd79};
ram[42382] = {-9'd76,-10'd76};
ram[42383] = {-9'd73,-10'd73};
ram[42384] = {-9'd70,-10'd70};
ram[42385] = {-9'd66,-10'd66};
ram[42386] = {-9'd63,-10'd63};
ram[42387] = {-9'd60,-10'd60};
ram[42388] = {-9'd57,-10'd57};
ram[42389] = {-9'd54,-10'd54};
ram[42390] = {-9'd51,-10'd51};
ram[42391] = {-9'd48,-10'd48};
ram[42392] = {-9'd44,-10'd44};
ram[42393] = {-9'd41,-10'd41};
ram[42394] = {-9'd38,-10'd38};
ram[42395] = {-9'd35,-10'd35};
ram[42396] = {-9'd32,-10'd32};
ram[42397] = {-9'd29,-10'd29};
ram[42398] = {-9'd26,-10'd26};
ram[42399] = {-9'd22,-10'd22};
ram[42400] = {-9'd19,-10'd19};
ram[42401] = {-9'd16,-10'd16};
ram[42402] = {-9'd13,-10'd13};
ram[42403] = {-9'd10,-10'd10};
ram[42404] = {-9'd7,-10'd7};
ram[42405] = {-9'd4,-10'd4};
ram[42406] = {9'd0,10'd0};
ram[42407] = {9'd3,10'd3};
ram[42408] = {9'd6,10'd6};
ram[42409] = {9'd9,10'd9};
ram[42410] = {9'd12,10'd12};
ram[42411] = {9'd15,10'd15};
ram[42412] = {9'd18,10'd18};
ram[42413] = {9'd21,10'd21};
ram[42414] = {9'd25,10'd25};
ram[42415] = {9'd28,10'd28};
ram[42416] = {9'd31,10'd31};
ram[42417] = {9'd34,10'd34};
ram[42418] = {9'd37,10'd37};
ram[42419] = {9'd40,10'd40};
ram[42420] = {9'd43,10'd43};
ram[42421] = {9'd47,10'd47};
ram[42422] = {9'd50,10'd50};
ram[42423] = {9'd53,10'd53};
ram[42424] = {9'd56,10'd56};
ram[42425] = {9'd59,10'd59};
ram[42426] = {9'd62,10'd62};
ram[42427] = {9'd65,10'd65};
ram[42428] = {9'd69,10'd69};
ram[42429] = {9'd72,10'd72};
ram[42430] = {9'd75,10'd75};
ram[42431] = {9'd78,10'd78};
ram[42432] = {9'd81,10'd81};
ram[42433] = {9'd84,10'd84};
ram[42434] = {9'd87,10'd87};
ram[42435] = {9'd91,10'd91};
ram[42436] = {9'd94,10'd94};
ram[42437] = {9'd97,10'd97};
ram[42438] = {-9'd100,10'd100};
ram[42439] = {-9'd97,10'd103};
ram[42440] = {-9'd94,10'd106};
ram[42441] = {-9'd91,10'd109};
ram[42442] = {-9'd88,10'd113};
ram[42443] = {-9'd85,10'd116};
ram[42444] = {-9'd81,10'd119};
ram[42445] = {-9'd78,10'd122};
ram[42446] = {-9'd75,10'd125};
ram[42447] = {-9'd72,10'd128};
ram[42448] = {-9'd69,10'd131};
ram[42449] = {-9'd66,10'd135};
ram[42450] = {-9'd63,10'd138};
ram[42451] = {-9'd59,10'd141};
ram[42452] = {-9'd56,10'd144};
ram[42453] = {-9'd53,10'd147};
ram[42454] = {-9'd50,10'd150};
ram[42455] = {-9'd47,10'd153};
ram[42456] = {-9'd44,10'd157};
ram[42457] = {-9'd41,10'd160};
ram[42458] = {-9'd37,10'd163};
ram[42459] = {-9'd34,10'd166};
ram[42460] = {-9'd31,10'd169};
ram[42461] = {-9'd28,10'd172};
ram[42462] = {-9'd25,10'd175};
ram[42463] = {-9'd22,10'd179};
ram[42464] = {-9'd19,10'd182};
ram[42465] = {-9'd15,10'd185};
ram[42466] = {-9'd12,10'd188};
ram[42467] = {-9'd9,10'd191};
ram[42468] = {-9'd6,10'd194};
ram[42469] = {-9'd3,10'd197};
ram[42470] = {9'd0,10'd201};
ram[42471] = {9'd3,10'd204};
ram[42472] = {9'd7,10'd207};
ram[42473] = {9'd10,10'd210};
ram[42474] = {9'd13,10'd213};
ram[42475] = {9'd16,10'd216};
ram[42476] = {9'd19,10'd219};
ram[42477] = {9'd22,10'd223};
ram[42478] = {9'd25,10'd226};
ram[42479] = {9'd29,10'd229};
ram[42480] = {9'd32,10'd232};
ram[42481] = {9'd35,10'd235};
ram[42482] = {9'd38,10'd238};
ram[42483] = {9'd41,10'd241};
ram[42484] = {9'd44,10'd245};
ram[42485] = {9'd47,10'd248};
ram[42486] = {9'd51,10'd251};
ram[42487] = {9'd54,10'd254};
ram[42488] = {9'd57,10'd257};
ram[42489] = {9'd60,10'd260};
ram[42490] = {9'd63,10'd263};
ram[42491] = {9'd66,10'd267};
ram[42492] = {9'd69,10'd270};
ram[42493] = {9'd73,10'd273};
ram[42494] = {9'd76,10'd276};
ram[42495] = {9'd79,10'd279};
ram[42496] = {9'd79,10'd279};
ram[42497] = {9'd82,10'd282};
ram[42498] = {9'd85,10'd285};
ram[42499] = {9'd88,10'd289};
ram[42500] = {9'd91,10'd292};
ram[42501] = {9'd95,10'd295};
ram[42502] = {9'd98,10'd298};
ram[42503] = {-9'd99,10'd301};
ram[42504] = {-9'd96,10'd304};
ram[42505] = {-9'd93,10'd307};
ram[42506] = {-9'd90,10'd311};
ram[42507] = {-9'd87,10'd314};
ram[42508] = {-9'd84,10'd317};
ram[42509] = {-9'd81,10'd320};
ram[42510] = {-9'd77,10'd323};
ram[42511] = {-9'd74,10'd326};
ram[42512] = {-9'd71,10'd329};
ram[42513] = {-9'd68,10'd333};
ram[42514] = {-9'd65,10'd336};
ram[42515] = {-9'd62,10'd339};
ram[42516] = {-9'd59,10'd342};
ram[42517] = {-9'd55,10'd345};
ram[42518] = {-9'd52,10'd348};
ram[42519] = {-9'd49,10'd351};
ram[42520] = {-9'd46,10'd354};
ram[42521] = {-9'd43,10'd358};
ram[42522] = {-9'd40,10'd361};
ram[42523] = {-9'd37,10'd364};
ram[42524] = {-9'd33,10'd367};
ram[42525] = {-9'd30,10'd370};
ram[42526] = {-9'd27,10'd373};
ram[42527] = {-9'd24,10'd376};
ram[42528] = {-9'd21,10'd380};
ram[42529] = {-9'd18,10'd383};
ram[42530] = {-9'd15,10'd386};
ram[42531] = {-9'd11,10'd389};
ram[42532] = {-9'd8,10'd392};
ram[42533] = {-9'd5,10'd395};
ram[42534] = {-9'd2,10'd398};
ram[42535] = {9'd1,-10'd399};
ram[42536] = {9'd4,-10'd396};
ram[42537] = {9'd7,-10'd393};
ram[42538] = {9'd10,-10'd390};
ram[42539] = {9'd14,-10'd387};
ram[42540] = {9'd17,-10'd384};
ram[42541] = {9'd20,-10'd381};
ram[42542] = {9'd23,-10'd377};
ram[42543] = {9'd26,-10'd374};
ram[42544] = {9'd29,-10'd371};
ram[42545] = {9'd32,-10'd368};
ram[42546] = {9'd36,-10'd365};
ram[42547] = {9'd39,-10'd362};
ram[42548] = {9'd42,-10'd359};
ram[42549] = {9'd45,-10'd355};
ram[42550] = {9'd48,-10'd352};
ram[42551] = {9'd51,-10'd349};
ram[42552] = {9'd54,-10'd346};
ram[42553] = {9'd58,-10'd343};
ram[42554] = {9'd61,-10'd340};
ram[42555] = {9'd64,-10'd337};
ram[42556] = {9'd67,-10'd334};
ram[42557] = {9'd70,-10'd330};
ram[42558] = {9'd73,-10'd327};
ram[42559] = {9'd76,-10'd324};
ram[42560] = {9'd80,-10'd321};
ram[42561] = {9'd83,-10'd318};
ram[42562] = {9'd86,-10'd315};
ram[42563] = {9'd89,-10'd312};
ram[42564] = {9'd92,-10'd308};
ram[42565] = {9'd95,-10'd305};
ram[42566] = {9'd98,-10'd302};
ram[42567] = {-9'd99,-10'd299};
ram[42568] = {-9'd96,-10'd296};
ram[42569] = {-9'd92,-10'd293};
ram[42570] = {-9'd89,-10'd290};
ram[42571] = {-9'd86,-10'd286};
ram[42572] = {-9'd83,-10'd283};
ram[42573] = {-9'd80,-10'd280};
ram[42574] = {-9'd77,-10'd277};
ram[42575] = {-9'd74,-10'd274};
ram[42576] = {-9'd70,-10'd271};
ram[42577] = {-9'd67,-10'd268};
ram[42578] = {-9'd64,-10'd264};
ram[42579] = {-9'd61,-10'd261};
ram[42580] = {-9'd58,-10'd258};
ram[42581] = {-9'd55,-10'd255};
ram[42582] = {-9'd52,-10'd252};
ram[42583] = {-9'd48,-10'd249};
ram[42584] = {-9'd45,-10'd246};
ram[42585] = {-9'd42,-10'd242};
ram[42586] = {-9'd39,-10'd239};
ram[42587] = {-9'd36,-10'd236};
ram[42588] = {-9'd33,-10'd233};
ram[42589] = {-9'd30,-10'd230};
ram[42590] = {-9'd26,-10'd227};
ram[42591] = {-9'd23,-10'd224};
ram[42592] = {-9'd20,-10'd220};
ram[42593] = {-9'd17,-10'd217};
ram[42594] = {-9'd14,-10'd214};
ram[42595] = {-9'd11,-10'd211};
ram[42596] = {-9'd8,-10'd208};
ram[42597] = {-9'd4,-10'd205};
ram[42598] = {-9'd1,-10'd202};
ram[42599] = {9'd2,-10'd198};
ram[42600] = {9'd5,-10'd195};
ram[42601] = {9'd8,-10'd192};
ram[42602] = {9'd11,-10'd189};
ram[42603] = {9'd14,-10'd186};
ram[42604] = {9'd18,-10'd183};
ram[42605] = {9'd21,-10'd180};
ram[42606] = {9'd24,-10'd176};
ram[42607] = {9'd27,-10'd173};
ram[42608] = {9'd30,-10'd170};
ram[42609] = {9'd33,-10'd167};
ram[42610] = {9'd36,-10'd164};
ram[42611] = {9'd40,-10'd161};
ram[42612] = {9'd43,-10'd158};
ram[42613] = {9'd46,-10'd154};
ram[42614] = {9'd49,-10'd151};
ram[42615] = {9'd52,-10'd148};
ram[42616] = {9'd55,-10'd145};
ram[42617] = {9'd58,-10'd142};
ram[42618] = {9'd62,-10'd139};
ram[42619] = {9'd65,-10'd136};
ram[42620] = {9'd68,-10'd132};
ram[42621] = {9'd71,-10'd129};
ram[42622] = {9'd74,-10'd126};
ram[42623] = {9'd77,-10'd123};
ram[42624] = {9'd77,-10'd123};
ram[42625] = {9'd80,-10'd120};
ram[42626] = {9'd84,-10'd117};
ram[42627] = {9'd87,-10'd114};
ram[42628] = {9'd90,-10'd110};
ram[42629] = {9'd93,-10'd107};
ram[42630] = {9'd96,-10'd104};
ram[42631] = {9'd99,-10'd101};
ram[42632] = {-9'd98,-10'd98};
ram[42633] = {-9'd95,-10'd95};
ram[42634] = {-9'd92,-10'd92};
ram[42635] = {-9'd88,-10'd88};
ram[42636] = {-9'd85,-10'd85};
ram[42637] = {-9'd82,-10'd82};
ram[42638] = {-9'd79,-10'd79};
ram[42639] = {-9'd76,-10'd76};
ram[42640] = {-9'd73,-10'd73};
ram[42641] = {-9'd70,-10'd70};
ram[42642] = {-9'd66,-10'd66};
ram[42643] = {-9'd63,-10'd63};
ram[42644] = {-9'd60,-10'd60};
ram[42645] = {-9'd57,-10'd57};
ram[42646] = {-9'd54,-10'd54};
ram[42647] = {-9'd51,-10'd51};
ram[42648] = {-9'd48,-10'd48};
ram[42649] = {-9'd44,-10'd44};
ram[42650] = {-9'd41,-10'd41};
ram[42651] = {-9'd38,-10'd38};
ram[42652] = {-9'd35,-10'd35};
ram[42653] = {-9'd32,-10'd32};
ram[42654] = {-9'd29,-10'd29};
ram[42655] = {-9'd26,-10'd26};
ram[42656] = {-9'd22,-10'd22};
ram[42657] = {-9'd19,-10'd19};
ram[42658] = {-9'd16,-10'd16};
ram[42659] = {-9'd13,-10'd13};
ram[42660] = {-9'd10,-10'd10};
ram[42661] = {-9'd7,-10'd7};
ram[42662] = {-9'd4,-10'd4};
ram[42663] = {9'd0,10'd0};
ram[42664] = {9'd3,10'd3};
ram[42665] = {9'd6,10'd6};
ram[42666] = {9'd9,10'd9};
ram[42667] = {9'd12,10'd12};
ram[42668] = {9'd15,10'd15};
ram[42669] = {9'd18,10'd18};
ram[42670] = {9'd21,10'd21};
ram[42671] = {9'd25,10'd25};
ram[42672] = {9'd28,10'd28};
ram[42673] = {9'd31,10'd31};
ram[42674] = {9'd34,10'd34};
ram[42675] = {9'd37,10'd37};
ram[42676] = {9'd40,10'd40};
ram[42677] = {9'd43,10'd43};
ram[42678] = {9'd47,10'd47};
ram[42679] = {9'd50,10'd50};
ram[42680] = {9'd53,10'd53};
ram[42681] = {9'd56,10'd56};
ram[42682] = {9'd59,10'd59};
ram[42683] = {9'd62,10'd62};
ram[42684] = {9'd65,10'd65};
ram[42685] = {9'd69,10'd69};
ram[42686] = {9'd72,10'd72};
ram[42687] = {9'd75,10'd75};
ram[42688] = {9'd78,10'd78};
ram[42689] = {9'd81,10'd81};
ram[42690] = {9'd84,10'd84};
ram[42691] = {9'd87,10'd87};
ram[42692] = {9'd91,10'd91};
ram[42693] = {9'd94,10'd94};
ram[42694] = {9'd97,10'd97};
ram[42695] = {-9'd100,10'd100};
ram[42696] = {-9'd97,10'd103};
ram[42697] = {-9'd94,10'd106};
ram[42698] = {-9'd91,10'd109};
ram[42699] = {-9'd88,10'd113};
ram[42700] = {-9'd85,10'd116};
ram[42701] = {-9'd81,10'd119};
ram[42702] = {-9'd78,10'd122};
ram[42703] = {-9'd75,10'd125};
ram[42704] = {-9'd72,10'd128};
ram[42705] = {-9'd69,10'd131};
ram[42706] = {-9'd66,10'd135};
ram[42707] = {-9'd63,10'd138};
ram[42708] = {-9'd59,10'd141};
ram[42709] = {-9'd56,10'd144};
ram[42710] = {-9'd53,10'd147};
ram[42711] = {-9'd50,10'd150};
ram[42712] = {-9'd47,10'd153};
ram[42713] = {-9'd44,10'd157};
ram[42714] = {-9'd41,10'd160};
ram[42715] = {-9'd37,10'd163};
ram[42716] = {-9'd34,10'd166};
ram[42717] = {-9'd31,10'd169};
ram[42718] = {-9'd28,10'd172};
ram[42719] = {-9'd25,10'd175};
ram[42720] = {-9'd22,10'd179};
ram[42721] = {-9'd19,10'd182};
ram[42722] = {-9'd15,10'd185};
ram[42723] = {-9'd12,10'd188};
ram[42724] = {-9'd9,10'd191};
ram[42725] = {-9'd6,10'd194};
ram[42726] = {-9'd3,10'd197};
ram[42727] = {9'd0,10'd201};
ram[42728] = {9'd3,10'd204};
ram[42729] = {9'd7,10'd207};
ram[42730] = {9'd10,10'd210};
ram[42731] = {9'd13,10'd213};
ram[42732] = {9'd16,10'd216};
ram[42733] = {9'd19,10'd219};
ram[42734] = {9'd22,10'd223};
ram[42735] = {9'd25,10'd226};
ram[42736] = {9'd29,10'd229};
ram[42737] = {9'd32,10'd232};
ram[42738] = {9'd35,10'd235};
ram[42739] = {9'd38,10'd238};
ram[42740] = {9'd41,10'd241};
ram[42741] = {9'd44,10'd245};
ram[42742] = {9'd47,10'd248};
ram[42743] = {9'd51,10'd251};
ram[42744] = {9'd54,10'd254};
ram[42745] = {9'd57,10'd257};
ram[42746] = {9'd60,10'd260};
ram[42747] = {9'd63,10'd263};
ram[42748] = {9'd66,10'd267};
ram[42749] = {9'd69,10'd270};
ram[42750] = {9'd73,10'd273};
ram[42751] = {9'd76,10'd276};
ram[42752] = {9'd76,10'd276};
ram[42753] = {9'd79,10'd279};
ram[42754] = {9'd82,10'd282};
ram[42755] = {9'd85,10'd285};
ram[42756] = {9'd88,10'd289};
ram[42757] = {9'd91,10'd292};
ram[42758] = {9'd95,10'd295};
ram[42759] = {9'd98,10'd298};
ram[42760] = {-9'd99,10'd301};
ram[42761] = {-9'd96,10'd304};
ram[42762] = {-9'd93,10'd307};
ram[42763] = {-9'd90,10'd311};
ram[42764] = {-9'd87,10'd314};
ram[42765] = {-9'd84,10'd317};
ram[42766] = {-9'd81,10'd320};
ram[42767] = {-9'd77,10'd323};
ram[42768] = {-9'd74,10'd326};
ram[42769] = {-9'd71,10'd329};
ram[42770] = {-9'd68,10'd333};
ram[42771] = {-9'd65,10'd336};
ram[42772] = {-9'd62,10'd339};
ram[42773] = {-9'd59,10'd342};
ram[42774] = {-9'd55,10'd345};
ram[42775] = {-9'd52,10'd348};
ram[42776] = {-9'd49,10'd351};
ram[42777] = {-9'd46,10'd354};
ram[42778] = {-9'd43,10'd358};
ram[42779] = {-9'd40,10'd361};
ram[42780] = {-9'd37,10'd364};
ram[42781] = {-9'd33,10'd367};
ram[42782] = {-9'd30,10'd370};
ram[42783] = {-9'd27,10'd373};
ram[42784] = {-9'd24,10'd376};
ram[42785] = {-9'd21,10'd380};
ram[42786] = {-9'd18,10'd383};
ram[42787] = {-9'd15,10'd386};
ram[42788] = {-9'd11,10'd389};
ram[42789] = {-9'd8,10'd392};
ram[42790] = {-9'd5,10'd395};
ram[42791] = {-9'd2,10'd398};
ram[42792] = {9'd1,-10'd399};
ram[42793] = {9'd4,-10'd396};
ram[42794] = {9'd7,-10'd393};
ram[42795] = {9'd10,-10'd390};
ram[42796] = {9'd14,-10'd387};
ram[42797] = {9'd17,-10'd384};
ram[42798] = {9'd20,-10'd381};
ram[42799] = {9'd23,-10'd377};
ram[42800] = {9'd26,-10'd374};
ram[42801] = {9'd29,-10'd371};
ram[42802] = {9'd32,-10'd368};
ram[42803] = {9'd36,-10'd365};
ram[42804] = {9'd39,-10'd362};
ram[42805] = {9'd42,-10'd359};
ram[42806] = {9'd45,-10'd355};
ram[42807] = {9'd48,-10'd352};
ram[42808] = {9'd51,-10'd349};
ram[42809] = {9'd54,-10'd346};
ram[42810] = {9'd58,-10'd343};
ram[42811] = {9'd61,-10'd340};
ram[42812] = {9'd64,-10'd337};
ram[42813] = {9'd67,-10'd334};
ram[42814] = {9'd70,-10'd330};
ram[42815] = {9'd73,-10'd327};
ram[42816] = {9'd76,-10'd324};
ram[42817] = {9'd80,-10'd321};
ram[42818] = {9'd83,-10'd318};
ram[42819] = {9'd86,-10'd315};
ram[42820] = {9'd89,-10'd312};
ram[42821] = {9'd92,-10'd308};
ram[42822] = {9'd95,-10'd305};
ram[42823] = {9'd98,-10'd302};
ram[42824] = {-9'd99,-10'd299};
ram[42825] = {-9'd96,-10'd296};
ram[42826] = {-9'd92,-10'd293};
ram[42827] = {-9'd89,-10'd290};
ram[42828] = {-9'd86,-10'd286};
ram[42829] = {-9'd83,-10'd283};
ram[42830] = {-9'd80,-10'd280};
ram[42831] = {-9'd77,-10'd277};
ram[42832] = {-9'd74,-10'd274};
ram[42833] = {-9'd70,-10'd271};
ram[42834] = {-9'd67,-10'd268};
ram[42835] = {-9'd64,-10'd264};
ram[42836] = {-9'd61,-10'd261};
ram[42837] = {-9'd58,-10'd258};
ram[42838] = {-9'd55,-10'd255};
ram[42839] = {-9'd52,-10'd252};
ram[42840] = {-9'd48,-10'd249};
ram[42841] = {-9'd45,-10'd246};
ram[42842] = {-9'd42,-10'd242};
ram[42843] = {-9'd39,-10'd239};
ram[42844] = {-9'd36,-10'd236};
ram[42845] = {-9'd33,-10'd233};
ram[42846] = {-9'd30,-10'd230};
ram[42847] = {-9'd26,-10'd227};
ram[42848] = {-9'd23,-10'd224};
ram[42849] = {-9'd20,-10'd220};
ram[42850] = {-9'd17,-10'd217};
ram[42851] = {-9'd14,-10'd214};
ram[42852] = {-9'd11,-10'd211};
ram[42853] = {-9'd8,-10'd208};
ram[42854] = {-9'd4,-10'd205};
ram[42855] = {-9'd1,-10'd202};
ram[42856] = {9'd2,-10'd198};
ram[42857] = {9'd5,-10'd195};
ram[42858] = {9'd8,-10'd192};
ram[42859] = {9'd11,-10'd189};
ram[42860] = {9'd14,-10'd186};
ram[42861] = {9'd18,-10'd183};
ram[42862] = {9'd21,-10'd180};
ram[42863] = {9'd24,-10'd176};
ram[42864] = {9'd27,-10'd173};
ram[42865] = {9'd30,-10'd170};
ram[42866] = {9'd33,-10'd167};
ram[42867] = {9'd36,-10'd164};
ram[42868] = {9'd40,-10'd161};
ram[42869] = {9'd43,-10'd158};
ram[42870] = {9'd46,-10'd154};
ram[42871] = {9'd49,-10'd151};
ram[42872] = {9'd52,-10'd148};
ram[42873] = {9'd55,-10'd145};
ram[42874] = {9'd58,-10'd142};
ram[42875] = {9'd62,-10'd139};
ram[42876] = {9'd65,-10'd136};
ram[42877] = {9'd68,-10'd132};
ram[42878] = {9'd71,-10'd129};
ram[42879] = {9'd74,-10'd126};
ram[42880] = {9'd74,-10'd126};
ram[42881] = {9'd77,-10'd123};
ram[42882] = {9'd80,-10'd120};
ram[42883] = {9'd84,-10'd117};
ram[42884] = {9'd87,-10'd114};
ram[42885] = {9'd90,-10'd110};
ram[42886] = {9'd93,-10'd107};
ram[42887] = {9'd96,-10'd104};
ram[42888] = {9'd99,-10'd101};
ram[42889] = {-9'd98,-10'd98};
ram[42890] = {-9'd95,-10'd95};
ram[42891] = {-9'd92,-10'd92};
ram[42892] = {-9'd88,-10'd88};
ram[42893] = {-9'd85,-10'd85};
ram[42894] = {-9'd82,-10'd82};
ram[42895] = {-9'd79,-10'd79};
ram[42896] = {-9'd76,-10'd76};
ram[42897] = {-9'd73,-10'd73};
ram[42898] = {-9'd70,-10'd70};
ram[42899] = {-9'd66,-10'd66};
ram[42900] = {-9'd63,-10'd63};
ram[42901] = {-9'd60,-10'd60};
ram[42902] = {-9'd57,-10'd57};
ram[42903] = {-9'd54,-10'd54};
ram[42904] = {-9'd51,-10'd51};
ram[42905] = {-9'd48,-10'd48};
ram[42906] = {-9'd44,-10'd44};
ram[42907] = {-9'd41,-10'd41};
ram[42908] = {-9'd38,-10'd38};
ram[42909] = {-9'd35,-10'd35};
ram[42910] = {-9'd32,-10'd32};
ram[42911] = {-9'd29,-10'd29};
ram[42912] = {-9'd26,-10'd26};
ram[42913] = {-9'd22,-10'd22};
ram[42914] = {-9'd19,-10'd19};
ram[42915] = {-9'd16,-10'd16};
ram[42916] = {-9'd13,-10'd13};
ram[42917] = {-9'd10,-10'd10};
ram[42918] = {-9'd7,-10'd7};
ram[42919] = {-9'd4,-10'd4};
ram[42920] = {9'd0,10'd0};
ram[42921] = {9'd3,10'd3};
ram[42922] = {9'd6,10'd6};
ram[42923] = {9'd9,10'd9};
ram[42924] = {9'd12,10'd12};
ram[42925] = {9'd15,10'd15};
ram[42926] = {9'd18,10'd18};
ram[42927] = {9'd21,10'd21};
ram[42928] = {9'd25,10'd25};
ram[42929] = {9'd28,10'd28};
ram[42930] = {9'd31,10'd31};
ram[42931] = {9'd34,10'd34};
ram[42932] = {9'd37,10'd37};
ram[42933] = {9'd40,10'd40};
ram[42934] = {9'd43,10'd43};
ram[42935] = {9'd47,10'd47};
ram[42936] = {9'd50,10'd50};
ram[42937] = {9'd53,10'd53};
ram[42938] = {9'd56,10'd56};
ram[42939] = {9'd59,10'd59};
ram[42940] = {9'd62,10'd62};
ram[42941] = {9'd65,10'd65};
ram[42942] = {9'd69,10'd69};
ram[42943] = {9'd72,10'd72};
ram[42944] = {9'd75,10'd75};
ram[42945] = {9'd78,10'd78};
ram[42946] = {9'd81,10'd81};
ram[42947] = {9'd84,10'd84};
ram[42948] = {9'd87,10'd87};
ram[42949] = {9'd91,10'd91};
ram[42950] = {9'd94,10'd94};
ram[42951] = {9'd97,10'd97};
ram[42952] = {-9'd100,10'd100};
ram[42953] = {-9'd97,10'd103};
ram[42954] = {-9'd94,10'd106};
ram[42955] = {-9'd91,10'd109};
ram[42956] = {-9'd88,10'd113};
ram[42957] = {-9'd85,10'd116};
ram[42958] = {-9'd81,10'd119};
ram[42959] = {-9'd78,10'd122};
ram[42960] = {-9'd75,10'd125};
ram[42961] = {-9'd72,10'd128};
ram[42962] = {-9'd69,10'd131};
ram[42963] = {-9'd66,10'd135};
ram[42964] = {-9'd63,10'd138};
ram[42965] = {-9'd59,10'd141};
ram[42966] = {-9'd56,10'd144};
ram[42967] = {-9'd53,10'd147};
ram[42968] = {-9'd50,10'd150};
ram[42969] = {-9'd47,10'd153};
ram[42970] = {-9'd44,10'd157};
ram[42971] = {-9'd41,10'd160};
ram[42972] = {-9'd37,10'd163};
ram[42973] = {-9'd34,10'd166};
ram[42974] = {-9'd31,10'd169};
ram[42975] = {-9'd28,10'd172};
ram[42976] = {-9'd25,10'd175};
ram[42977] = {-9'd22,10'd179};
ram[42978] = {-9'd19,10'd182};
ram[42979] = {-9'd15,10'd185};
ram[42980] = {-9'd12,10'd188};
ram[42981] = {-9'd9,10'd191};
ram[42982] = {-9'd6,10'd194};
ram[42983] = {-9'd3,10'd197};
ram[42984] = {9'd0,10'd201};
ram[42985] = {9'd3,10'd204};
ram[42986] = {9'd7,10'd207};
ram[42987] = {9'd10,10'd210};
ram[42988] = {9'd13,10'd213};
ram[42989] = {9'd16,10'd216};
ram[42990] = {9'd19,10'd219};
ram[42991] = {9'd22,10'd223};
ram[42992] = {9'd25,10'd226};
ram[42993] = {9'd29,10'd229};
ram[42994] = {9'd32,10'd232};
ram[42995] = {9'd35,10'd235};
ram[42996] = {9'd38,10'd238};
ram[42997] = {9'd41,10'd241};
ram[42998] = {9'd44,10'd245};
ram[42999] = {9'd47,10'd248};
ram[43000] = {9'd51,10'd251};
ram[43001] = {9'd54,10'd254};
ram[43002] = {9'd57,10'd257};
ram[43003] = {9'd60,10'd260};
ram[43004] = {9'd63,10'd263};
ram[43005] = {9'd66,10'd267};
ram[43006] = {9'd69,10'd270};
ram[43007] = {9'd73,10'd273};
ram[43008] = {9'd73,10'd273};
ram[43009] = {9'd76,10'd276};
ram[43010] = {9'd79,10'd279};
ram[43011] = {9'd82,10'd282};
ram[43012] = {9'd85,10'd285};
ram[43013] = {9'd88,10'd289};
ram[43014] = {9'd91,10'd292};
ram[43015] = {9'd95,10'd295};
ram[43016] = {9'd98,10'd298};
ram[43017] = {-9'd99,10'd301};
ram[43018] = {-9'd96,10'd304};
ram[43019] = {-9'd93,10'd307};
ram[43020] = {-9'd90,10'd311};
ram[43021] = {-9'd87,10'd314};
ram[43022] = {-9'd84,10'd317};
ram[43023] = {-9'd81,10'd320};
ram[43024] = {-9'd77,10'd323};
ram[43025] = {-9'd74,10'd326};
ram[43026] = {-9'd71,10'd329};
ram[43027] = {-9'd68,10'd333};
ram[43028] = {-9'd65,10'd336};
ram[43029] = {-9'd62,10'd339};
ram[43030] = {-9'd59,10'd342};
ram[43031] = {-9'd55,10'd345};
ram[43032] = {-9'd52,10'd348};
ram[43033] = {-9'd49,10'd351};
ram[43034] = {-9'd46,10'd354};
ram[43035] = {-9'd43,10'd358};
ram[43036] = {-9'd40,10'd361};
ram[43037] = {-9'd37,10'd364};
ram[43038] = {-9'd33,10'd367};
ram[43039] = {-9'd30,10'd370};
ram[43040] = {-9'd27,10'd373};
ram[43041] = {-9'd24,10'd376};
ram[43042] = {-9'd21,10'd380};
ram[43043] = {-9'd18,10'd383};
ram[43044] = {-9'd15,10'd386};
ram[43045] = {-9'd11,10'd389};
ram[43046] = {-9'd8,10'd392};
ram[43047] = {-9'd5,10'd395};
ram[43048] = {-9'd2,10'd398};
ram[43049] = {9'd1,-10'd399};
ram[43050] = {9'd4,-10'd396};
ram[43051] = {9'd7,-10'd393};
ram[43052] = {9'd10,-10'd390};
ram[43053] = {9'd14,-10'd387};
ram[43054] = {9'd17,-10'd384};
ram[43055] = {9'd20,-10'd381};
ram[43056] = {9'd23,-10'd377};
ram[43057] = {9'd26,-10'd374};
ram[43058] = {9'd29,-10'd371};
ram[43059] = {9'd32,-10'd368};
ram[43060] = {9'd36,-10'd365};
ram[43061] = {9'd39,-10'd362};
ram[43062] = {9'd42,-10'd359};
ram[43063] = {9'd45,-10'd355};
ram[43064] = {9'd48,-10'd352};
ram[43065] = {9'd51,-10'd349};
ram[43066] = {9'd54,-10'd346};
ram[43067] = {9'd58,-10'd343};
ram[43068] = {9'd61,-10'd340};
ram[43069] = {9'd64,-10'd337};
ram[43070] = {9'd67,-10'd334};
ram[43071] = {9'd70,-10'd330};
ram[43072] = {9'd73,-10'd327};
ram[43073] = {9'd76,-10'd324};
ram[43074] = {9'd80,-10'd321};
ram[43075] = {9'd83,-10'd318};
ram[43076] = {9'd86,-10'd315};
ram[43077] = {9'd89,-10'd312};
ram[43078] = {9'd92,-10'd308};
ram[43079] = {9'd95,-10'd305};
ram[43080] = {9'd98,-10'd302};
ram[43081] = {-9'd99,-10'd299};
ram[43082] = {-9'd96,-10'd296};
ram[43083] = {-9'd92,-10'd293};
ram[43084] = {-9'd89,-10'd290};
ram[43085] = {-9'd86,-10'd286};
ram[43086] = {-9'd83,-10'd283};
ram[43087] = {-9'd80,-10'd280};
ram[43088] = {-9'd77,-10'd277};
ram[43089] = {-9'd74,-10'd274};
ram[43090] = {-9'd70,-10'd271};
ram[43091] = {-9'd67,-10'd268};
ram[43092] = {-9'd64,-10'd264};
ram[43093] = {-9'd61,-10'd261};
ram[43094] = {-9'd58,-10'd258};
ram[43095] = {-9'd55,-10'd255};
ram[43096] = {-9'd52,-10'd252};
ram[43097] = {-9'd48,-10'd249};
ram[43098] = {-9'd45,-10'd246};
ram[43099] = {-9'd42,-10'd242};
ram[43100] = {-9'd39,-10'd239};
ram[43101] = {-9'd36,-10'd236};
ram[43102] = {-9'd33,-10'd233};
ram[43103] = {-9'd30,-10'd230};
ram[43104] = {-9'd26,-10'd227};
ram[43105] = {-9'd23,-10'd224};
ram[43106] = {-9'd20,-10'd220};
ram[43107] = {-9'd17,-10'd217};
ram[43108] = {-9'd14,-10'd214};
ram[43109] = {-9'd11,-10'd211};
ram[43110] = {-9'd8,-10'd208};
ram[43111] = {-9'd4,-10'd205};
ram[43112] = {-9'd1,-10'd202};
ram[43113] = {9'd2,-10'd198};
ram[43114] = {9'd5,-10'd195};
ram[43115] = {9'd8,-10'd192};
ram[43116] = {9'd11,-10'd189};
ram[43117] = {9'd14,-10'd186};
ram[43118] = {9'd18,-10'd183};
ram[43119] = {9'd21,-10'd180};
ram[43120] = {9'd24,-10'd176};
ram[43121] = {9'd27,-10'd173};
ram[43122] = {9'd30,-10'd170};
ram[43123] = {9'd33,-10'd167};
ram[43124] = {9'd36,-10'd164};
ram[43125] = {9'd40,-10'd161};
ram[43126] = {9'd43,-10'd158};
ram[43127] = {9'd46,-10'd154};
ram[43128] = {9'd49,-10'd151};
ram[43129] = {9'd52,-10'd148};
ram[43130] = {9'd55,-10'd145};
ram[43131] = {9'd58,-10'd142};
ram[43132] = {9'd62,-10'd139};
ram[43133] = {9'd65,-10'd136};
ram[43134] = {9'd68,-10'd132};
ram[43135] = {9'd71,-10'd129};
ram[43136] = {9'd71,-10'd129};
ram[43137] = {9'd74,-10'd126};
ram[43138] = {9'd77,-10'd123};
ram[43139] = {9'd80,-10'd120};
ram[43140] = {9'd84,-10'd117};
ram[43141] = {9'd87,-10'd114};
ram[43142] = {9'd90,-10'd110};
ram[43143] = {9'd93,-10'd107};
ram[43144] = {9'd96,-10'd104};
ram[43145] = {9'd99,-10'd101};
ram[43146] = {-9'd98,-10'd98};
ram[43147] = {-9'd95,-10'd95};
ram[43148] = {-9'd92,-10'd92};
ram[43149] = {-9'd88,-10'd88};
ram[43150] = {-9'd85,-10'd85};
ram[43151] = {-9'd82,-10'd82};
ram[43152] = {-9'd79,-10'd79};
ram[43153] = {-9'd76,-10'd76};
ram[43154] = {-9'd73,-10'd73};
ram[43155] = {-9'd70,-10'd70};
ram[43156] = {-9'd66,-10'd66};
ram[43157] = {-9'd63,-10'd63};
ram[43158] = {-9'd60,-10'd60};
ram[43159] = {-9'd57,-10'd57};
ram[43160] = {-9'd54,-10'd54};
ram[43161] = {-9'd51,-10'd51};
ram[43162] = {-9'd48,-10'd48};
ram[43163] = {-9'd44,-10'd44};
ram[43164] = {-9'd41,-10'd41};
ram[43165] = {-9'd38,-10'd38};
ram[43166] = {-9'd35,-10'd35};
ram[43167] = {-9'd32,-10'd32};
ram[43168] = {-9'd29,-10'd29};
ram[43169] = {-9'd26,-10'd26};
ram[43170] = {-9'd22,-10'd22};
ram[43171] = {-9'd19,-10'd19};
ram[43172] = {-9'd16,-10'd16};
ram[43173] = {-9'd13,-10'd13};
ram[43174] = {-9'd10,-10'd10};
ram[43175] = {-9'd7,-10'd7};
ram[43176] = {-9'd4,-10'd4};
ram[43177] = {9'd0,10'd0};
ram[43178] = {9'd3,10'd3};
ram[43179] = {9'd6,10'd6};
ram[43180] = {9'd9,10'd9};
ram[43181] = {9'd12,10'd12};
ram[43182] = {9'd15,10'd15};
ram[43183] = {9'd18,10'd18};
ram[43184] = {9'd21,10'd21};
ram[43185] = {9'd25,10'd25};
ram[43186] = {9'd28,10'd28};
ram[43187] = {9'd31,10'd31};
ram[43188] = {9'd34,10'd34};
ram[43189] = {9'd37,10'd37};
ram[43190] = {9'd40,10'd40};
ram[43191] = {9'd43,10'd43};
ram[43192] = {9'd47,10'd47};
ram[43193] = {9'd50,10'd50};
ram[43194] = {9'd53,10'd53};
ram[43195] = {9'd56,10'd56};
ram[43196] = {9'd59,10'd59};
ram[43197] = {9'd62,10'd62};
ram[43198] = {9'd65,10'd65};
ram[43199] = {9'd69,10'd69};
ram[43200] = {9'd72,10'd72};
ram[43201] = {9'd75,10'd75};
ram[43202] = {9'd78,10'd78};
ram[43203] = {9'd81,10'd81};
ram[43204] = {9'd84,10'd84};
ram[43205] = {9'd87,10'd87};
ram[43206] = {9'd91,10'd91};
ram[43207] = {9'd94,10'd94};
ram[43208] = {9'd97,10'd97};
ram[43209] = {-9'd100,10'd100};
ram[43210] = {-9'd97,10'd103};
ram[43211] = {-9'd94,10'd106};
ram[43212] = {-9'd91,10'd109};
ram[43213] = {-9'd88,10'd113};
ram[43214] = {-9'd85,10'd116};
ram[43215] = {-9'd81,10'd119};
ram[43216] = {-9'd78,10'd122};
ram[43217] = {-9'd75,10'd125};
ram[43218] = {-9'd72,10'd128};
ram[43219] = {-9'd69,10'd131};
ram[43220] = {-9'd66,10'd135};
ram[43221] = {-9'd63,10'd138};
ram[43222] = {-9'd59,10'd141};
ram[43223] = {-9'd56,10'd144};
ram[43224] = {-9'd53,10'd147};
ram[43225] = {-9'd50,10'd150};
ram[43226] = {-9'd47,10'd153};
ram[43227] = {-9'd44,10'd157};
ram[43228] = {-9'd41,10'd160};
ram[43229] = {-9'd37,10'd163};
ram[43230] = {-9'd34,10'd166};
ram[43231] = {-9'd31,10'd169};
ram[43232] = {-9'd28,10'd172};
ram[43233] = {-9'd25,10'd175};
ram[43234] = {-9'd22,10'd179};
ram[43235] = {-9'd19,10'd182};
ram[43236] = {-9'd15,10'd185};
ram[43237] = {-9'd12,10'd188};
ram[43238] = {-9'd9,10'd191};
ram[43239] = {-9'd6,10'd194};
ram[43240] = {-9'd3,10'd197};
ram[43241] = {9'd0,10'd201};
ram[43242] = {9'd3,10'd204};
ram[43243] = {9'd7,10'd207};
ram[43244] = {9'd10,10'd210};
ram[43245] = {9'd13,10'd213};
ram[43246] = {9'd16,10'd216};
ram[43247] = {9'd19,10'd219};
ram[43248] = {9'd22,10'd223};
ram[43249] = {9'd25,10'd226};
ram[43250] = {9'd29,10'd229};
ram[43251] = {9'd32,10'd232};
ram[43252] = {9'd35,10'd235};
ram[43253] = {9'd38,10'd238};
ram[43254] = {9'd41,10'd241};
ram[43255] = {9'd44,10'd245};
ram[43256] = {9'd47,10'd248};
ram[43257] = {9'd51,10'd251};
ram[43258] = {9'd54,10'd254};
ram[43259] = {9'd57,10'd257};
ram[43260] = {9'd60,10'd260};
ram[43261] = {9'd63,10'd263};
ram[43262] = {9'd66,10'd267};
ram[43263] = {9'd69,10'd270};
ram[43264] = {9'd69,10'd270};
ram[43265] = {9'd73,10'd273};
ram[43266] = {9'd76,10'd276};
ram[43267] = {9'd79,10'd279};
ram[43268] = {9'd82,10'd282};
ram[43269] = {9'd85,10'd285};
ram[43270] = {9'd88,10'd289};
ram[43271] = {9'd91,10'd292};
ram[43272] = {9'd95,10'd295};
ram[43273] = {9'd98,10'd298};
ram[43274] = {-9'd99,10'd301};
ram[43275] = {-9'd96,10'd304};
ram[43276] = {-9'd93,10'd307};
ram[43277] = {-9'd90,10'd311};
ram[43278] = {-9'd87,10'd314};
ram[43279] = {-9'd84,10'd317};
ram[43280] = {-9'd81,10'd320};
ram[43281] = {-9'd77,10'd323};
ram[43282] = {-9'd74,10'd326};
ram[43283] = {-9'd71,10'd329};
ram[43284] = {-9'd68,10'd333};
ram[43285] = {-9'd65,10'd336};
ram[43286] = {-9'd62,10'd339};
ram[43287] = {-9'd59,10'd342};
ram[43288] = {-9'd55,10'd345};
ram[43289] = {-9'd52,10'd348};
ram[43290] = {-9'd49,10'd351};
ram[43291] = {-9'd46,10'd354};
ram[43292] = {-9'd43,10'd358};
ram[43293] = {-9'd40,10'd361};
ram[43294] = {-9'd37,10'd364};
ram[43295] = {-9'd33,10'd367};
ram[43296] = {-9'd30,10'd370};
ram[43297] = {-9'd27,10'd373};
ram[43298] = {-9'd24,10'd376};
ram[43299] = {-9'd21,10'd380};
ram[43300] = {-9'd18,10'd383};
ram[43301] = {-9'd15,10'd386};
ram[43302] = {-9'd11,10'd389};
ram[43303] = {-9'd8,10'd392};
ram[43304] = {-9'd5,10'd395};
ram[43305] = {-9'd2,10'd398};
ram[43306] = {9'd1,-10'd399};
ram[43307] = {9'd4,-10'd396};
ram[43308] = {9'd7,-10'd393};
ram[43309] = {9'd10,-10'd390};
ram[43310] = {9'd14,-10'd387};
ram[43311] = {9'd17,-10'd384};
ram[43312] = {9'd20,-10'd381};
ram[43313] = {9'd23,-10'd377};
ram[43314] = {9'd26,-10'd374};
ram[43315] = {9'd29,-10'd371};
ram[43316] = {9'd32,-10'd368};
ram[43317] = {9'd36,-10'd365};
ram[43318] = {9'd39,-10'd362};
ram[43319] = {9'd42,-10'd359};
ram[43320] = {9'd45,-10'd355};
ram[43321] = {9'd48,-10'd352};
ram[43322] = {9'd51,-10'd349};
ram[43323] = {9'd54,-10'd346};
ram[43324] = {9'd58,-10'd343};
ram[43325] = {9'd61,-10'd340};
ram[43326] = {9'd64,-10'd337};
ram[43327] = {9'd67,-10'd334};
ram[43328] = {9'd70,-10'd330};
ram[43329] = {9'd73,-10'd327};
ram[43330] = {9'd76,-10'd324};
ram[43331] = {9'd80,-10'd321};
ram[43332] = {9'd83,-10'd318};
ram[43333] = {9'd86,-10'd315};
ram[43334] = {9'd89,-10'd312};
ram[43335] = {9'd92,-10'd308};
ram[43336] = {9'd95,-10'd305};
ram[43337] = {9'd98,-10'd302};
ram[43338] = {-9'd99,-10'd299};
ram[43339] = {-9'd96,-10'd296};
ram[43340] = {-9'd92,-10'd293};
ram[43341] = {-9'd89,-10'd290};
ram[43342] = {-9'd86,-10'd286};
ram[43343] = {-9'd83,-10'd283};
ram[43344] = {-9'd80,-10'd280};
ram[43345] = {-9'd77,-10'd277};
ram[43346] = {-9'd74,-10'd274};
ram[43347] = {-9'd70,-10'd271};
ram[43348] = {-9'd67,-10'd268};
ram[43349] = {-9'd64,-10'd264};
ram[43350] = {-9'd61,-10'd261};
ram[43351] = {-9'd58,-10'd258};
ram[43352] = {-9'd55,-10'd255};
ram[43353] = {-9'd52,-10'd252};
ram[43354] = {-9'd48,-10'd249};
ram[43355] = {-9'd45,-10'd246};
ram[43356] = {-9'd42,-10'd242};
ram[43357] = {-9'd39,-10'd239};
ram[43358] = {-9'd36,-10'd236};
ram[43359] = {-9'd33,-10'd233};
ram[43360] = {-9'd30,-10'd230};
ram[43361] = {-9'd26,-10'd227};
ram[43362] = {-9'd23,-10'd224};
ram[43363] = {-9'd20,-10'd220};
ram[43364] = {-9'd17,-10'd217};
ram[43365] = {-9'd14,-10'd214};
ram[43366] = {-9'd11,-10'd211};
ram[43367] = {-9'd8,-10'd208};
ram[43368] = {-9'd4,-10'd205};
ram[43369] = {-9'd1,-10'd202};
ram[43370] = {9'd2,-10'd198};
ram[43371] = {9'd5,-10'd195};
ram[43372] = {9'd8,-10'd192};
ram[43373] = {9'd11,-10'd189};
ram[43374] = {9'd14,-10'd186};
ram[43375] = {9'd18,-10'd183};
ram[43376] = {9'd21,-10'd180};
ram[43377] = {9'd24,-10'd176};
ram[43378] = {9'd27,-10'd173};
ram[43379] = {9'd30,-10'd170};
ram[43380] = {9'd33,-10'd167};
ram[43381] = {9'd36,-10'd164};
ram[43382] = {9'd40,-10'd161};
ram[43383] = {9'd43,-10'd158};
ram[43384] = {9'd46,-10'd154};
ram[43385] = {9'd49,-10'd151};
ram[43386] = {9'd52,-10'd148};
ram[43387] = {9'd55,-10'd145};
ram[43388] = {9'd58,-10'd142};
ram[43389] = {9'd62,-10'd139};
ram[43390] = {9'd65,-10'd136};
ram[43391] = {9'd68,-10'd132};
ram[43392] = {9'd68,-10'd132};
ram[43393] = {9'd71,-10'd129};
ram[43394] = {9'd74,-10'd126};
ram[43395] = {9'd77,-10'd123};
ram[43396] = {9'd80,-10'd120};
ram[43397] = {9'd84,-10'd117};
ram[43398] = {9'd87,-10'd114};
ram[43399] = {9'd90,-10'd110};
ram[43400] = {9'd93,-10'd107};
ram[43401] = {9'd96,-10'd104};
ram[43402] = {9'd99,-10'd101};
ram[43403] = {-9'd98,-10'd98};
ram[43404] = {-9'd95,-10'd95};
ram[43405] = {-9'd92,-10'd92};
ram[43406] = {-9'd88,-10'd88};
ram[43407] = {-9'd85,-10'd85};
ram[43408] = {-9'd82,-10'd82};
ram[43409] = {-9'd79,-10'd79};
ram[43410] = {-9'd76,-10'd76};
ram[43411] = {-9'd73,-10'd73};
ram[43412] = {-9'd70,-10'd70};
ram[43413] = {-9'd66,-10'd66};
ram[43414] = {-9'd63,-10'd63};
ram[43415] = {-9'd60,-10'd60};
ram[43416] = {-9'd57,-10'd57};
ram[43417] = {-9'd54,-10'd54};
ram[43418] = {-9'd51,-10'd51};
ram[43419] = {-9'd48,-10'd48};
ram[43420] = {-9'd44,-10'd44};
ram[43421] = {-9'd41,-10'd41};
ram[43422] = {-9'd38,-10'd38};
ram[43423] = {-9'd35,-10'd35};
ram[43424] = {-9'd32,-10'd32};
ram[43425] = {-9'd29,-10'd29};
ram[43426] = {-9'd26,-10'd26};
ram[43427] = {-9'd22,-10'd22};
ram[43428] = {-9'd19,-10'd19};
ram[43429] = {-9'd16,-10'd16};
ram[43430] = {-9'd13,-10'd13};
ram[43431] = {-9'd10,-10'd10};
ram[43432] = {-9'd7,-10'd7};
ram[43433] = {-9'd4,-10'd4};
ram[43434] = {9'd0,10'd0};
ram[43435] = {9'd3,10'd3};
ram[43436] = {9'd6,10'd6};
ram[43437] = {9'd9,10'd9};
ram[43438] = {9'd12,10'd12};
ram[43439] = {9'd15,10'd15};
ram[43440] = {9'd18,10'd18};
ram[43441] = {9'd21,10'd21};
ram[43442] = {9'd25,10'd25};
ram[43443] = {9'd28,10'd28};
ram[43444] = {9'd31,10'd31};
ram[43445] = {9'd34,10'd34};
ram[43446] = {9'd37,10'd37};
ram[43447] = {9'd40,10'd40};
ram[43448] = {9'd43,10'd43};
ram[43449] = {9'd47,10'd47};
ram[43450] = {9'd50,10'd50};
ram[43451] = {9'd53,10'd53};
ram[43452] = {9'd56,10'd56};
ram[43453] = {9'd59,10'd59};
ram[43454] = {9'd62,10'd62};
ram[43455] = {9'd65,10'd65};
ram[43456] = {9'd69,10'd69};
ram[43457] = {9'd72,10'd72};
ram[43458] = {9'd75,10'd75};
ram[43459] = {9'd78,10'd78};
ram[43460] = {9'd81,10'd81};
ram[43461] = {9'd84,10'd84};
ram[43462] = {9'd87,10'd87};
ram[43463] = {9'd91,10'd91};
ram[43464] = {9'd94,10'd94};
ram[43465] = {9'd97,10'd97};
ram[43466] = {-9'd100,10'd100};
ram[43467] = {-9'd97,10'd103};
ram[43468] = {-9'd94,10'd106};
ram[43469] = {-9'd91,10'd109};
ram[43470] = {-9'd88,10'd113};
ram[43471] = {-9'd85,10'd116};
ram[43472] = {-9'd81,10'd119};
ram[43473] = {-9'd78,10'd122};
ram[43474] = {-9'd75,10'd125};
ram[43475] = {-9'd72,10'd128};
ram[43476] = {-9'd69,10'd131};
ram[43477] = {-9'd66,10'd135};
ram[43478] = {-9'd63,10'd138};
ram[43479] = {-9'd59,10'd141};
ram[43480] = {-9'd56,10'd144};
ram[43481] = {-9'd53,10'd147};
ram[43482] = {-9'd50,10'd150};
ram[43483] = {-9'd47,10'd153};
ram[43484] = {-9'd44,10'd157};
ram[43485] = {-9'd41,10'd160};
ram[43486] = {-9'd37,10'd163};
ram[43487] = {-9'd34,10'd166};
ram[43488] = {-9'd31,10'd169};
ram[43489] = {-9'd28,10'd172};
ram[43490] = {-9'd25,10'd175};
ram[43491] = {-9'd22,10'd179};
ram[43492] = {-9'd19,10'd182};
ram[43493] = {-9'd15,10'd185};
ram[43494] = {-9'd12,10'd188};
ram[43495] = {-9'd9,10'd191};
ram[43496] = {-9'd6,10'd194};
ram[43497] = {-9'd3,10'd197};
ram[43498] = {9'd0,10'd201};
ram[43499] = {9'd3,10'd204};
ram[43500] = {9'd7,10'd207};
ram[43501] = {9'd10,10'd210};
ram[43502] = {9'd13,10'd213};
ram[43503] = {9'd16,10'd216};
ram[43504] = {9'd19,10'd219};
ram[43505] = {9'd22,10'd223};
ram[43506] = {9'd25,10'd226};
ram[43507] = {9'd29,10'd229};
ram[43508] = {9'd32,10'd232};
ram[43509] = {9'd35,10'd235};
ram[43510] = {9'd38,10'd238};
ram[43511] = {9'd41,10'd241};
ram[43512] = {9'd44,10'd245};
ram[43513] = {9'd47,10'd248};
ram[43514] = {9'd51,10'd251};
ram[43515] = {9'd54,10'd254};
ram[43516] = {9'd57,10'd257};
ram[43517] = {9'd60,10'd260};
ram[43518] = {9'd63,10'd263};
ram[43519] = {9'd66,10'd267};
ram[43520] = {9'd66,10'd267};
ram[43521] = {9'd69,10'd270};
ram[43522] = {9'd73,10'd273};
ram[43523] = {9'd76,10'd276};
ram[43524] = {9'd79,10'd279};
ram[43525] = {9'd82,10'd282};
ram[43526] = {9'd85,10'd285};
ram[43527] = {9'd88,10'd289};
ram[43528] = {9'd91,10'd292};
ram[43529] = {9'd95,10'd295};
ram[43530] = {9'd98,10'd298};
ram[43531] = {-9'd99,10'd301};
ram[43532] = {-9'd96,10'd304};
ram[43533] = {-9'd93,10'd307};
ram[43534] = {-9'd90,10'd311};
ram[43535] = {-9'd87,10'd314};
ram[43536] = {-9'd84,10'd317};
ram[43537] = {-9'd81,10'd320};
ram[43538] = {-9'd77,10'd323};
ram[43539] = {-9'd74,10'd326};
ram[43540] = {-9'd71,10'd329};
ram[43541] = {-9'd68,10'd333};
ram[43542] = {-9'd65,10'd336};
ram[43543] = {-9'd62,10'd339};
ram[43544] = {-9'd59,10'd342};
ram[43545] = {-9'd55,10'd345};
ram[43546] = {-9'd52,10'd348};
ram[43547] = {-9'd49,10'd351};
ram[43548] = {-9'd46,10'd354};
ram[43549] = {-9'd43,10'd358};
ram[43550] = {-9'd40,10'd361};
ram[43551] = {-9'd37,10'd364};
ram[43552] = {-9'd33,10'd367};
ram[43553] = {-9'd30,10'd370};
ram[43554] = {-9'd27,10'd373};
ram[43555] = {-9'd24,10'd376};
ram[43556] = {-9'd21,10'd380};
ram[43557] = {-9'd18,10'd383};
ram[43558] = {-9'd15,10'd386};
ram[43559] = {-9'd11,10'd389};
ram[43560] = {-9'd8,10'd392};
ram[43561] = {-9'd5,10'd395};
ram[43562] = {-9'd2,10'd398};
ram[43563] = {9'd1,-10'd399};
ram[43564] = {9'd4,-10'd396};
ram[43565] = {9'd7,-10'd393};
ram[43566] = {9'd10,-10'd390};
ram[43567] = {9'd14,-10'd387};
ram[43568] = {9'd17,-10'd384};
ram[43569] = {9'd20,-10'd381};
ram[43570] = {9'd23,-10'd377};
ram[43571] = {9'd26,-10'd374};
ram[43572] = {9'd29,-10'd371};
ram[43573] = {9'd32,-10'd368};
ram[43574] = {9'd36,-10'd365};
ram[43575] = {9'd39,-10'd362};
ram[43576] = {9'd42,-10'd359};
ram[43577] = {9'd45,-10'd355};
ram[43578] = {9'd48,-10'd352};
ram[43579] = {9'd51,-10'd349};
ram[43580] = {9'd54,-10'd346};
ram[43581] = {9'd58,-10'd343};
ram[43582] = {9'd61,-10'd340};
ram[43583] = {9'd64,-10'd337};
ram[43584] = {9'd67,-10'd334};
ram[43585] = {9'd70,-10'd330};
ram[43586] = {9'd73,-10'd327};
ram[43587] = {9'd76,-10'd324};
ram[43588] = {9'd80,-10'd321};
ram[43589] = {9'd83,-10'd318};
ram[43590] = {9'd86,-10'd315};
ram[43591] = {9'd89,-10'd312};
ram[43592] = {9'd92,-10'd308};
ram[43593] = {9'd95,-10'd305};
ram[43594] = {9'd98,-10'd302};
ram[43595] = {-9'd99,-10'd299};
ram[43596] = {-9'd96,-10'd296};
ram[43597] = {-9'd92,-10'd293};
ram[43598] = {-9'd89,-10'd290};
ram[43599] = {-9'd86,-10'd286};
ram[43600] = {-9'd83,-10'd283};
ram[43601] = {-9'd80,-10'd280};
ram[43602] = {-9'd77,-10'd277};
ram[43603] = {-9'd74,-10'd274};
ram[43604] = {-9'd70,-10'd271};
ram[43605] = {-9'd67,-10'd268};
ram[43606] = {-9'd64,-10'd264};
ram[43607] = {-9'd61,-10'd261};
ram[43608] = {-9'd58,-10'd258};
ram[43609] = {-9'd55,-10'd255};
ram[43610] = {-9'd52,-10'd252};
ram[43611] = {-9'd48,-10'd249};
ram[43612] = {-9'd45,-10'd246};
ram[43613] = {-9'd42,-10'd242};
ram[43614] = {-9'd39,-10'd239};
ram[43615] = {-9'd36,-10'd236};
ram[43616] = {-9'd33,-10'd233};
ram[43617] = {-9'd30,-10'd230};
ram[43618] = {-9'd26,-10'd227};
ram[43619] = {-9'd23,-10'd224};
ram[43620] = {-9'd20,-10'd220};
ram[43621] = {-9'd17,-10'd217};
ram[43622] = {-9'd14,-10'd214};
ram[43623] = {-9'd11,-10'd211};
ram[43624] = {-9'd8,-10'd208};
ram[43625] = {-9'd4,-10'd205};
ram[43626] = {-9'd1,-10'd202};
ram[43627] = {9'd2,-10'd198};
ram[43628] = {9'd5,-10'd195};
ram[43629] = {9'd8,-10'd192};
ram[43630] = {9'd11,-10'd189};
ram[43631] = {9'd14,-10'd186};
ram[43632] = {9'd18,-10'd183};
ram[43633] = {9'd21,-10'd180};
ram[43634] = {9'd24,-10'd176};
ram[43635] = {9'd27,-10'd173};
ram[43636] = {9'd30,-10'd170};
ram[43637] = {9'd33,-10'd167};
ram[43638] = {9'd36,-10'd164};
ram[43639] = {9'd40,-10'd161};
ram[43640] = {9'd43,-10'd158};
ram[43641] = {9'd46,-10'd154};
ram[43642] = {9'd49,-10'd151};
ram[43643] = {9'd52,-10'd148};
ram[43644] = {9'd55,-10'd145};
ram[43645] = {9'd58,-10'd142};
ram[43646] = {9'd62,-10'd139};
ram[43647] = {9'd65,-10'd136};
ram[43648] = {9'd65,-10'd136};
ram[43649] = {9'd68,-10'd132};
ram[43650] = {9'd71,-10'd129};
ram[43651] = {9'd74,-10'd126};
ram[43652] = {9'd77,-10'd123};
ram[43653] = {9'd80,-10'd120};
ram[43654] = {9'd84,-10'd117};
ram[43655] = {9'd87,-10'd114};
ram[43656] = {9'd90,-10'd110};
ram[43657] = {9'd93,-10'd107};
ram[43658] = {9'd96,-10'd104};
ram[43659] = {9'd99,-10'd101};
ram[43660] = {-9'd98,-10'd98};
ram[43661] = {-9'd95,-10'd95};
ram[43662] = {-9'd92,-10'd92};
ram[43663] = {-9'd88,-10'd88};
ram[43664] = {-9'd85,-10'd85};
ram[43665] = {-9'd82,-10'd82};
ram[43666] = {-9'd79,-10'd79};
ram[43667] = {-9'd76,-10'd76};
ram[43668] = {-9'd73,-10'd73};
ram[43669] = {-9'd70,-10'd70};
ram[43670] = {-9'd66,-10'd66};
ram[43671] = {-9'd63,-10'd63};
ram[43672] = {-9'd60,-10'd60};
ram[43673] = {-9'd57,-10'd57};
ram[43674] = {-9'd54,-10'd54};
ram[43675] = {-9'd51,-10'd51};
ram[43676] = {-9'd48,-10'd48};
ram[43677] = {-9'd44,-10'd44};
ram[43678] = {-9'd41,-10'd41};
ram[43679] = {-9'd38,-10'd38};
ram[43680] = {-9'd35,-10'd35};
ram[43681] = {-9'd32,-10'd32};
ram[43682] = {-9'd29,-10'd29};
ram[43683] = {-9'd26,-10'd26};
ram[43684] = {-9'd22,-10'd22};
ram[43685] = {-9'd19,-10'd19};
ram[43686] = {-9'd16,-10'd16};
ram[43687] = {-9'd13,-10'd13};
ram[43688] = {-9'd10,-10'd10};
ram[43689] = {-9'd7,-10'd7};
ram[43690] = {-9'd4,-10'd4};
ram[43691] = {9'd0,10'd0};
ram[43692] = {9'd3,10'd3};
ram[43693] = {9'd6,10'd6};
ram[43694] = {9'd9,10'd9};
ram[43695] = {9'd12,10'd12};
ram[43696] = {9'd15,10'd15};
ram[43697] = {9'd18,10'd18};
ram[43698] = {9'd21,10'd21};
ram[43699] = {9'd25,10'd25};
ram[43700] = {9'd28,10'd28};
ram[43701] = {9'd31,10'd31};
ram[43702] = {9'd34,10'd34};
ram[43703] = {9'd37,10'd37};
ram[43704] = {9'd40,10'd40};
ram[43705] = {9'd43,10'd43};
ram[43706] = {9'd47,10'd47};
ram[43707] = {9'd50,10'd50};
ram[43708] = {9'd53,10'd53};
ram[43709] = {9'd56,10'd56};
ram[43710] = {9'd59,10'd59};
ram[43711] = {9'd62,10'd62};
ram[43712] = {9'd65,10'd65};
ram[43713] = {9'd69,10'd69};
ram[43714] = {9'd72,10'd72};
ram[43715] = {9'd75,10'd75};
ram[43716] = {9'd78,10'd78};
ram[43717] = {9'd81,10'd81};
ram[43718] = {9'd84,10'd84};
ram[43719] = {9'd87,10'd87};
ram[43720] = {9'd91,10'd91};
ram[43721] = {9'd94,10'd94};
ram[43722] = {9'd97,10'd97};
ram[43723] = {-9'd100,10'd100};
ram[43724] = {-9'd97,10'd103};
ram[43725] = {-9'd94,10'd106};
ram[43726] = {-9'd91,10'd109};
ram[43727] = {-9'd88,10'd113};
ram[43728] = {-9'd85,10'd116};
ram[43729] = {-9'd81,10'd119};
ram[43730] = {-9'd78,10'd122};
ram[43731] = {-9'd75,10'd125};
ram[43732] = {-9'd72,10'd128};
ram[43733] = {-9'd69,10'd131};
ram[43734] = {-9'd66,10'd135};
ram[43735] = {-9'd63,10'd138};
ram[43736] = {-9'd59,10'd141};
ram[43737] = {-9'd56,10'd144};
ram[43738] = {-9'd53,10'd147};
ram[43739] = {-9'd50,10'd150};
ram[43740] = {-9'd47,10'd153};
ram[43741] = {-9'd44,10'd157};
ram[43742] = {-9'd41,10'd160};
ram[43743] = {-9'd37,10'd163};
ram[43744] = {-9'd34,10'd166};
ram[43745] = {-9'd31,10'd169};
ram[43746] = {-9'd28,10'd172};
ram[43747] = {-9'd25,10'd175};
ram[43748] = {-9'd22,10'd179};
ram[43749] = {-9'd19,10'd182};
ram[43750] = {-9'd15,10'd185};
ram[43751] = {-9'd12,10'd188};
ram[43752] = {-9'd9,10'd191};
ram[43753] = {-9'd6,10'd194};
ram[43754] = {-9'd3,10'd197};
ram[43755] = {9'd0,10'd201};
ram[43756] = {9'd3,10'd204};
ram[43757] = {9'd7,10'd207};
ram[43758] = {9'd10,10'd210};
ram[43759] = {9'd13,10'd213};
ram[43760] = {9'd16,10'd216};
ram[43761] = {9'd19,10'd219};
ram[43762] = {9'd22,10'd223};
ram[43763] = {9'd25,10'd226};
ram[43764] = {9'd29,10'd229};
ram[43765] = {9'd32,10'd232};
ram[43766] = {9'd35,10'd235};
ram[43767] = {9'd38,10'd238};
ram[43768] = {9'd41,10'd241};
ram[43769] = {9'd44,10'd245};
ram[43770] = {9'd47,10'd248};
ram[43771] = {9'd51,10'd251};
ram[43772] = {9'd54,10'd254};
ram[43773] = {9'd57,10'd257};
ram[43774] = {9'd60,10'd260};
ram[43775] = {9'd63,10'd263};
ram[43776] = {9'd63,10'd263};
ram[43777] = {9'd66,10'd267};
ram[43778] = {9'd69,10'd270};
ram[43779] = {9'd73,10'd273};
ram[43780] = {9'd76,10'd276};
ram[43781] = {9'd79,10'd279};
ram[43782] = {9'd82,10'd282};
ram[43783] = {9'd85,10'd285};
ram[43784] = {9'd88,10'd289};
ram[43785] = {9'd91,10'd292};
ram[43786] = {9'd95,10'd295};
ram[43787] = {9'd98,10'd298};
ram[43788] = {-9'd99,10'd301};
ram[43789] = {-9'd96,10'd304};
ram[43790] = {-9'd93,10'd307};
ram[43791] = {-9'd90,10'd311};
ram[43792] = {-9'd87,10'd314};
ram[43793] = {-9'd84,10'd317};
ram[43794] = {-9'd81,10'd320};
ram[43795] = {-9'd77,10'd323};
ram[43796] = {-9'd74,10'd326};
ram[43797] = {-9'd71,10'd329};
ram[43798] = {-9'd68,10'd333};
ram[43799] = {-9'd65,10'd336};
ram[43800] = {-9'd62,10'd339};
ram[43801] = {-9'd59,10'd342};
ram[43802] = {-9'd55,10'd345};
ram[43803] = {-9'd52,10'd348};
ram[43804] = {-9'd49,10'd351};
ram[43805] = {-9'd46,10'd354};
ram[43806] = {-9'd43,10'd358};
ram[43807] = {-9'd40,10'd361};
ram[43808] = {-9'd37,10'd364};
ram[43809] = {-9'd33,10'd367};
ram[43810] = {-9'd30,10'd370};
ram[43811] = {-9'd27,10'd373};
ram[43812] = {-9'd24,10'd376};
ram[43813] = {-9'd21,10'd380};
ram[43814] = {-9'd18,10'd383};
ram[43815] = {-9'd15,10'd386};
ram[43816] = {-9'd11,10'd389};
ram[43817] = {-9'd8,10'd392};
ram[43818] = {-9'd5,10'd395};
ram[43819] = {-9'd2,10'd398};
ram[43820] = {9'd1,-10'd399};
ram[43821] = {9'd4,-10'd396};
ram[43822] = {9'd7,-10'd393};
ram[43823] = {9'd10,-10'd390};
ram[43824] = {9'd14,-10'd387};
ram[43825] = {9'd17,-10'd384};
ram[43826] = {9'd20,-10'd381};
ram[43827] = {9'd23,-10'd377};
ram[43828] = {9'd26,-10'd374};
ram[43829] = {9'd29,-10'd371};
ram[43830] = {9'd32,-10'd368};
ram[43831] = {9'd36,-10'd365};
ram[43832] = {9'd39,-10'd362};
ram[43833] = {9'd42,-10'd359};
ram[43834] = {9'd45,-10'd355};
ram[43835] = {9'd48,-10'd352};
ram[43836] = {9'd51,-10'd349};
ram[43837] = {9'd54,-10'd346};
ram[43838] = {9'd58,-10'd343};
ram[43839] = {9'd61,-10'd340};
ram[43840] = {9'd64,-10'd337};
ram[43841] = {9'd67,-10'd334};
ram[43842] = {9'd70,-10'd330};
ram[43843] = {9'd73,-10'd327};
ram[43844] = {9'd76,-10'd324};
ram[43845] = {9'd80,-10'd321};
ram[43846] = {9'd83,-10'd318};
ram[43847] = {9'd86,-10'd315};
ram[43848] = {9'd89,-10'd312};
ram[43849] = {9'd92,-10'd308};
ram[43850] = {9'd95,-10'd305};
ram[43851] = {9'd98,-10'd302};
ram[43852] = {-9'd99,-10'd299};
ram[43853] = {-9'd96,-10'd296};
ram[43854] = {-9'd92,-10'd293};
ram[43855] = {-9'd89,-10'd290};
ram[43856] = {-9'd86,-10'd286};
ram[43857] = {-9'd83,-10'd283};
ram[43858] = {-9'd80,-10'd280};
ram[43859] = {-9'd77,-10'd277};
ram[43860] = {-9'd74,-10'd274};
ram[43861] = {-9'd70,-10'd271};
ram[43862] = {-9'd67,-10'd268};
ram[43863] = {-9'd64,-10'd264};
ram[43864] = {-9'd61,-10'd261};
ram[43865] = {-9'd58,-10'd258};
ram[43866] = {-9'd55,-10'd255};
ram[43867] = {-9'd52,-10'd252};
ram[43868] = {-9'd48,-10'd249};
ram[43869] = {-9'd45,-10'd246};
ram[43870] = {-9'd42,-10'd242};
ram[43871] = {-9'd39,-10'd239};
ram[43872] = {-9'd36,-10'd236};
ram[43873] = {-9'd33,-10'd233};
ram[43874] = {-9'd30,-10'd230};
ram[43875] = {-9'd26,-10'd227};
ram[43876] = {-9'd23,-10'd224};
ram[43877] = {-9'd20,-10'd220};
ram[43878] = {-9'd17,-10'd217};
ram[43879] = {-9'd14,-10'd214};
ram[43880] = {-9'd11,-10'd211};
ram[43881] = {-9'd8,-10'd208};
ram[43882] = {-9'd4,-10'd205};
ram[43883] = {-9'd1,-10'd202};
ram[43884] = {9'd2,-10'd198};
ram[43885] = {9'd5,-10'd195};
ram[43886] = {9'd8,-10'd192};
ram[43887] = {9'd11,-10'd189};
ram[43888] = {9'd14,-10'd186};
ram[43889] = {9'd18,-10'd183};
ram[43890] = {9'd21,-10'd180};
ram[43891] = {9'd24,-10'd176};
ram[43892] = {9'd27,-10'd173};
ram[43893] = {9'd30,-10'd170};
ram[43894] = {9'd33,-10'd167};
ram[43895] = {9'd36,-10'd164};
ram[43896] = {9'd40,-10'd161};
ram[43897] = {9'd43,-10'd158};
ram[43898] = {9'd46,-10'd154};
ram[43899] = {9'd49,-10'd151};
ram[43900] = {9'd52,-10'd148};
ram[43901] = {9'd55,-10'd145};
ram[43902] = {9'd58,-10'd142};
ram[43903] = {9'd62,-10'd139};
ram[43904] = {9'd62,-10'd139};
ram[43905] = {9'd65,-10'd136};
ram[43906] = {9'd68,-10'd132};
ram[43907] = {9'd71,-10'd129};
ram[43908] = {9'd74,-10'd126};
ram[43909] = {9'd77,-10'd123};
ram[43910] = {9'd80,-10'd120};
ram[43911] = {9'd84,-10'd117};
ram[43912] = {9'd87,-10'd114};
ram[43913] = {9'd90,-10'd110};
ram[43914] = {9'd93,-10'd107};
ram[43915] = {9'd96,-10'd104};
ram[43916] = {9'd99,-10'd101};
ram[43917] = {-9'd98,-10'd98};
ram[43918] = {-9'd95,-10'd95};
ram[43919] = {-9'd92,-10'd92};
ram[43920] = {-9'd88,-10'd88};
ram[43921] = {-9'd85,-10'd85};
ram[43922] = {-9'd82,-10'd82};
ram[43923] = {-9'd79,-10'd79};
ram[43924] = {-9'd76,-10'd76};
ram[43925] = {-9'd73,-10'd73};
ram[43926] = {-9'd70,-10'd70};
ram[43927] = {-9'd66,-10'd66};
ram[43928] = {-9'd63,-10'd63};
ram[43929] = {-9'd60,-10'd60};
ram[43930] = {-9'd57,-10'd57};
ram[43931] = {-9'd54,-10'd54};
ram[43932] = {-9'd51,-10'd51};
ram[43933] = {-9'd48,-10'd48};
ram[43934] = {-9'd44,-10'd44};
ram[43935] = {-9'd41,-10'd41};
ram[43936] = {-9'd38,-10'd38};
ram[43937] = {-9'd35,-10'd35};
ram[43938] = {-9'd32,-10'd32};
ram[43939] = {-9'd29,-10'd29};
ram[43940] = {-9'd26,-10'd26};
ram[43941] = {-9'd22,-10'd22};
ram[43942] = {-9'd19,-10'd19};
ram[43943] = {-9'd16,-10'd16};
ram[43944] = {-9'd13,-10'd13};
ram[43945] = {-9'd10,-10'd10};
ram[43946] = {-9'd7,-10'd7};
ram[43947] = {-9'd4,-10'd4};
ram[43948] = {9'd0,10'd0};
ram[43949] = {9'd3,10'd3};
ram[43950] = {9'd6,10'd6};
ram[43951] = {9'd9,10'd9};
ram[43952] = {9'd12,10'd12};
ram[43953] = {9'd15,10'd15};
ram[43954] = {9'd18,10'd18};
ram[43955] = {9'd21,10'd21};
ram[43956] = {9'd25,10'd25};
ram[43957] = {9'd28,10'd28};
ram[43958] = {9'd31,10'd31};
ram[43959] = {9'd34,10'd34};
ram[43960] = {9'd37,10'd37};
ram[43961] = {9'd40,10'd40};
ram[43962] = {9'd43,10'd43};
ram[43963] = {9'd47,10'd47};
ram[43964] = {9'd50,10'd50};
ram[43965] = {9'd53,10'd53};
ram[43966] = {9'd56,10'd56};
ram[43967] = {9'd59,10'd59};
ram[43968] = {9'd62,10'd62};
ram[43969] = {9'd65,10'd65};
ram[43970] = {9'd69,10'd69};
ram[43971] = {9'd72,10'd72};
ram[43972] = {9'd75,10'd75};
ram[43973] = {9'd78,10'd78};
ram[43974] = {9'd81,10'd81};
ram[43975] = {9'd84,10'd84};
ram[43976] = {9'd87,10'd87};
ram[43977] = {9'd91,10'd91};
ram[43978] = {9'd94,10'd94};
ram[43979] = {9'd97,10'd97};
ram[43980] = {-9'd100,10'd100};
ram[43981] = {-9'd97,10'd103};
ram[43982] = {-9'd94,10'd106};
ram[43983] = {-9'd91,10'd109};
ram[43984] = {-9'd88,10'd113};
ram[43985] = {-9'd85,10'd116};
ram[43986] = {-9'd81,10'd119};
ram[43987] = {-9'd78,10'd122};
ram[43988] = {-9'd75,10'd125};
ram[43989] = {-9'd72,10'd128};
ram[43990] = {-9'd69,10'd131};
ram[43991] = {-9'd66,10'd135};
ram[43992] = {-9'd63,10'd138};
ram[43993] = {-9'd59,10'd141};
ram[43994] = {-9'd56,10'd144};
ram[43995] = {-9'd53,10'd147};
ram[43996] = {-9'd50,10'd150};
ram[43997] = {-9'd47,10'd153};
ram[43998] = {-9'd44,10'd157};
ram[43999] = {-9'd41,10'd160};
ram[44000] = {-9'd37,10'd163};
ram[44001] = {-9'd34,10'd166};
ram[44002] = {-9'd31,10'd169};
ram[44003] = {-9'd28,10'd172};
ram[44004] = {-9'd25,10'd175};
ram[44005] = {-9'd22,10'd179};
ram[44006] = {-9'd19,10'd182};
ram[44007] = {-9'd15,10'd185};
ram[44008] = {-9'd12,10'd188};
ram[44009] = {-9'd9,10'd191};
ram[44010] = {-9'd6,10'd194};
ram[44011] = {-9'd3,10'd197};
ram[44012] = {9'd0,10'd201};
ram[44013] = {9'd3,10'd204};
ram[44014] = {9'd7,10'd207};
ram[44015] = {9'd10,10'd210};
ram[44016] = {9'd13,10'd213};
ram[44017] = {9'd16,10'd216};
ram[44018] = {9'd19,10'd219};
ram[44019] = {9'd22,10'd223};
ram[44020] = {9'd25,10'd226};
ram[44021] = {9'd29,10'd229};
ram[44022] = {9'd32,10'd232};
ram[44023] = {9'd35,10'd235};
ram[44024] = {9'd38,10'd238};
ram[44025] = {9'd41,10'd241};
ram[44026] = {9'd44,10'd245};
ram[44027] = {9'd47,10'd248};
ram[44028] = {9'd51,10'd251};
ram[44029] = {9'd54,10'd254};
ram[44030] = {9'd57,10'd257};
ram[44031] = {9'd60,10'd260};
ram[44032] = {9'd60,10'd260};
ram[44033] = {9'd63,10'd263};
ram[44034] = {9'd66,10'd267};
ram[44035] = {9'd69,10'd270};
ram[44036] = {9'd73,10'd273};
ram[44037] = {9'd76,10'd276};
ram[44038] = {9'd79,10'd279};
ram[44039] = {9'd82,10'd282};
ram[44040] = {9'd85,10'd285};
ram[44041] = {9'd88,10'd289};
ram[44042] = {9'd91,10'd292};
ram[44043] = {9'd95,10'd295};
ram[44044] = {9'd98,10'd298};
ram[44045] = {-9'd99,10'd301};
ram[44046] = {-9'd96,10'd304};
ram[44047] = {-9'd93,10'd307};
ram[44048] = {-9'd90,10'd311};
ram[44049] = {-9'd87,10'd314};
ram[44050] = {-9'd84,10'd317};
ram[44051] = {-9'd81,10'd320};
ram[44052] = {-9'd77,10'd323};
ram[44053] = {-9'd74,10'd326};
ram[44054] = {-9'd71,10'd329};
ram[44055] = {-9'd68,10'd333};
ram[44056] = {-9'd65,10'd336};
ram[44057] = {-9'd62,10'd339};
ram[44058] = {-9'd59,10'd342};
ram[44059] = {-9'd55,10'd345};
ram[44060] = {-9'd52,10'd348};
ram[44061] = {-9'd49,10'd351};
ram[44062] = {-9'd46,10'd354};
ram[44063] = {-9'd43,10'd358};
ram[44064] = {-9'd40,10'd361};
ram[44065] = {-9'd37,10'd364};
ram[44066] = {-9'd33,10'd367};
ram[44067] = {-9'd30,10'd370};
ram[44068] = {-9'd27,10'd373};
ram[44069] = {-9'd24,10'd376};
ram[44070] = {-9'd21,10'd380};
ram[44071] = {-9'd18,10'd383};
ram[44072] = {-9'd15,10'd386};
ram[44073] = {-9'd11,10'd389};
ram[44074] = {-9'd8,10'd392};
ram[44075] = {-9'd5,10'd395};
ram[44076] = {-9'd2,10'd398};
ram[44077] = {9'd1,-10'd399};
ram[44078] = {9'd4,-10'd396};
ram[44079] = {9'd7,-10'd393};
ram[44080] = {9'd10,-10'd390};
ram[44081] = {9'd14,-10'd387};
ram[44082] = {9'd17,-10'd384};
ram[44083] = {9'd20,-10'd381};
ram[44084] = {9'd23,-10'd377};
ram[44085] = {9'd26,-10'd374};
ram[44086] = {9'd29,-10'd371};
ram[44087] = {9'd32,-10'd368};
ram[44088] = {9'd36,-10'd365};
ram[44089] = {9'd39,-10'd362};
ram[44090] = {9'd42,-10'd359};
ram[44091] = {9'd45,-10'd355};
ram[44092] = {9'd48,-10'd352};
ram[44093] = {9'd51,-10'd349};
ram[44094] = {9'd54,-10'd346};
ram[44095] = {9'd58,-10'd343};
ram[44096] = {9'd61,-10'd340};
ram[44097] = {9'd64,-10'd337};
ram[44098] = {9'd67,-10'd334};
ram[44099] = {9'd70,-10'd330};
ram[44100] = {9'd73,-10'd327};
ram[44101] = {9'd76,-10'd324};
ram[44102] = {9'd80,-10'd321};
ram[44103] = {9'd83,-10'd318};
ram[44104] = {9'd86,-10'd315};
ram[44105] = {9'd89,-10'd312};
ram[44106] = {9'd92,-10'd308};
ram[44107] = {9'd95,-10'd305};
ram[44108] = {9'd98,-10'd302};
ram[44109] = {-9'd99,-10'd299};
ram[44110] = {-9'd96,-10'd296};
ram[44111] = {-9'd92,-10'd293};
ram[44112] = {-9'd89,-10'd290};
ram[44113] = {-9'd86,-10'd286};
ram[44114] = {-9'd83,-10'd283};
ram[44115] = {-9'd80,-10'd280};
ram[44116] = {-9'd77,-10'd277};
ram[44117] = {-9'd74,-10'd274};
ram[44118] = {-9'd70,-10'd271};
ram[44119] = {-9'd67,-10'd268};
ram[44120] = {-9'd64,-10'd264};
ram[44121] = {-9'd61,-10'd261};
ram[44122] = {-9'd58,-10'd258};
ram[44123] = {-9'd55,-10'd255};
ram[44124] = {-9'd52,-10'd252};
ram[44125] = {-9'd48,-10'd249};
ram[44126] = {-9'd45,-10'd246};
ram[44127] = {-9'd42,-10'd242};
ram[44128] = {-9'd39,-10'd239};
ram[44129] = {-9'd36,-10'd236};
ram[44130] = {-9'd33,-10'd233};
ram[44131] = {-9'd30,-10'd230};
ram[44132] = {-9'd26,-10'd227};
ram[44133] = {-9'd23,-10'd224};
ram[44134] = {-9'd20,-10'd220};
ram[44135] = {-9'd17,-10'd217};
ram[44136] = {-9'd14,-10'd214};
ram[44137] = {-9'd11,-10'd211};
ram[44138] = {-9'd8,-10'd208};
ram[44139] = {-9'd4,-10'd205};
ram[44140] = {-9'd1,-10'd202};
ram[44141] = {9'd2,-10'd198};
ram[44142] = {9'd5,-10'd195};
ram[44143] = {9'd8,-10'd192};
ram[44144] = {9'd11,-10'd189};
ram[44145] = {9'd14,-10'd186};
ram[44146] = {9'd18,-10'd183};
ram[44147] = {9'd21,-10'd180};
ram[44148] = {9'd24,-10'd176};
ram[44149] = {9'd27,-10'd173};
ram[44150] = {9'd30,-10'd170};
ram[44151] = {9'd33,-10'd167};
ram[44152] = {9'd36,-10'd164};
ram[44153] = {9'd40,-10'd161};
ram[44154] = {9'd43,-10'd158};
ram[44155] = {9'd46,-10'd154};
ram[44156] = {9'd49,-10'd151};
ram[44157] = {9'd52,-10'd148};
ram[44158] = {9'd55,-10'd145};
ram[44159] = {9'd58,-10'd142};
ram[44160] = {9'd58,-10'd142};
ram[44161] = {9'd62,-10'd139};
ram[44162] = {9'd65,-10'd136};
ram[44163] = {9'd68,-10'd132};
ram[44164] = {9'd71,-10'd129};
ram[44165] = {9'd74,-10'd126};
ram[44166] = {9'd77,-10'd123};
ram[44167] = {9'd80,-10'd120};
ram[44168] = {9'd84,-10'd117};
ram[44169] = {9'd87,-10'd114};
ram[44170] = {9'd90,-10'd110};
ram[44171] = {9'd93,-10'd107};
ram[44172] = {9'd96,-10'd104};
ram[44173] = {9'd99,-10'd101};
ram[44174] = {-9'd98,-10'd98};
ram[44175] = {-9'd95,-10'd95};
ram[44176] = {-9'd92,-10'd92};
ram[44177] = {-9'd88,-10'd88};
ram[44178] = {-9'd85,-10'd85};
ram[44179] = {-9'd82,-10'd82};
ram[44180] = {-9'd79,-10'd79};
ram[44181] = {-9'd76,-10'd76};
ram[44182] = {-9'd73,-10'd73};
ram[44183] = {-9'd70,-10'd70};
ram[44184] = {-9'd66,-10'd66};
ram[44185] = {-9'd63,-10'd63};
ram[44186] = {-9'd60,-10'd60};
ram[44187] = {-9'd57,-10'd57};
ram[44188] = {-9'd54,-10'd54};
ram[44189] = {-9'd51,-10'd51};
ram[44190] = {-9'd48,-10'd48};
ram[44191] = {-9'd44,-10'd44};
ram[44192] = {-9'd41,-10'd41};
ram[44193] = {-9'd38,-10'd38};
ram[44194] = {-9'd35,-10'd35};
ram[44195] = {-9'd32,-10'd32};
ram[44196] = {-9'd29,-10'd29};
ram[44197] = {-9'd26,-10'd26};
ram[44198] = {-9'd22,-10'd22};
ram[44199] = {-9'd19,-10'd19};
ram[44200] = {-9'd16,-10'd16};
ram[44201] = {-9'd13,-10'd13};
ram[44202] = {-9'd10,-10'd10};
ram[44203] = {-9'd7,-10'd7};
ram[44204] = {-9'd4,-10'd4};
ram[44205] = {9'd0,10'd0};
ram[44206] = {9'd3,10'd3};
ram[44207] = {9'd6,10'd6};
ram[44208] = {9'd9,10'd9};
ram[44209] = {9'd12,10'd12};
ram[44210] = {9'd15,10'd15};
ram[44211] = {9'd18,10'd18};
ram[44212] = {9'd21,10'd21};
ram[44213] = {9'd25,10'd25};
ram[44214] = {9'd28,10'd28};
ram[44215] = {9'd31,10'd31};
ram[44216] = {9'd34,10'd34};
ram[44217] = {9'd37,10'd37};
ram[44218] = {9'd40,10'd40};
ram[44219] = {9'd43,10'd43};
ram[44220] = {9'd47,10'd47};
ram[44221] = {9'd50,10'd50};
ram[44222] = {9'd53,10'd53};
ram[44223] = {9'd56,10'd56};
ram[44224] = {9'd59,10'd59};
ram[44225] = {9'd62,10'd62};
ram[44226] = {9'd65,10'd65};
ram[44227] = {9'd69,10'd69};
ram[44228] = {9'd72,10'd72};
ram[44229] = {9'd75,10'd75};
ram[44230] = {9'd78,10'd78};
ram[44231] = {9'd81,10'd81};
ram[44232] = {9'd84,10'd84};
ram[44233] = {9'd87,10'd87};
ram[44234] = {9'd91,10'd91};
ram[44235] = {9'd94,10'd94};
ram[44236] = {9'd97,10'd97};
ram[44237] = {-9'd100,10'd100};
ram[44238] = {-9'd97,10'd103};
ram[44239] = {-9'd94,10'd106};
ram[44240] = {-9'd91,10'd109};
ram[44241] = {-9'd88,10'd113};
ram[44242] = {-9'd85,10'd116};
ram[44243] = {-9'd81,10'd119};
ram[44244] = {-9'd78,10'd122};
ram[44245] = {-9'd75,10'd125};
ram[44246] = {-9'd72,10'd128};
ram[44247] = {-9'd69,10'd131};
ram[44248] = {-9'd66,10'd135};
ram[44249] = {-9'd63,10'd138};
ram[44250] = {-9'd59,10'd141};
ram[44251] = {-9'd56,10'd144};
ram[44252] = {-9'd53,10'd147};
ram[44253] = {-9'd50,10'd150};
ram[44254] = {-9'd47,10'd153};
ram[44255] = {-9'd44,10'd157};
ram[44256] = {-9'd41,10'd160};
ram[44257] = {-9'd37,10'd163};
ram[44258] = {-9'd34,10'd166};
ram[44259] = {-9'd31,10'd169};
ram[44260] = {-9'd28,10'd172};
ram[44261] = {-9'd25,10'd175};
ram[44262] = {-9'd22,10'd179};
ram[44263] = {-9'd19,10'd182};
ram[44264] = {-9'd15,10'd185};
ram[44265] = {-9'd12,10'd188};
ram[44266] = {-9'd9,10'd191};
ram[44267] = {-9'd6,10'd194};
ram[44268] = {-9'd3,10'd197};
ram[44269] = {9'd0,10'd201};
ram[44270] = {9'd3,10'd204};
ram[44271] = {9'd7,10'd207};
ram[44272] = {9'd10,10'd210};
ram[44273] = {9'd13,10'd213};
ram[44274] = {9'd16,10'd216};
ram[44275] = {9'd19,10'd219};
ram[44276] = {9'd22,10'd223};
ram[44277] = {9'd25,10'd226};
ram[44278] = {9'd29,10'd229};
ram[44279] = {9'd32,10'd232};
ram[44280] = {9'd35,10'd235};
ram[44281] = {9'd38,10'd238};
ram[44282] = {9'd41,10'd241};
ram[44283] = {9'd44,10'd245};
ram[44284] = {9'd47,10'd248};
ram[44285] = {9'd51,10'd251};
ram[44286] = {9'd54,10'd254};
ram[44287] = {9'd57,10'd257};
ram[44288] = {9'd57,10'd257};
ram[44289] = {9'd60,10'd260};
ram[44290] = {9'd63,10'd263};
ram[44291] = {9'd66,10'd267};
ram[44292] = {9'd69,10'd270};
ram[44293] = {9'd73,10'd273};
ram[44294] = {9'd76,10'd276};
ram[44295] = {9'd79,10'd279};
ram[44296] = {9'd82,10'd282};
ram[44297] = {9'd85,10'd285};
ram[44298] = {9'd88,10'd289};
ram[44299] = {9'd91,10'd292};
ram[44300] = {9'd95,10'd295};
ram[44301] = {9'd98,10'd298};
ram[44302] = {-9'd99,10'd301};
ram[44303] = {-9'd96,10'd304};
ram[44304] = {-9'd93,10'd307};
ram[44305] = {-9'd90,10'd311};
ram[44306] = {-9'd87,10'd314};
ram[44307] = {-9'd84,10'd317};
ram[44308] = {-9'd81,10'd320};
ram[44309] = {-9'd77,10'd323};
ram[44310] = {-9'd74,10'd326};
ram[44311] = {-9'd71,10'd329};
ram[44312] = {-9'd68,10'd333};
ram[44313] = {-9'd65,10'd336};
ram[44314] = {-9'd62,10'd339};
ram[44315] = {-9'd59,10'd342};
ram[44316] = {-9'd55,10'd345};
ram[44317] = {-9'd52,10'd348};
ram[44318] = {-9'd49,10'd351};
ram[44319] = {-9'd46,10'd354};
ram[44320] = {-9'd43,10'd358};
ram[44321] = {-9'd40,10'd361};
ram[44322] = {-9'd37,10'd364};
ram[44323] = {-9'd33,10'd367};
ram[44324] = {-9'd30,10'd370};
ram[44325] = {-9'd27,10'd373};
ram[44326] = {-9'd24,10'd376};
ram[44327] = {-9'd21,10'd380};
ram[44328] = {-9'd18,10'd383};
ram[44329] = {-9'd15,10'd386};
ram[44330] = {-9'd11,10'd389};
ram[44331] = {-9'd8,10'd392};
ram[44332] = {-9'd5,10'd395};
ram[44333] = {-9'd2,10'd398};
ram[44334] = {9'd1,-10'd399};
ram[44335] = {9'd4,-10'd396};
ram[44336] = {9'd7,-10'd393};
ram[44337] = {9'd10,-10'd390};
ram[44338] = {9'd14,-10'd387};
ram[44339] = {9'd17,-10'd384};
ram[44340] = {9'd20,-10'd381};
ram[44341] = {9'd23,-10'd377};
ram[44342] = {9'd26,-10'd374};
ram[44343] = {9'd29,-10'd371};
ram[44344] = {9'd32,-10'd368};
ram[44345] = {9'd36,-10'd365};
ram[44346] = {9'd39,-10'd362};
ram[44347] = {9'd42,-10'd359};
ram[44348] = {9'd45,-10'd355};
ram[44349] = {9'd48,-10'd352};
ram[44350] = {9'd51,-10'd349};
ram[44351] = {9'd54,-10'd346};
ram[44352] = {9'd58,-10'd343};
ram[44353] = {9'd61,-10'd340};
ram[44354] = {9'd64,-10'd337};
ram[44355] = {9'd67,-10'd334};
ram[44356] = {9'd70,-10'd330};
ram[44357] = {9'd73,-10'd327};
ram[44358] = {9'd76,-10'd324};
ram[44359] = {9'd80,-10'd321};
ram[44360] = {9'd83,-10'd318};
ram[44361] = {9'd86,-10'd315};
ram[44362] = {9'd89,-10'd312};
ram[44363] = {9'd92,-10'd308};
ram[44364] = {9'd95,-10'd305};
ram[44365] = {9'd98,-10'd302};
ram[44366] = {-9'd99,-10'd299};
ram[44367] = {-9'd96,-10'd296};
ram[44368] = {-9'd92,-10'd293};
ram[44369] = {-9'd89,-10'd290};
ram[44370] = {-9'd86,-10'd286};
ram[44371] = {-9'd83,-10'd283};
ram[44372] = {-9'd80,-10'd280};
ram[44373] = {-9'd77,-10'd277};
ram[44374] = {-9'd74,-10'd274};
ram[44375] = {-9'd70,-10'd271};
ram[44376] = {-9'd67,-10'd268};
ram[44377] = {-9'd64,-10'd264};
ram[44378] = {-9'd61,-10'd261};
ram[44379] = {-9'd58,-10'd258};
ram[44380] = {-9'd55,-10'd255};
ram[44381] = {-9'd52,-10'd252};
ram[44382] = {-9'd48,-10'd249};
ram[44383] = {-9'd45,-10'd246};
ram[44384] = {-9'd42,-10'd242};
ram[44385] = {-9'd39,-10'd239};
ram[44386] = {-9'd36,-10'd236};
ram[44387] = {-9'd33,-10'd233};
ram[44388] = {-9'd30,-10'd230};
ram[44389] = {-9'd26,-10'd227};
ram[44390] = {-9'd23,-10'd224};
ram[44391] = {-9'd20,-10'd220};
ram[44392] = {-9'd17,-10'd217};
ram[44393] = {-9'd14,-10'd214};
ram[44394] = {-9'd11,-10'd211};
ram[44395] = {-9'd8,-10'd208};
ram[44396] = {-9'd4,-10'd205};
ram[44397] = {-9'd1,-10'd202};
ram[44398] = {9'd2,-10'd198};
ram[44399] = {9'd5,-10'd195};
ram[44400] = {9'd8,-10'd192};
ram[44401] = {9'd11,-10'd189};
ram[44402] = {9'd14,-10'd186};
ram[44403] = {9'd18,-10'd183};
ram[44404] = {9'd21,-10'd180};
ram[44405] = {9'd24,-10'd176};
ram[44406] = {9'd27,-10'd173};
ram[44407] = {9'd30,-10'd170};
ram[44408] = {9'd33,-10'd167};
ram[44409] = {9'd36,-10'd164};
ram[44410] = {9'd40,-10'd161};
ram[44411] = {9'd43,-10'd158};
ram[44412] = {9'd46,-10'd154};
ram[44413] = {9'd49,-10'd151};
ram[44414] = {9'd52,-10'd148};
ram[44415] = {9'd55,-10'd145};
ram[44416] = {9'd55,-10'd145};
ram[44417] = {9'd58,-10'd142};
ram[44418] = {9'd62,-10'd139};
ram[44419] = {9'd65,-10'd136};
ram[44420] = {9'd68,-10'd132};
ram[44421] = {9'd71,-10'd129};
ram[44422] = {9'd74,-10'd126};
ram[44423] = {9'd77,-10'd123};
ram[44424] = {9'd80,-10'd120};
ram[44425] = {9'd84,-10'd117};
ram[44426] = {9'd87,-10'd114};
ram[44427] = {9'd90,-10'd110};
ram[44428] = {9'd93,-10'd107};
ram[44429] = {9'd96,-10'd104};
ram[44430] = {9'd99,-10'd101};
ram[44431] = {-9'd98,-10'd98};
ram[44432] = {-9'd95,-10'd95};
ram[44433] = {-9'd92,-10'd92};
ram[44434] = {-9'd88,-10'd88};
ram[44435] = {-9'd85,-10'd85};
ram[44436] = {-9'd82,-10'd82};
ram[44437] = {-9'd79,-10'd79};
ram[44438] = {-9'd76,-10'd76};
ram[44439] = {-9'd73,-10'd73};
ram[44440] = {-9'd70,-10'd70};
ram[44441] = {-9'd66,-10'd66};
ram[44442] = {-9'd63,-10'd63};
ram[44443] = {-9'd60,-10'd60};
ram[44444] = {-9'd57,-10'd57};
ram[44445] = {-9'd54,-10'd54};
ram[44446] = {-9'd51,-10'd51};
ram[44447] = {-9'd48,-10'd48};
ram[44448] = {-9'd44,-10'd44};
ram[44449] = {-9'd41,-10'd41};
ram[44450] = {-9'd38,-10'd38};
ram[44451] = {-9'd35,-10'd35};
ram[44452] = {-9'd32,-10'd32};
ram[44453] = {-9'd29,-10'd29};
ram[44454] = {-9'd26,-10'd26};
ram[44455] = {-9'd22,-10'd22};
ram[44456] = {-9'd19,-10'd19};
ram[44457] = {-9'd16,-10'd16};
ram[44458] = {-9'd13,-10'd13};
ram[44459] = {-9'd10,-10'd10};
ram[44460] = {-9'd7,-10'd7};
ram[44461] = {-9'd4,-10'd4};
ram[44462] = {9'd0,10'd0};
ram[44463] = {9'd3,10'd3};
ram[44464] = {9'd6,10'd6};
ram[44465] = {9'd9,10'd9};
ram[44466] = {9'd12,10'd12};
ram[44467] = {9'd15,10'd15};
ram[44468] = {9'd18,10'd18};
ram[44469] = {9'd21,10'd21};
ram[44470] = {9'd25,10'd25};
ram[44471] = {9'd28,10'd28};
ram[44472] = {9'd31,10'd31};
ram[44473] = {9'd34,10'd34};
ram[44474] = {9'd37,10'd37};
ram[44475] = {9'd40,10'd40};
ram[44476] = {9'd43,10'd43};
ram[44477] = {9'd47,10'd47};
ram[44478] = {9'd50,10'd50};
ram[44479] = {9'd53,10'd53};
ram[44480] = {9'd56,10'd56};
ram[44481] = {9'd59,10'd59};
ram[44482] = {9'd62,10'd62};
ram[44483] = {9'd65,10'd65};
ram[44484] = {9'd69,10'd69};
ram[44485] = {9'd72,10'd72};
ram[44486] = {9'd75,10'd75};
ram[44487] = {9'd78,10'd78};
ram[44488] = {9'd81,10'd81};
ram[44489] = {9'd84,10'd84};
ram[44490] = {9'd87,10'd87};
ram[44491] = {9'd91,10'd91};
ram[44492] = {9'd94,10'd94};
ram[44493] = {9'd97,10'd97};
ram[44494] = {-9'd100,10'd100};
ram[44495] = {-9'd97,10'd103};
ram[44496] = {-9'd94,10'd106};
ram[44497] = {-9'd91,10'd109};
ram[44498] = {-9'd88,10'd113};
ram[44499] = {-9'd85,10'd116};
ram[44500] = {-9'd81,10'd119};
ram[44501] = {-9'd78,10'd122};
ram[44502] = {-9'd75,10'd125};
ram[44503] = {-9'd72,10'd128};
ram[44504] = {-9'd69,10'd131};
ram[44505] = {-9'd66,10'd135};
ram[44506] = {-9'd63,10'd138};
ram[44507] = {-9'd59,10'd141};
ram[44508] = {-9'd56,10'd144};
ram[44509] = {-9'd53,10'd147};
ram[44510] = {-9'd50,10'd150};
ram[44511] = {-9'd47,10'd153};
ram[44512] = {-9'd44,10'd157};
ram[44513] = {-9'd41,10'd160};
ram[44514] = {-9'd37,10'd163};
ram[44515] = {-9'd34,10'd166};
ram[44516] = {-9'd31,10'd169};
ram[44517] = {-9'd28,10'd172};
ram[44518] = {-9'd25,10'd175};
ram[44519] = {-9'd22,10'd179};
ram[44520] = {-9'd19,10'd182};
ram[44521] = {-9'd15,10'd185};
ram[44522] = {-9'd12,10'd188};
ram[44523] = {-9'd9,10'd191};
ram[44524] = {-9'd6,10'd194};
ram[44525] = {-9'd3,10'd197};
ram[44526] = {9'd0,10'd201};
ram[44527] = {9'd3,10'd204};
ram[44528] = {9'd7,10'd207};
ram[44529] = {9'd10,10'd210};
ram[44530] = {9'd13,10'd213};
ram[44531] = {9'd16,10'd216};
ram[44532] = {9'd19,10'd219};
ram[44533] = {9'd22,10'd223};
ram[44534] = {9'd25,10'd226};
ram[44535] = {9'd29,10'd229};
ram[44536] = {9'd32,10'd232};
ram[44537] = {9'd35,10'd235};
ram[44538] = {9'd38,10'd238};
ram[44539] = {9'd41,10'd241};
ram[44540] = {9'd44,10'd245};
ram[44541] = {9'd47,10'd248};
ram[44542] = {9'd51,10'd251};
ram[44543] = {9'd54,10'd254};
ram[44544] = {9'd54,10'd254};
ram[44545] = {9'd57,10'd257};
ram[44546] = {9'd60,10'd260};
ram[44547] = {9'd63,10'd263};
ram[44548] = {9'd66,10'd267};
ram[44549] = {9'd69,10'd270};
ram[44550] = {9'd73,10'd273};
ram[44551] = {9'd76,10'd276};
ram[44552] = {9'd79,10'd279};
ram[44553] = {9'd82,10'd282};
ram[44554] = {9'd85,10'd285};
ram[44555] = {9'd88,10'd289};
ram[44556] = {9'd91,10'd292};
ram[44557] = {9'd95,10'd295};
ram[44558] = {9'd98,10'd298};
ram[44559] = {-9'd99,10'd301};
ram[44560] = {-9'd96,10'd304};
ram[44561] = {-9'd93,10'd307};
ram[44562] = {-9'd90,10'd311};
ram[44563] = {-9'd87,10'd314};
ram[44564] = {-9'd84,10'd317};
ram[44565] = {-9'd81,10'd320};
ram[44566] = {-9'd77,10'd323};
ram[44567] = {-9'd74,10'd326};
ram[44568] = {-9'd71,10'd329};
ram[44569] = {-9'd68,10'd333};
ram[44570] = {-9'd65,10'd336};
ram[44571] = {-9'd62,10'd339};
ram[44572] = {-9'd59,10'd342};
ram[44573] = {-9'd55,10'd345};
ram[44574] = {-9'd52,10'd348};
ram[44575] = {-9'd49,10'd351};
ram[44576] = {-9'd46,10'd354};
ram[44577] = {-9'd43,10'd358};
ram[44578] = {-9'd40,10'd361};
ram[44579] = {-9'd37,10'd364};
ram[44580] = {-9'd33,10'd367};
ram[44581] = {-9'd30,10'd370};
ram[44582] = {-9'd27,10'd373};
ram[44583] = {-9'd24,10'd376};
ram[44584] = {-9'd21,10'd380};
ram[44585] = {-9'd18,10'd383};
ram[44586] = {-9'd15,10'd386};
ram[44587] = {-9'd11,10'd389};
ram[44588] = {-9'd8,10'd392};
ram[44589] = {-9'd5,10'd395};
ram[44590] = {-9'd2,10'd398};
ram[44591] = {9'd1,-10'd399};
ram[44592] = {9'd4,-10'd396};
ram[44593] = {9'd7,-10'd393};
ram[44594] = {9'd10,-10'd390};
ram[44595] = {9'd14,-10'd387};
ram[44596] = {9'd17,-10'd384};
ram[44597] = {9'd20,-10'd381};
ram[44598] = {9'd23,-10'd377};
ram[44599] = {9'd26,-10'd374};
ram[44600] = {9'd29,-10'd371};
ram[44601] = {9'd32,-10'd368};
ram[44602] = {9'd36,-10'd365};
ram[44603] = {9'd39,-10'd362};
ram[44604] = {9'd42,-10'd359};
ram[44605] = {9'd45,-10'd355};
ram[44606] = {9'd48,-10'd352};
ram[44607] = {9'd51,-10'd349};
ram[44608] = {9'd54,-10'd346};
ram[44609] = {9'd58,-10'd343};
ram[44610] = {9'd61,-10'd340};
ram[44611] = {9'd64,-10'd337};
ram[44612] = {9'd67,-10'd334};
ram[44613] = {9'd70,-10'd330};
ram[44614] = {9'd73,-10'd327};
ram[44615] = {9'd76,-10'd324};
ram[44616] = {9'd80,-10'd321};
ram[44617] = {9'd83,-10'd318};
ram[44618] = {9'd86,-10'd315};
ram[44619] = {9'd89,-10'd312};
ram[44620] = {9'd92,-10'd308};
ram[44621] = {9'd95,-10'd305};
ram[44622] = {9'd98,-10'd302};
ram[44623] = {-9'd99,-10'd299};
ram[44624] = {-9'd96,-10'd296};
ram[44625] = {-9'd92,-10'd293};
ram[44626] = {-9'd89,-10'd290};
ram[44627] = {-9'd86,-10'd286};
ram[44628] = {-9'd83,-10'd283};
ram[44629] = {-9'd80,-10'd280};
ram[44630] = {-9'd77,-10'd277};
ram[44631] = {-9'd74,-10'd274};
ram[44632] = {-9'd70,-10'd271};
ram[44633] = {-9'd67,-10'd268};
ram[44634] = {-9'd64,-10'd264};
ram[44635] = {-9'd61,-10'd261};
ram[44636] = {-9'd58,-10'd258};
ram[44637] = {-9'd55,-10'd255};
ram[44638] = {-9'd52,-10'd252};
ram[44639] = {-9'd48,-10'd249};
ram[44640] = {-9'd45,-10'd246};
ram[44641] = {-9'd42,-10'd242};
ram[44642] = {-9'd39,-10'd239};
ram[44643] = {-9'd36,-10'd236};
ram[44644] = {-9'd33,-10'd233};
ram[44645] = {-9'd30,-10'd230};
ram[44646] = {-9'd26,-10'd227};
ram[44647] = {-9'd23,-10'd224};
ram[44648] = {-9'd20,-10'd220};
ram[44649] = {-9'd17,-10'd217};
ram[44650] = {-9'd14,-10'd214};
ram[44651] = {-9'd11,-10'd211};
ram[44652] = {-9'd8,-10'd208};
ram[44653] = {-9'd4,-10'd205};
ram[44654] = {-9'd1,-10'd202};
ram[44655] = {9'd2,-10'd198};
ram[44656] = {9'd5,-10'd195};
ram[44657] = {9'd8,-10'd192};
ram[44658] = {9'd11,-10'd189};
ram[44659] = {9'd14,-10'd186};
ram[44660] = {9'd18,-10'd183};
ram[44661] = {9'd21,-10'd180};
ram[44662] = {9'd24,-10'd176};
ram[44663] = {9'd27,-10'd173};
ram[44664] = {9'd30,-10'd170};
ram[44665] = {9'd33,-10'd167};
ram[44666] = {9'd36,-10'd164};
ram[44667] = {9'd40,-10'd161};
ram[44668] = {9'd43,-10'd158};
ram[44669] = {9'd46,-10'd154};
ram[44670] = {9'd49,-10'd151};
ram[44671] = {9'd52,-10'd148};
ram[44672] = {9'd52,-10'd148};
ram[44673] = {9'd55,-10'd145};
ram[44674] = {9'd58,-10'd142};
ram[44675] = {9'd62,-10'd139};
ram[44676] = {9'd65,-10'd136};
ram[44677] = {9'd68,-10'd132};
ram[44678] = {9'd71,-10'd129};
ram[44679] = {9'd74,-10'd126};
ram[44680] = {9'd77,-10'd123};
ram[44681] = {9'd80,-10'd120};
ram[44682] = {9'd84,-10'd117};
ram[44683] = {9'd87,-10'd114};
ram[44684] = {9'd90,-10'd110};
ram[44685] = {9'd93,-10'd107};
ram[44686] = {9'd96,-10'd104};
ram[44687] = {9'd99,-10'd101};
ram[44688] = {-9'd98,-10'd98};
ram[44689] = {-9'd95,-10'd95};
ram[44690] = {-9'd92,-10'd92};
ram[44691] = {-9'd88,-10'd88};
ram[44692] = {-9'd85,-10'd85};
ram[44693] = {-9'd82,-10'd82};
ram[44694] = {-9'd79,-10'd79};
ram[44695] = {-9'd76,-10'd76};
ram[44696] = {-9'd73,-10'd73};
ram[44697] = {-9'd70,-10'd70};
ram[44698] = {-9'd66,-10'd66};
ram[44699] = {-9'd63,-10'd63};
ram[44700] = {-9'd60,-10'd60};
ram[44701] = {-9'd57,-10'd57};
ram[44702] = {-9'd54,-10'd54};
ram[44703] = {-9'd51,-10'd51};
ram[44704] = {-9'd48,-10'd48};
ram[44705] = {-9'd44,-10'd44};
ram[44706] = {-9'd41,-10'd41};
ram[44707] = {-9'd38,-10'd38};
ram[44708] = {-9'd35,-10'd35};
ram[44709] = {-9'd32,-10'd32};
ram[44710] = {-9'd29,-10'd29};
ram[44711] = {-9'd26,-10'd26};
ram[44712] = {-9'd22,-10'd22};
ram[44713] = {-9'd19,-10'd19};
ram[44714] = {-9'd16,-10'd16};
ram[44715] = {-9'd13,-10'd13};
ram[44716] = {-9'd10,-10'd10};
ram[44717] = {-9'd7,-10'd7};
ram[44718] = {-9'd4,-10'd4};
ram[44719] = {9'd0,10'd0};
ram[44720] = {9'd3,10'd3};
ram[44721] = {9'd6,10'd6};
ram[44722] = {9'd9,10'd9};
ram[44723] = {9'd12,10'd12};
ram[44724] = {9'd15,10'd15};
ram[44725] = {9'd18,10'd18};
ram[44726] = {9'd21,10'd21};
ram[44727] = {9'd25,10'd25};
ram[44728] = {9'd28,10'd28};
ram[44729] = {9'd31,10'd31};
ram[44730] = {9'd34,10'd34};
ram[44731] = {9'd37,10'd37};
ram[44732] = {9'd40,10'd40};
ram[44733] = {9'd43,10'd43};
ram[44734] = {9'd47,10'd47};
ram[44735] = {9'd50,10'd50};
ram[44736] = {9'd53,10'd53};
ram[44737] = {9'd56,10'd56};
ram[44738] = {9'd59,10'd59};
ram[44739] = {9'd62,10'd62};
ram[44740] = {9'd65,10'd65};
ram[44741] = {9'd69,10'd69};
ram[44742] = {9'd72,10'd72};
ram[44743] = {9'd75,10'd75};
ram[44744] = {9'd78,10'd78};
ram[44745] = {9'd81,10'd81};
ram[44746] = {9'd84,10'd84};
ram[44747] = {9'd87,10'd87};
ram[44748] = {9'd91,10'd91};
ram[44749] = {9'd94,10'd94};
ram[44750] = {9'd97,10'd97};
ram[44751] = {-9'd100,10'd100};
ram[44752] = {-9'd97,10'd103};
ram[44753] = {-9'd94,10'd106};
ram[44754] = {-9'd91,10'd109};
ram[44755] = {-9'd88,10'd113};
ram[44756] = {-9'd85,10'd116};
ram[44757] = {-9'd81,10'd119};
ram[44758] = {-9'd78,10'd122};
ram[44759] = {-9'd75,10'd125};
ram[44760] = {-9'd72,10'd128};
ram[44761] = {-9'd69,10'd131};
ram[44762] = {-9'd66,10'd135};
ram[44763] = {-9'd63,10'd138};
ram[44764] = {-9'd59,10'd141};
ram[44765] = {-9'd56,10'd144};
ram[44766] = {-9'd53,10'd147};
ram[44767] = {-9'd50,10'd150};
ram[44768] = {-9'd47,10'd153};
ram[44769] = {-9'd44,10'd157};
ram[44770] = {-9'd41,10'd160};
ram[44771] = {-9'd37,10'd163};
ram[44772] = {-9'd34,10'd166};
ram[44773] = {-9'd31,10'd169};
ram[44774] = {-9'd28,10'd172};
ram[44775] = {-9'd25,10'd175};
ram[44776] = {-9'd22,10'd179};
ram[44777] = {-9'd19,10'd182};
ram[44778] = {-9'd15,10'd185};
ram[44779] = {-9'd12,10'd188};
ram[44780] = {-9'd9,10'd191};
ram[44781] = {-9'd6,10'd194};
ram[44782] = {-9'd3,10'd197};
ram[44783] = {9'd0,10'd201};
ram[44784] = {9'd3,10'd204};
ram[44785] = {9'd7,10'd207};
ram[44786] = {9'd10,10'd210};
ram[44787] = {9'd13,10'd213};
ram[44788] = {9'd16,10'd216};
ram[44789] = {9'd19,10'd219};
ram[44790] = {9'd22,10'd223};
ram[44791] = {9'd25,10'd226};
ram[44792] = {9'd29,10'd229};
ram[44793] = {9'd32,10'd232};
ram[44794] = {9'd35,10'd235};
ram[44795] = {9'd38,10'd238};
ram[44796] = {9'd41,10'd241};
ram[44797] = {9'd44,10'd245};
ram[44798] = {9'd47,10'd248};
ram[44799] = {9'd51,10'd251};
ram[44800] = {9'd51,10'd251};
ram[44801] = {9'd54,10'd254};
ram[44802] = {9'd57,10'd257};
ram[44803] = {9'd60,10'd260};
ram[44804] = {9'd63,10'd263};
ram[44805] = {9'd66,10'd267};
ram[44806] = {9'd69,10'd270};
ram[44807] = {9'd73,10'd273};
ram[44808] = {9'd76,10'd276};
ram[44809] = {9'd79,10'd279};
ram[44810] = {9'd82,10'd282};
ram[44811] = {9'd85,10'd285};
ram[44812] = {9'd88,10'd289};
ram[44813] = {9'd91,10'd292};
ram[44814] = {9'd95,10'd295};
ram[44815] = {9'd98,10'd298};
ram[44816] = {-9'd99,10'd301};
ram[44817] = {-9'd96,10'd304};
ram[44818] = {-9'd93,10'd307};
ram[44819] = {-9'd90,10'd311};
ram[44820] = {-9'd87,10'd314};
ram[44821] = {-9'd84,10'd317};
ram[44822] = {-9'd81,10'd320};
ram[44823] = {-9'd77,10'd323};
ram[44824] = {-9'd74,10'd326};
ram[44825] = {-9'd71,10'd329};
ram[44826] = {-9'd68,10'd333};
ram[44827] = {-9'd65,10'd336};
ram[44828] = {-9'd62,10'd339};
ram[44829] = {-9'd59,10'd342};
ram[44830] = {-9'd55,10'd345};
ram[44831] = {-9'd52,10'd348};
ram[44832] = {-9'd49,10'd351};
ram[44833] = {-9'd46,10'd354};
ram[44834] = {-9'd43,10'd358};
ram[44835] = {-9'd40,10'd361};
ram[44836] = {-9'd37,10'd364};
ram[44837] = {-9'd33,10'd367};
ram[44838] = {-9'd30,10'd370};
ram[44839] = {-9'd27,10'd373};
ram[44840] = {-9'd24,10'd376};
ram[44841] = {-9'd21,10'd380};
ram[44842] = {-9'd18,10'd383};
ram[44843] = {-9'd15,10'd386};
ram[44844] = {-9'd11,10'd389};
ram[44845] = {-9'd8,10'd392};
ram[44846] = {-9'd5,10'd395};
ram[44847] = {-9'd2,10'd398};
ram[44848] = {9'd1,-10'd399};
ram[44849] = {9'd4,-10'd396};
ram[44850] = {9'd7,-10'd393};
ram[44851] = {9'd10,-10'd390};
ram[44852] = {9'd14,-10'd387};
ram[44853] = {9'd17,-10'd384};
ram[44854] = {9'd20,-10'd381};
ram[44855] = {9'd23,-10'd377};
ram[44856] = {9'd26,-10'd374};
ram[44857] = {9'd29,-10'd371};
ram[44858] = {9'd32,-10'd368};
ram[44859] = {9'd36,-10'd365};
ram[44860] = {9'd39,-10'd362};
ram[44861] = {9'd42,-10'd359};
ram[44862] = {9'd45,-10'd355};
ram[44863] = {9'd48,-10'd352};
ram[44864] = {9'd51,-10'd349};
ram[44865] = {9'd54,-10'd346};
ram[44866] = {9'd58,-10'd343};
ram[44867] = {9'd61,-10'd340};
ram[44868] = {9'd64,-10'd337};
ram[44869] = {9'd67,-10'd334};
ram[44870] = {9'd70,-10'd330};
ram[44871] = {9'd73,-10'd327};
ram[44872] = {9'd76,-10'd324};
ram[44873] = {9'd80,-10'd321};
ram[44874] = {9'd83,-10'd318};
ram[44875] = {9'd86,-10'd315};
ram[44876] = {9'd89,-10'd312};
ram[44877] = {9'd92,-10'd308};
ram[44878] = {9'd95,-10'd305};
ram[44879] = {9'd98,-10'd302};
ram[44880] = {-9'd99,-10'd299};
ram[44881] = {-9'd96,-10'd296};
ram[44882] = {-9'd92,-10'd293};
ram[44883] = {-9'd89,-10'd290};
ram[44884] = {-9'd86,-10'd286};
ram[44885] = {-9'd83,-10'd283};
ram[44886] = {-9'd80,-10'd280};
ram[44887] = {-9'd77,-10'd277};
ram[44888] = {-9'd74,-10'd274};
ram[44889] = {-9'd70,-10'd271};
ram[44890] = {-9'd67,-10'd268};
ram[44891] = {-9'd64,-10'd264};
ram[44892] = {-9'd61,-10'd261};
ram[44893] = {-9'd58,-10'd258};
ram[44894] = {-9'd55,-10'd255};
ram[44895] = {-9'd52,-10'd252};
ram[44896] = {-9'd48,-10'd249};
ram[44897] = {-9'd45,-10'd246};
ram[44898] = {-9'd42,-10'd242};
ram[44899] = {-9'd39,-10'd239};
ram[44900] = {-9'd36,-10'd236};
ram[44901] = {-9'd33,-10'd233};
ram[44902] = {-9'd30,-10'd230};
ram[44903] = {-9'd26,-10'd227};
ram[44904] = {-9'd23,-10'd224};
ram[44905] = {-9'd20,-10'd220};
ram[44906] = {-9'd17,-10'd217};
ram[44907] = {-9'd14,-10'd214};
ram[44908] = {-9'd11,-10'd211};
ram[44909] = {-9'd8,-10'd208};
ram[44910] = {-9'd4,-10'd205};
ram[44911] = {-9'd1,-10'd202};
ram[44912] = {9'd2,-10'd198};
ram[44913] = {9'd5,-10'd195};
ram[44914] = {9'd8,-10'd192};
ram[44915] = {9'd11,-10'd189};
ram[44916] = {9'd14,-10'd186};
ram[44917] = {9'd18,-10'd183};
ram[44918] = {9'd21,-10'd180};
ram[44919] = {9'd24,-10'd176};
ram[44920] = {9'd27,-10'd173};
ram[44921] = {9'd30,-10'd170};
ram[44922] = {9'd33,-10'd167};
ram[44923] = {9'd36,-10'd164};
ram[44924] = {9'd40,-10'd161};
ram[44925] = {9'd43,-10'd158};
ram[44926] = {9'd46,-10'd154};
ram[44927] = {9'd49,-10'd151};
ram[44928] = {9'd49,-10'd151};
ram[44929] = {9'd52,-10'd148};
ram[44930] = {9'd55,-10'd145};
ram[44931] = {9'd58,-10'd142};
ram[44932] = {9'd62,-10'd139};
ram[44933] = {9'd65,-10'd136};
ram[44934] = {9'd68,-10'd132};
ram[44935] = {9'd71,-10'd129};
ram[44936] = {9'd74,-10'd126};
ram[44937] = {9'd77,-10'd123};
ram[44938] = {9'd80,-10'd120};
ram[44939] = {9'd84,-10'd117};
ram[44940] = {9'd87,-10'd114};
ram[44941] = {9'd90,-10'd110};
ram[44942] = {9'd93,-10'd107};
ram[44943] = {9'd96,-10'd104};
ram[44944] = {9'd99,-10'd101};
ram[44945] = {-9'd98,-10'd98};
ram[44946] = {-9'd95,-10'd95};
ram[44947] = {-9'd92,-10'd92};
ram[44948] = {-9'd88,-10'd88};
ram[44949] = {-9'd85,-10'd85};
ram[44950] = {-9'd82,-10'd82};
ram[44951] = {-9'd79,-10'd79};
ram[44952] = {-9'd76,-10'd76};
ram[44953] = {-9'd73,-10'd73};
ram[44954] = {-9'd70,-10'd70};
ram[44955] = {-9'd66,-10'd66};
ram[44956] = {-9'd63,-10'd63};
ram[44957] = {-9'd60,-10'd60};
ram[44958] = {-9'd57,-10'd57};
ram[44959] = {-9'd54,-10'd54};
ram[44960] = {-9'd51,-10'd51};
ram[44961] = {-9'd48,-10'd48};
ram[44962] = {-9'd44,-10'd44};
ram[44963] = {-9'd41,-10'd41};
ram[44964] = {-9'd38,-10'd38};
ram[44965] = {-9'd35,-10'd35};
ram[44966] = {-9'd32,-10'd32};
ram[44967] = {-9'd29,-10'd29};
ram[44968] = {-9'd26,-10'd26};
ram[44969] = {-9'd22,-10'd22};
ram[44970] = {-9'd19,-10'd19};
ram[44971] = {-9'd16,-10'd16};
ram[44972] = {-9'd13,-10'd13};
ram[44973] = {-9'd10,-10'd10};
ram[44974] = {-9'd7,-10'd7};
ram[44975] = {-9'd4,-10'd4};
ram[44976] = {9'd0,10'd0};
ram[44977] = {9'd3,10'd3};
ram[44978] = {9'd6,10'd6};
ram[44979] = {9'd9,10'd9};
ram[44980] = {9'd12,10'd12};
ram[44981] = {9'd15,10'd15};
ram[44982] = {9'd18,10'd18};
ram[44983] = {9'd21,10'd21};
ram[44984] = {9'd25,10'd25};
ram[44985] = {9'd28,10'd28};
ram[44986] = {9'd31,10'd31};
ram[44987] = {9'd34,10'd34};
ram[44988] = {9'd37,10'd37};
ram[44989] = {9'd40,10'd40};
ram[44990] = {9'd43,10'd43};
ram[44991] = {9'd47,10'd47};
ram[44992] = {9'd50,10'd50};
ram[44993] = {9'd53,10'd53};
ram[44994] = {9'd56,10'd56};
ram[44995] = {9'd59,10'd59};
ram[44996] = {9'd62,10'd62};
ram[44997] = {9'd65,10'd65};
ram[44998] = {9'd69,10'd69};
ram[44999] = {9'd72,10'd72};
ram[45000] = {9'd75,10'd75};
ram[45001] = {9'd78,10'd78};
ram[45002] = {9'd81,10'd81};
ram[45003] = {9'd84,10'd84};
ram[45004] = {9'd87,10'd87};
ram[45005] = {9'd91,10'd91};
ram[45006] = {9'd94,10'd94};
ram[45007] = {9'd97,10'd97};
ram[45008] = {-9'd100,10'd100};
ram[45009] = {-9'd97,10'd103};
ram[45010] = {-9'd94,10'd106};
ram[45011] = {-9'd91,10'd109};
ram[45012] = {-9'd88,10'd113};
ram[45013] = {-9'd85,10'd116};
ram[45014] = {-9'd81,10'd119};
ram[45015] = {-9'd78,10'd122};
ram[45016] = {-9'd75,10'd125};
ram[45017] = {-9'd72,10'd128};
ram[45018] = {-9'd69,10'd131};
ram[45019] = {-9'd66,10'd135};
ram[45020] = {-9'd63,10'd138};
ram[45021] = {-9'd59,10'd141};
ram[45022] = {-9'd56,10'd144};
ram[45023] = {-9'd53,10'd147};
ram[45024] = {-9'd50,10'd150};
ram[45025] = {-9'd47,10'd153};
ram[45026] = {-9'd44,10'd157};
ram[45027] = {-9'd41,10'd160};
ram[45028] = {-9'd37,10'd163};
ram[45029] = {-9'd34,10'd166};
ram[45030] = {-9'd31,10'd169};
ram[45031] = {-9'd28,10'd172};
ram[45032] = {-9'd25,10'd175};
ram[45033] = {-9'd22,10'd179};
ram[45034] = {-9'd19,10'd182};
ram[45035] = {-9'd15,10'd185};
ram[45036] = {-9'd12,10'd188};
ram[45037] = {-9'd9,10'd191};
ram[45038] = {-9'd6,10'd194};
ram[45039] = {-9'd3,10'd197};
ram[45040] = {9'd0,10'd201};
ram[45041] = {9'd3,10'd204};
ram[45042] = {9'd7,10'd207};
ram[45043] = {9'd10,10'd210};
ram[45044] = {9'd13,10'd213};
ram[45045] = {9'd16,10'd216};
ram[45046] = {9'd19,10'd219};
ram[45047] = {9'd22,10'd223};
ram[45048] = {9'd25,10'd226};
ram[45049] = {9'd29,10'd229};
ram[45050] = {9'd32,10'd232};
ram[45051] = {9'd35,10'd235};
ram[45052] = {9'd38,10'd238};
ram[45053] = {9'd41,10'd241};
ram[45054] = {9'd44,10'd245};
ram[45055] = {9'd47,10'd248};
ram[45056] = {9'd47,10'd248};
ram[45057] = {9'd51,10'd251};
ram[45058] = {9'd54,10'd254};
ram[45059] = {9'd57,10'd257};
ram[45060] = {9'd60,10'd260};
ram[45061] = {9'd63,10'd263};
ram[45062] = {9'd66,10'd267};
ram[45063] = {9'd69,10'd270};
ram[45064] = {9'd73,10'd273};
ram[45065] = {9'd76,10'd276};
ram[45066] = {9'd79,10'd279};
ram[45067] = {9'd82,10'd282};
ram[45068] = {9'd85,10'd285};
ram[45069] = {9'd88,10'd289};
ram[45070] = {9'd91,10'd292};
ram[45071] = {9'd95,10'd295};
ram[45072] = {9'd98,10'd298};
ram[45073] = {-9'd99,10'd301};
ram[45074] = {-9'd96,10'd304};
ram[45075] = {-9'd93,10'd307};
ram[45076] = {-9'd90,10'd311};
ram[45077] = {-9'd87,10'd314};
ram[45078] = {-9'd84,10'd317};
ram[45079] = {-9'd81,10'd320};
ram[45080] = {-9'd77,10'd323};
ram[45081] = {-9'd74,10'd326};
ram[45082] = {-9'd71,10'd329};
ram[45083] = {-9'd68,10'd333};
ram[45084] = {-9'd65,10'd336};
ram[45085] = {-9'd62,10'd339};
ram[45086] = {-9'd59,10'd342};
ram[45087] = {-9'd55,10'd345};
ram[45088] = {-9'd52,10'd348};
ram[45089] = {-9'd49,10'd351};
ram[45090] = {-9'd46,10'd354};
ram[45091] = {-9'd43,10'd358};
ram[45092] = {-9'd40,10'd361};
ram[45093] = {-9'd37,10'd364};
ram[45094] = {-9'd33,10'd367};
ram[45095] = {-9'd30,10'd370};
ram[45096] = {-9'd27,10'd373};
ram[45097] = {-9'd24,10'd376};
ram[45098] = {-9'd21,10'd380};
ram[45099] = {-9'd18,10'd383};
ram[45100] = {-9'd15,10'd386};
ram[45101] = {-9'd11,10'd389};
ram[45102] = {-9'd8,10'd392};
ram[45103] = {-9'd5,10'd395};
ram[45104] = {-9'd2,10'd398};
ram[45105] = {9'd1,-10'd399};
ram[45106] = {9'd4,-10'd396};
ram[45107] = {9'd7,-10'd393};
ram[45108] = {9'd10,-10'd390};
ram[45109] = {9'd14,-10'd387};
ram[45110] = {9'd17,-10'd384};
ram[45111] = {9'd20,-10'd381};
ram[45112] = {9'd23,-10'd377};
ram[45113] = {9'd26,-10'd374};
ram[45114] = {9'd29,-10'd371};
ram[45115] = {9'd32,-10'd368};
ram[45116] = {9'd36,-10'd365};
ram[45117] = {9'd39,-10'd362};
ram[45118] = {9'd42,-10'd359};
ram[45119] = {9'd45,-10'd355};
ram[45120] = {9'd48,-10'd352};
ram[45121] = {9'd51,-10'd349};
ram[45122] = {9'd54,-10'd346};
ram[45123] = {9'd58,-10'd343};
ram[45124] = {9'd61,-10'd340};
ram[45125] = {9'd64,-10'd337};
ram[45126] = {9'd67,-10'd334};
ram[45127] = {9'd70,-10'd330};
ram[45128] = {9'd73,-10'd327};
ram[45129] = {9'd76,-10'd324};
ram[45130] = {9'd80,-10'd321};
ram[45131] = {9'd83,-10'd318};
ram[45132] = {9'd86,-10'd315};
ram[45133] = {9'd89,-10'd312};
ram[45134] = {9'd92,-10'd308};
ram[45135] = {9'd95,-10'd305};
ram[45136] = {9'd98,-10'd302};
ram[45137] = {-9'd99,-10'd299};
ram[45138] = {-9'd96,-10'd296};
ram[45139] = {-9'd92,-10'd293};
ram[45140] = {-9'd89,-10'd290};
ram[45141] = {-9'd86,-10'd286};
ram[45142] = {-9'd83,-10'd283};
ram[45143] = {-9'd80,-10'd280};
ram[45144] = {-9'd77,-10'd277};
ram[45145] = {-9'd74,-10'd274};
ram[45146] = {-9'd70,-10'd271};
ram[45147] = {-9'd67,-10'd268};
ram[45148] = {-9'd64,-10'd264};
ram[45149] = {-9'd61,-10'd261};
ram[45150] = {-9'd58,-10'd258};
ram[45151] = {-9'd55,-10'd255};
ram[45152] = {-9'd52,-10'd252};
ram[45153] = {-9'd48,-10'd249};
ram[45154] = {-9'd45,-10'd246};
ram[45155] = {-9'd42,-10'd242};
ram[45156] = {-9'd39,-10'd239};
ram[45157] = {-9'd36,-10'd236};
ram[45158] = {-9'd33,-10'd233};
ram[45159] = {-9'd30,-10'd230};
ram[45160] = {-9'd26,-10'd227};
ram[45161] = {-9'd23,-10'd224};
ram[45162] = {-9'd20,-10'd220};
ram[45163] = {-9'd17,-10'd217};
ram[45164] = {-9'd14,-10'd214};
ram[45165] = {-9'd11,-10'd211};
ram[45166] = {-9'd8,-10'd208};
ram[45167] = {-9'd4,-10'd205};
ram[45168] = {-9'd1,-10'd202};
ram[45169] = {9'd2,-10'd198};
ram[45170] = {9'd5,-10'd195};
ram[45171] = {9'd8,-10'd192};
ram[45172] = {9'd11,-10'd189};
ram[45173] = {9'd14,-10'd186};
ram[45174] = {9'd18,-10'd183};
ram[45175] = {9'd21,-10'd180};
ram[45176] = {9'd24,-10'd176};
ram[45177] = {9'd27,-10'd173};
ram[45178] = {9'd30,-10'd170};
ram[45179] = {9'd33,-10'd167};
ram[45180] = {9'd36,-10'd164};
ram[45181] = {9'd40,-10'd161};
ram[45182] = {9'd43,-10'd158};
ram[45183] = {9'd46,-10'd154};
ram[45184] = {9'd46,-10'd154};
ram[45185] = {9'd49,-10'd151};
ram[45186] = {9'd52,-10'd148};
ram[45187] = {9'd55,-10'd145};
ram[45188] = {9'd58,-10'd142};
ram[45189] = {9'd62,-10'd139};
ram[45190] = {9'd65,-10'd136};
ram[45191] = {9'd68,-10'd132};
ram[45192] = {9'd71,-10'd129};
ram[45193] = {9'd74,-10'd126};
ram[45194] = {9'd77,-10'd123};
ram[45195] = {9'd80,-10'd120};
ram[45196] = {9'd84,-10'd117};
ram[45197] = {9'd87,-10'd114};
ram[45198] = {9'd90,-10'd110};
ram[45199] = {9'd93,-10'd107};
ram[45200] = {9'd96,-10'd104};
ram[45201] = {9'd99,-10'd101};
ram[45202] = {-9'd98,-10'd98};
ram[45203] = {-9'd95,-10'd95};
ram[45204] = {-9'd92,-10'd92};
ram[45205] = {-9'd88,-10'd88};
ram[45206] = {-9'd85,-10'd85};
ram[45207] = {-9'd82,-10'd82};
ram[45208] = {-9'd79,-10'd79};
ram[45209] = {-9'd76,-10'd76};
ram[45210] = {-9'd73,-10'd73};
ram[45211] = {-9'd70,-10'd70};
ram[45212] = {-9'd66,-10'd66};
ram[45213] = {-9'd63,-10'd63};
ram[45214] = {-9'd60,-10'd60};
ram[45215] = {-9'd57,-10'd57};
ram[45216] = {-9'd54,-10'd54};
ram[45217] = {-9'd51,-10'd51};
ram[45218] = {-9'd48,-10'd48};
ram[45219] = {-9'd44,-10'd44};
ram[45220] = {-9'd41,-10'd41};
ram[45221] = {-9'd38,-10'd38};
ram[45222] = {-9'd35,-10'd35};
ram[45223] = {-9'd32,-10'd32};
ram[45224] = {-9'd29,-10'd29};
ram[45225] = {-9'd26,-10'd26};
ram[45226] = {-9'd22,-10'd22};
ram[45227] = {-9'd19,-10'd19};
ram[45228] = {-9'd16,-10'd16};
ram[45229] = {-9'd13,-10'd13};
ram[45230] = {-9'd10,-10'd10};
ram[45231] = {-9'd7,-10'd7};
ram[45232] = {-9'd4,-10'd4};
ram[45233] = {9'd0,10'd0};
ram[45234] = {9'd3,10'd3};
ram[45235] = {9'd6,10'd6};
ram[45236] = {9'd9,10'd9};
ram[45237] = {9'd12,10'd12};
ram[45238] = {9'd15,10'd15};
ram[45239] = {9'd18,10'd18};
ram[45240] = {9'd21,10'd21};
ram[45241] = {9'd25,10'd25};
ram[45242] = {9'd28,10'd28};
ram[45243] = {9'd31,10'd31};
ram[45244] = {9'd34,10'd34};
ram[45245] = {9'd37,10'd37};
ram[45246] = {9'd40,10'd40};
ram[45247] = {9'd43,10'd43};
ram[45248] = {9'd47,10'd47};
ram[45249] = {9'd50,10'd50};
ram[45250] = {9'd53,10'd53};
ram[45251] = {9'd56,10'd56};
ram[45252] = {9'd59,10'd59};
ram[45253] = {9'd62,10'd62};
ram[45254] = {9'd65,10'd65};
ram[45255] = {9'd69,10'd69};
ram[45256] = {9'd72,10'd72};
ram[45257] = {9'd75,10'd75};
ram[45258] = {9'd78,10'd78};
ram[45259] = {9'd81,10'd81};
ram[45260] = {9'd84,10'd84};
ram[45261] = {9'd87,10'd87};
ram[45262] = {9'd91,10'd91};
ram[45263] = {9'd94,10'd94};
ram[45264] = {9'd97,10'd97};
ram[45265] = {-9'd100,10'd100};
ram[45266] = {-9'd97,10'd103};
ram[45267] = {-9'd94,10'd106};
ram[45268] = {-9'd91,10'd109};
ram[45269] = {-9'd88,10'd113};
ram[45270] = {-9'd85,10'd116};
ram[45271] = {-9'd81,10'd119};
ram[45272] = {-9'd78,10'd122};
ram[45273] = {-9'd75,10'd125};
ram[45274] = {-9'd72,10'd128};
ram[45275] = {-9'd69,10'd131};
ram[45276] = {-9'd66,10'd135};
ram[45277] = {-9'd63,10'd138};
ram[45278] = {-9'd59,10'd141};
ram[45279] = {-9'd56,10'd144};
ram[45280] = {-9'd53,10'd147};
ram[45281] = {-9'd50,10'd150};
ram[45282] = {-9'd47,10'd153};
ram[45283] = {-9'd44,10'd157};
ram[45284] = {-9'd41,10'd160};
ram[45285] = {-9'd37,10'd163};
ram[45286] = {-9'd34,10'd166};
ram[45287] = {-9'd31,10'd169};
ram[45288] = {-9'd28,10'd172};
ram[45289] = {-9'd25,10'd175};
ram[45290] = {-9'd22,10'd179};
ram[45291] = {-9'd19,10'd182};
ram[45292] = {-9'd15,10'd185};
ram[45293] = {-9'd12,10'd188};
ram[45294] = {-9'd9,10'd191};
ram[45295] = {-9'd6,10'd194};
ram[45296] = {-9'd3,10'd197};
ram[45297] = {9'd0,10'd201};
ram[45298] = {9'd3,10'd204};
ram[45299] = {9'd7,10'd207};
ram[45300] = {9'd10,10'd210};
ram[45301] = {9'd13,10'd213};
ram[45302] = {9'd16,10'd216};
ram[45303] = {9'd19,10'd219};
ram[45304] = {9'd22,10'd223};
ram[45305] = {9'd25,10'd226};
ram[45306] = {9'd29,10'd229};
ram[45307] = {9'd32,10'd232};
ram[45308] = {9'd35,10'd235};
ram[45309] = {9'd38,10'd238};
ram[45310] = {9'd41,10'd241};
ram[45311] = {9'd44,10'd245};
ram[45312] = {9'd44,10'd245};
ram[45313] = {9'd47,10'd248};
ram[45314] = {9'd51,10'd251};
ram[45315] = {9'd54,10'd254};
ram[45316] = {9'd57,10'd257};
ram[45317] = {9'd60,10'd260};
ram[45318] = {9'd63,10'd263};
ram[45319] = {9'd66,10'd267};
ram[45320] = {9'd69,10'd270};
ram[45321] = {9'd73,10'd273};
ram[45322] = {9'd76,10'd276};
ram[45323] = {9'd79,10'd279};
ram[45324] = {9'd82,10'd282};
ram[45325] = {9'd85,10'd285};
ram[45326] = {9'd88,10'd289};
ram[45327] = {9'd91,10'd292};
ram[45328] = {9'd95,10'd295};
ram[45329] = {9'd98,10'd298};
ram[45330] = {-9'd99,10'd301};
ram[45331] = {-9'd96,10'd304};
ram[45332] = {-9'd93,10'd307};
ram[45333] = {-9'd90,10'd311};
ram[45334] = {-9'd87,10'd314};
ram[45335] = {-9'd84,10'd317};
ram[45336] = {-9'd81,10'd320};
ram[45337] = {-9'd77,10'd323};
ram[45338] = {-9'd74,10'd326};
ram[45339] = {-9'd71,10'd329};
ram[45340] = {-9'd68,10'd333};
ram[45341] = {-9'd65,10'd336};
ram[45342] = {-9'd62,10'd339};
ram[45343] = {-9'd59,10'd342};
ram[45344] = {-9'd55,10'd345};
ram[45345] = {-9'd52,10'd348};
ram[45346] = {-9'd49,10'd351};
ram[45347] = {-9'd46,10'd354};
ram[45348] = {-9'd43,10'd358};
ram[45349] = {-9'd40,10'd361};
ram[45350] = {-9'd37,10'd364};
ram[45351] = {-9'd33,10'd367};
ram[45352] = {-9'd30,10'd370};
ram[45353] = {-9'd27,10'd373};
ram[45354] = {-9'd24,10'd376};
ram[45355] = {-9'd21,10'd380};
ram[45356] = {-9'd18,10'd383};
ram[45357] = {-9'd15,10'd386};
ram[45358] = {-9'd11,10'd389};
ram[45359] = {-9'd8,10'd392};
ram[45360] = {-9'd5,10'd395};
ram[45361] = {-9'd2,10'd398};
ram[45362] = {9'd1,-10'd399};
ram[45363] = {9'd4,-10'd396};
ram[45364] = {9'd7,-10'd393};
ram[45365] = {9'd10,-10'd390};
ram[45366] = {9'd14,-10'd387};
ram[45367] = {9'd17,-10'd384};
ram[45368] = {9'd20,-10'd381};
ram[45369] = {9'd23,-10'd377};
ram[45370] = {9'd26,-10'd374};
ram[45371] = {9'd29,-10'd371};
ram[45372] = {9'd32,-10'd368};
ram[45373] = {9'd36,-10'd365};
ram[45374] = {9'd39,-10'd362};
ram[45375] = {9'd42,-10'd359};
ram[45376] = {9'd45,-10'd355};
ram[45377] = {9'd48,-10'd352};
ram[45378] = {9'd51,-10'd349};
ram[45379] = {9'd54,-10'd346};
ram[45380] = {9'd58,-10'd343};
ram[45381] = {9'd61,-10'd340};
ram[45382] = {9'd64,-10'd337};
ram[45383] = {9'd67,-10'd334};
ram[45384] = {9'd70,-10'd330};
ram[45385] = {9'd73,-10'd327};
ram[45386] = {9'd76,-10'd324};
ram[45387] = {9'd80,-10'd321};
ram[45388] = {9'd83,-10'd318};
ram[45389] = {9'd86,-10'd315};
ram[45390] = {9'd89,-10'd312};
ram[45391] = {9'd92,-10'd308};
ram[45392] = {9'd95,-10'd305};
ram[45393] = {9'd98,-10'd302};
ram[45394] = {-9'd99,-10'd299};
ram[45395] = {-9'd96,-10'd296};
ram[45396] = {-9'd92,-10'd293};
ram[45397] = {-9'd89,-10'd290};
ram[45398] = {-9'd86,-10'd286};
ram[45399] = {-9'd83,-10'd283};
ram[45400] = {-9'd80,-10'd280};
ram[45401] = {-9'd77,-10'd277};
ram[45402] = {-9'd74,-10'd274};
ram[45403] = {-9'd70,-10'd271};
ram[45404] = {-9'd67,-10'd268};
ram[45405] = {-9'd64,-10'd264};
ram[45406] = {-9'd61,-10'd261};
ram[45407] = {-9'd58,-10'd258};
ram[45408] = {-9'd55,-10'd255};
ram[45409] = {-9'd52,-10'd252};
ram[45410] = {-9'd48,-10'd249};
ram[45411] = {-9'd45,-10'd246};
ram[45412] = {-9'd42,-10'd242};
ram[45413] = {-9'd39,-10'd239};
ram[45414] = {-9'd36,-10'd236};
ram[45415] = {-9'd33,-10'd233};
ram[45416] = {-9'd30,-10'd230};
ram[45417] = {-9'd26,-10'd227};
ram[45418] = {-9'd23,-10'd224};
ram[45419] = {-9'd20,-10'd220};
ram[45420] = {-9'd17,-10'd217};
ram[45421] = {-9'd14,-10'd214};
ram[45422] = {-9'd11,-10'd211};
ram[45423] = {-9'd8,-10'd208};
ram[45424] = {-9'd4,-10'd205};
ram[45425] = {-9'd1,-10'd202};
ram[45426] = {9'd2,-10'd198};
ram[45427] = {9'd5,-10'd195};
ram[45428] = {9'd8,-10'd192};
ram[45429] = {9'd11,-10'd189};
ram[45430] = {9'd14,-10'd186};
ram[45431] = {9'd18,-10'd183};
ram[45432] = {9'd21,-10'd180};
ram[45433] = {9'd24,-10'd176};
ram[45434] = {9'd27,-10'd173};
ram[45435] = {9'd30,-10'd170};
ram[45436] = {9'd33,-10'd167};
ram[45437] = {9'd36,-10'd164};
ram[45438] = {9'd40,-10'd161};
ram[45439] = {9'd43,-10'd158};
ram[45440] = {9'd43,-10'd158};
ram[45441] = {9'd46,-10'd154};
ram[45442] = {9'd49,-10'd151};
ram[45443] = {9'd52,-10'd148};
ram[45444] = {9'd55,-10'd145};
ram[45445] = {9'd58,-10'd142};
ram[45446] = {9'd62,-10'd139};
ram[45447] = {9'd65,-10'd136};
ram[45448] = {9'd68,-10'd132};
ram[45449] = {9'd71,-10'd129};
ram[45450] = {9'd74,-10'd126};
ram[45451] = {9'd77,-10'd123};
ram[45452] = {9'd80,-10'd120};
ram[45453] = {9'd84,-10'd117};
ram[45454] = {9'd87,-10'd114};
ram[45455] = {9'd90,-10'd110};
ram[45456] = {9'd93,-10'd107};
ram[45457] = {9'd96,-10'd104};
ram[45458] = {9'd99,-10'd101};
ram[45459] = {-9'd98,-10'd98};
ram[45460] = {-9'd95,-10'd95};
ram[45461] = {-9'd92,-10'd92};
ram[45462] = {-9'd88,-10'd88};
ram[45463] = {-9'd85,-10'd85};
ram[45464] = {-9'd82,-10'd82};
ram[45465] = {-9'd79,-10'd79};
ram[45466] = {-9'd76,-10'd76};
ram[45467] = {-9'd73,-10'd73};
ram[45468] = {-9'd70,-10'd70};
ram[45469] = {-9'd66,-10'd66};
ram[45470] = {-9'd63,-10'd63};
ram[45471] = {-9'd60,-10'd60};
ram[45472] = {-9'd57,-10'd57};
ram[45473] = {-9'd54,-10'd54};
ram[45474] = {-9'd51,-10'd51};
ram[45475] = {-9'd48,-10'd48};
ram[45476] = {-9'd44,-10'd44};
ram[45477] = {-9'd41,-10'd41};
ram[45478] = {-9'd38,-10'd38};
ram[45479] = {-9'd35,-10'd35};
ram[45480] = {-9'd32,-10'd32};
ram[45481] = {-9'd29,-10'd29};
ram[45482] = {-9'd26,-10'd26};
ram[45483] = {-9'd22,-10'd22};
ram[45484] = {-9'd19,-10'd19};
ram[45485] = {-9'd16,-10'd16};
ram[45486] = {-9'd13,-10'd13};
ram[45487] = {-9'd10,-10'd10};
ram[45488] = {-9'd7,-10'd7};
ram[45489] = {-9'd4,-10'd4};
ram[45490] = {9'd0,10'd0};
ram[45491] = {9'd3,10'd3};
ram[45492] = {9'd6,10'd6};
ram[45493] = {9'd9,10'd9};
ram[45494] = {9'd12,10'd12};
ram[45495] = {9'd15,10'd15};
ram[45496] = {9'd18,10'd18};
ram[45497] = {9'd21,10'd21};
ram[45498] = {9'd25,10'd25};
ram[45499] = {9'd28,10'd28};
ram[45500] = {9'd31,10'd31};
ram[45501] = {9'd34,10'd34};
ram[45502] = {9'd37,10'd37};
ram[45503] = {9'd40,10'd40};
ram[45504] = {9'd43,10'd43};
ram[45505] = {9'd47,10'd47};
ram[45506] = {9'd50,10'd50};
ram[45507] = {9'd53,10'd53};
ram[45508] = {9'd56,10'd56};
ram[45509] = {9'd59,10'd59};
ram[45510] = {9'd62,10'd62};
ram[45511] = {9'd65,10'd65};
ram[45512] = {9'd69,10'd69};
ram[45513] = {9'd72,10'd72};
ram[45514] = {9'd75,10'd75};
ram[45515] = {9'd78,10'd78};
ram[45516] = {9'd81,10'd81};
ram[45517] = {9'd84,10'd84};
ram[45518] = {9'd87,10'd87};
ram[45519] = {9'd91,10'd91};
ram[45520] = {9'd94,10'd94};
ram[45521] = {9'd97,10'd97};
ram[45522] = {-9'd100,10'd100};
ram[45523] = {-9'd97,10'd103};
ram[45524] = {-9'd94,10'd106};
ram[45525] = {-9'd91,10'd109};
ram[45526] = {-9'd88,10'd113};
ram[45527] = {-9'd85,10'd116};
ram[45528] = {-9'd81,10'd119};
ram[45529] = {-9'd78,10'd122};
ram[45530] = {-9'd75,10'd125};
ram[45531] = {-9'd72,10'd128};
ram[45532] = {-9'd69,10'd131};
ram[45533] = {-9'd66,10'd135};
ram[45534] = {-9'd63,10'd138};
ram[45535] = {-9'd59,10'd141};
ram[45536] = {-9'd56,10'd144};
ram[45537] = {-9'd53,10'd147};
ram[45538] = {-9'd50,10'd150};
ram[45539] = {-9'd47,10'd153};
ram[45540] = {-9'd44,10'd157};
ram[45541] = {-9'd41,10'd160};
ram[45542] = {-9'd37,10'd163};
ram[45543] = {-9'd34,10'd166};
ram[45544] = {-9'd31,10'd169};
ram[45545] = {-9'd28,10'd172};
ram[45546] = {-9'd25,10'd175};
ram[45547] = {-9'd22,10'd179};
ram[45548] = {-9'd19,10'd182};
ram[45549] = {-9'd15,10'd185};
ram[45550] = {-9'd12,10'd188};
ram[45551] = {-9'd9,10'd191};
ram[45552] = {-9'd6,10'd194};
ram[45553] = {-9'd3,10'd197};
ram[45554] = {9'd0,10'd201};
ram[45555] = {9'd3,10'd204};
ram[45556] = {9'd7,10'd207};
ram[45557] = {9'd10,10'd210};
ram[45558] = {9'd13,10'd213};
ram[45559] = {9'd16,10'd216};
ram[45560] = {9'd19,10'd219};
ram[45561] = {9'd22,10'd223};
ram[45562] = {9'd25,10'd226};
ram[45563] = {9'd29,10'd229};
ram[45564] = {9'd32,10'd232};
ram[45565] = {9'd35,10'd235};
ram[45566] = {9'd38,10'd238};
ram[45567] = {9'd41,10'd241};
ram[45568] = {9'd41,10'd241};
ram[45569] = {9'd44,10'd245};
ram[45570] = {9'd47,10'd248};
ram[45571] = {9'd51,10'd251};
ram[45572] = {9'd54,10'd254};
ram[45573] = {9'd57,10'd257};
ram[45574] = {9'd60,10'd260};
ram[45575] = {9'd63,10'd263};
ram[45576] = {9'd66,10'd267};
ram[45577] = {9'd69,10'd270};
ram[45578] = {9'd73,10'd273};
ram[45579] = {9'd76,10'd276};
ram[45580] = {9'd79,10'd279};
ram[45581] = {9'd82,10'd282};
ram[45582] = {9'd85,10'd285};
ram[45583] = {9'd88,10'd289};
ram[45584] = {9'd91,10'd292};
ram[45585] = {9'd95,10'd295};
ram[45586] = {9'd98,10'd298};
ram[45587] = {-9'd99,10'd301};
ram[45588] = {-9'd96,10'd304};
ram[45589] = {-9'd93,10'd307};
ram[45590] = {-9'd90,10'd311};
ram[45591] = {-9'd87,10'd314};
ram[45592] = {-9'd84,10'd317};
ram[45593] = {-9'd81,10'd320};
ram[45594] = {-9'd77,10'd323};
ram[45595] = {-9'd74,10'd326};
ram[45596] = {-9'd71,10'd329};
ram[45597] = {-9'd68,10'd333};
ram[45598] = {-9'd65,10'd336};
ram[45599] = {-9'd62,10'd339};
ram[45600] = {-9'd59,10'd342};
ram[45601] = {-9'd55,10'd345};
ram[45602] = {-9'd52,10'd348};
ram[45603] = {-9'd49,10'd351};
ram[45604] = {-9'd46,10'd354};
ram[45605] = {-9'd43,10'd358};
ram[45606] = {-9'd40,10'd361};
ram[45607] = {-9'd37,10'd364};
ram[45608] = {-9'd33,10'd367};
ram[45609] = {-9'd30,10'd370};
ram[45610] = {-9'd27,10'd373};
ram[45611] = {-9'd24,10'd376};
ram[45612] = {-9'd21,10'd380};
ram[45613] = {-9'd18,10'd383};
ram[45614] = {-9'd15,10'd386};
ram[45615] = {-9'd11,10'd389};
ram[45616] = {-9'd8,10'd392};
ram[45617] = {-9'd5,10'd395};
ram[45618] = {-9'd2,10'd398};
ram[45619] = {9'd1,-10'd399};
ram[45620] = {9'd4,-10'd396};
ram[45621] = {9'd7,-10'd393};
ram[45622] = {9'd10,-10'd390};
ram[45623] = {9'd14,-10'd387};
ram[45624] = {9'd17,-10'd384};
ram[45625] = {9'd20,-10'd381};
ram[45626] = {9'd23,-10'd377};
ram[45627] = {9'd26,-10'd374};
ram[45628] = {9'd29,-10'd371};
ram[45629] = {9'd32,-10'd368};
ram[45630] = {9'd36,-10'd365};
ram[45631] = {9'd39,-10'd362};
ram[45632] = {9'd42,-10'd359};
ram[45633] = {9'd45,-10'd355};
ram[45634] = {9'd48,-10'd352};
ram[45635] = {9'd51,-10'd349};
ram[45636] = {9'd54,-10'd346};
ram[45637] = {9'd58,-10'd343};
ram[45638] = {9'd61,-10'd340};
ram[45639] = {9'd64,-10'd337};
ram[45640] = {9'd67,-10'd334};
ram[45641] = {9'd70,-10'd330};
ram[45642] = {9'd73,-10'd327};
ram[45643] = {9'd76,-10'd324};
ram[45644] = {9'd80,-10'd321};
ram[45645] = {9'd83,-10'd318};
ram[45646] = {9'd86,-10'd315};
ram[45647] = {9'd89,-10'd312};
ram[45648] = {9'd92,-10'd308};
ram[45649] = {9'd95,-10'd305};
ram[45650] = {9'd98,-10'd302};
ram[45651] = {-9'd99,-10'd299};
ram[45652] = {-9'd96,-10'd296};
ram[45653] = {-9'd92,-10'd293};
ram[45654] = {-9'd89,-10'd290};
ram[45655] = {-9'd86,-10'd286};
ram[45656] = {-9'd83,-10'd283};
ram[45657] = {-9'd80,-10'd280};
ram[45658] = {-9'd77,-10'd277};
ram[45659] = {-9'd74,-10'd274};
ram[45660] = {-9'd70,-10'd271};
ram[45661] = {-9'd67,-10'd268};
ram[45662] = {-9'd64,-10'd264};
ram[45663] = {-9'd61,-10'd261};
ram[45664] = {-9'd58,-10'd258};
ram[45665] = {-9'd55,-10'd255};
ram[45666] = {-9'd52,-10'd252};
ram[45667] = {-9'd48,-10'd249};
ram[45668] = {-9'd45,-10'd246};
ram[45669] = {-9'd42,-10'd242};
ram[45670] = {-9'd39,-10'd239};
ram[45671] = {-9'd36,-10'd236};
ram[45672] = {-9'd33,-10'd233};
ram[45673] = {-9'd30,-10'd230};
ram[45674] = {-9'd26,-10'd227};
ram[45675] = {-9'd23,-10'd224};
ram[45676] = {-9'd20,-10'd220};
ram[45677] = {-9'd17,-10'd217};
ram[45678] = {-9'd14,-10'd214};
ram[45679] = {-9'd11,-10'd211};
ram[45680] = {-9'd8,-10'd208};
ram[45681] = {-9'd4,-10'd205};
ram[45682] = {-9'd1,-10'd202};
ram[45683] = {9'd2,-10'd198};
ram[45684] = {9'd5,-10'd195};
ram[45685] = {9'd8,-10'd192};
ram[45686] = {9'd11,-10'd189};
ram[45687] = {9'd14,-10'd186};
ram[45688] = {9'd18,-10'd183};
ram[45689] = {9'd21,-10'd180};
ram[45690] = {9'd24,-10'd176};
ram[45691] = {9'd27,-10'd173};
ram[45692] = {9'd30,-10'd170};
ram[45693] = {9'd33,-10'd167};
ram[45694] = {9'd36,-10'd164};
ram[45695] = {9'd40,-10'd161};
ram[45696] = {9'd40,-10'd161};
ram[45697] = {9'd43,-10'd158};
ram[45698] = {9'd46,-10'd154};
ram[45699] = {9'd49,-10'd151};
ram[45700] = {9'd52,-10'd148};
ram[45701] = {9'd55,-10'd145};
ram[45702] = {9'd58,-10'd142};
ram[45703] = {9'd62,-10'd139};
ram[45704] = {9'd65,-10'd136};
ram[45705] = {9'd68,-10'd132};
ram[45706] = {9'd71,-10'd129};
ram[45707] = {9'd74,-10'd126};
ram[45708] = {9'd77,-10'd123};
ram[45709] = {9'd80,-10'd120};
ram[45710] = {9'd84,-10'd117};
ram[45711] = {9'd87,-10'd114};
ram[45712] = {9'd90,-10'd110};
ram[45713] = {9'd93,-10'd107};
ram[45714] = {9'd96,-10'd104};
ram[45715] = {9'd99,-10'd101};
ram[45716] = {-9'd98,-10'd98};
ram[45717] = {-9'd95,-10'd95};
ram[45718] = {-9'd92,-10'd92};
ram[45719] = {-9'd88,-10'd88};
ram[45720] = {-9'd85,-10'd85};
ram[45721] = {-9'd82,-10'd82};
ram[45722] = {-9'd79,-10'd79};
ram[45723] = {-9'd76,-10'd76};
ram[45724] = {-9'd73,-10'd73};
ram[45725] = {-9'd70,-10'd70};
ram[45726] = {-9'd66,-10'd66};
ram[45727] = {-9'd63,-10'd63};
ram[45728] = {-9'd60,-10'd60};
ram[45729] = {-9'd57,-10'd57};
ram[45730] = {-9'd54,-10'd54};
ram[45731] = {-9'd51,-10'd51};
ram[45732] = {-9'd48,-10'd48};
ram[45733] = {-9'd44,-10'd44};
ram[45734] = {-9'd41,-10'd41};
ram[45735] = {-9'd38,-10'd38};
ram[45736] = {-9'd35,-10'd35};
ram[45737] = {-9'd32,-10'd32};
ram[45738] = {-9'd29,-10'd29};
ram[45739] = {-9'd26,-10'd26};
ram[45740] = {-9'd22,-10'd22};
ram[45741] = {-9'd19,-10'd19};
ram[45742] = {-9'd16,-10'd16};
ram[45743] = {-9'd13,-10'd13};
ram[45744] = {-9'd10,-10'd10};
ram[45745] = {-9'd7,-10'd7};
ram[45746] = {-9'd4,-10'd4};
ram[45747] = {9'd0,10'd0};
ram[45748] = {9'd3,10'd3};
ram[45749] = {9'd6,10'd6};
ram[45750] = {9'd9,10'd9};
ram[45751] = {9'd12,10'd12};
ram[45752] = {9'd15,10'd15};
ram[45753] = {9'd18,10'd18};
ram[45754] = {9'd21,10'd21};
ram[45755] = {9'd25,10'd25};
ram[45756] = {9'd28,10'd28};
ram[45757] = {9'd31,10'd31};
ram[45758] = {9'd34,10'd34};
ram[45759] = {9'd37,10'd37};
ram[45760] = {9'd40,10'd40};
ram[45761] = {9'd43,10'd43};
ram[45762] = {9'd47,10'd47};
ram[45763] = {9'd50,10'd50};
ram[45764] = {9'd53,10'd53};
ram[45765] = {9'd56,10'd56};
ram[45766] = {9'd59,10'd59};
ram[45767] = {9'd62,10'd62};
ram[45768] = {9'd65,10'd65};
ram[45769] = {9'd69,10'd69};
ram[45770] = {9'd72,10'd72};
ram[45771] = {9'd75,10'd75};
ram[45772] = {9'd78,10'd78};
ram[45773] = {9'd81,10'd81};
ram[45774] = {9'd84,10'd84};
ram[45775] = {9'd87,10'd87};
ram[45776] = {9'd91,10'd91};
ram[45777] = {9'd94,10'd94};
ram[45778] = {9'd97,10'd97};
ram[45779] = {-9'd100,10'd100};
ram[45780] = {-9'd97,10'd103};
ram[45781] = {-9'd94,10'd106};
ram[45782] = {-9'd91,10'd109};
ram[45783] = {-9'd88,10'd113};
ram[45784] = {-9'd85,10'd116};
ram[45785] = {-9'd81,10'd119};
ram[45786] = {-9'd78,10'd122};
ram[45787] = {-9'd75,10'd125};
ram[45788] = {-9'd72,10'd128};
ram[45789] = {-9'd69,10'd131};
ram[45790] = {-9'd66,10'd135};
ram[45791] = {-9'd63,10'd138};
ram[45792] = {-9'd59,10'd141};
ram[45793] = {-9'd56,10'd144};
ram[45794] = {-9'd53,10'd147};
ram[45795] = {-9'd50,10'd150};
ram[45796] = {-9'd47,10'd153};
ram[45797] = {-9'd44,10'd157};
ram[45798] = {-9'd41,10'd160};
ram[45799] = {-9'd37,10'd163};
ram[45800] = {-9'd34,10'd166};
ram[45801] = {-9'd31,10'd169};
ram[45802] = {-9'd28,10'd172};
ram[45803] = {-9'd25,10'd175};
ram[45804] = {-9'd22,10'd179};
ram[45805] = {-9'd19,10'd182};
ram[45806] = {-9'd15,10'd185};
ram[45807] = {-9'd12,10'd188};
ram[45808] = {-9'd9,10'd191};
ram[45809] = {-9'd6,10'd194};
ram[45810] = {-9'd3,10'd197};
ram[45811] = {9'd0,10'd201};
ram[45812] = {9'd3,10'd204};
ram[45813] = {9'd7,10'd207};
ram[45814] = {9'd10,10'd210};
ram[45815] = {9'd13,10'd213};
ram[45816] = {9'd16,10'd216};
ram[45817] = {9'd19,10'd219};
ram[45818] = {9'd22,10'd223};
ram[45819] = {9'd25,10'd226};
ram[45820] = {9'd29,10'd229};
ram[45821] = {9'd32,10'd232};
ram[45822] = {9'd35,10'd235};
ram[45823] = {9'd38,10'd238};
ram[45824] = {9'd38,10'd238};
ram[45825] = {9'd41,10'd241};
ram[45826] = {9'd44,10'd245};
ram[45827] = {9'd47,10'd248};
ram[45828] = {9'd51,10'd251};
ram[45829] = {9'd54,10'd254};
ram[45830] = {9'd57,10'd257};
ram[45831] = {9'd60,10'd260};
ram[45832] = {9'd63,10'd263};
ram[45833] = {9'd66,10'd267};
ram[45834] = {9'd69,10'd270};
ram[45835] = {9'd73,10'd273};
ram[45836] = {9'd76,10'd276};
ram[45837] = {9'd79,10'd279};
ram[45838] = {9'd82,10'd282};
ram[45839] = {9'd85,10'd285};
ram[45840] = {9'd88,10'd289};
ram[45841] = {9'd91,10'd292};
ram[45842] = {9'd95,10'd295};
ram[45843] = {9'd98,10'd298};
ram[45844] = {-9'd99,10'd301};
ram[45845] = {-9'd96,10'd304};
ram[45846] = {-9'd93,10'd307};
ram[45847] = {-9'd90,10'd311};
ram[45848] = {-9'd87,10'd314};
ram[45849] = {-9'd84,10'd317};
ram[45850] = {-9'd81,10'd320};
ram[45851] = {-9'd77,10'd323};
ram[45852] = {-9'd74,10'd326};
ram[45853] = {-9'd71,10'd329};
ram[45854] = {-9'd68,10'd333};
ram[45855] = {-9'd65,10'd336};
ram[45856] = {-9'd62,10'd339};
ram[45857] = {-9'd59,10'd342};
ram[45858] = {-9'd55,10'd345};
ram[45859] = {-9'd52,10'd348};
ram[45860] = {-9'd49,10'd351};
ram[45861] = {-9'd46,10'd354};
ram[45862] = {-9'd43,10'd358};
ram[45863] = {-9'd40,10'd361};
ram[45864] = {-9'd37,10'd364};
ram[45865] = {-9'd33,10'd367};
ram[45866] = {-9'd30,10'd370};
ram[45867] = {-9'd27,10'd373};
ram[45868] = {-9'd24,10'd376};
ram[45869] = {-9'd21,10'd380};
ram[45870] = {-9'd18,10'd383};
ram[45871] = {-9'd15,10'd386};
ram[45872] = {-9'd11,10'd389};
ram[45873] = {-9'd8,10'd392};
ram[45874] = {-9'd5,10'd395};
ram[45875] = {-9'd2,10'd398};
ram[45876] = {9'd1,-10'd399};
ram[45877] = {9'd4,-10'd396};
ram[45878] = {9'd7,-10'd393};
ram[45879] = {9'd10,-10'd390};
ram[45880] = {9'd14,-10'd387};
ram[45881] = {9'd17,-10'd384};
ram[45882] = {9'd20,-10'd381};
ram[45883] = {9'd23,-10'd377};
ram[45884] = {9'd26,-10'd374};
ram[45885] = {9'd29,-10'd371};
ram[45886] = {9'd32,-10'd368};
ram[45887] = {9'd36,-10'd365};
ram[45888] = {9'd39,-10'd362};
ram[45889] = {9'd42,-10'd359};
ram[45890] = {9'd45,-10'd355};
ram[45891] = {9'd48,-10'd352};
ram[45892] = {9'd51,-10'd349};
ram[45893] = {9'd54,-10'd346};
ram[45894] = {9'd58,-10'd343};
ram[45895] = {9'd61,-10'd340};
ram[45896] = {9'd64,-10'd337};
ram[45897] = {9'd67,-10'd334};
ram[45898] = {9'd70,-10'd330};
ram[45899] = {9'd73,-10'd327};
ram[45900] = {9'd76,-10'd324};
ram[45901] = {9'd80,-10'd321};
ram[45902] = {9'd83,-10'd318};
ram[45903] = {9'd86,-10'd315};
ram[45904] = {9'd89,-10'd312};
ram[45905] = {9'd92,-10'd308};
ram[45906] = {9'd95,-10'd305};
ram[45907] = {9'd98,-10'd302};
ram[45908] = {-9'd99,-10'd299};
ram[45909] = {-9'd96,-10'd296};
ram[45910] = {-9'd92,-10'd293};
ram[45911] = {-9'd89,-10'd290};
ram[45912] = {-9'd86,-10'd286};
ram[45913] = {-9'd83,-10'd283};
ram[45914] = {-9'd80,-10'd280};
ram[45915] = {-9'd77,-10'd277};
ram[45916] = {-9'd74,-10'd274};
ram[45917] = {-9'd70,-10'd271};
ram[45918] = {-9'd67,-10'd268};
ram[45919] = {-9'd64,-10'd264};
ram[45920] = {-9'd61,-10'd261};
ram[45921] = {-9'd58,-10'd258};
ram[45922] = {-9'd55,-10'd255};
ram[45923] = {-9'd52,-10'd252};
ram[45924] = {-9'd48,-10'd249};
ram[45925] = {-9'd45,-10'd246};
ram[45926] = {-9'd42,-10'd242};
ram[45927] = {-9'd39,-10'd239};
ram[45928] = {-9'd36,-10'd236};
ram[45929] = {-9'd33,-10'd233};
ram[45930] = {-9'd30,-10'd230};
ram[45931] = {-9'd26,-10'd227};
ram[45932] = {-9'd23,-10'd224};
ram[45933] = {-9'd20,-10'd220};
ram[45934] = {-9'd17,-10'd217};
ram[45935] = {-9'd14,-10'd214};
ram[45936] = {-9'd11,-10'd211};
ram[45937] = {-9'd8,-10'd208};
ram[45938] = {-9'd4,-10'd205};
ram[45939] = {-9'd1,-10'd202};
ram[45940] = {9'd2,-10'd198};
ram[45941] = {9'd5,-10'd195};
ram[45942] = {9'd8,-10'd192};
ram[45943] = {9'd11,-10'd189};
ram[45944] = {9'd14,-10'd186};
ram[45945] = {9'd18,-10'd183};
ram[45946] = {9'd21,-10'd180};
ram[45947] = {9'd24,-10'd176};
ram[45948] = {9'd27,-10'd173};
ram[45949] = {9'd30,-10'd170};
ram[45950] = {9'd33,-10'd167};
ram[45951] = {9'd36,-10'd164};
ram[45952] = {9'd36,-10'd164};
ram[45953] = {9'd40,-10'd161};
ram[45954] = {9'd43,-10'd158};
ram[45955] = {9'd46,-10'd154};
ram[45956] = {9'd49,-10'd151};
ram[45957] = {9'd52,-10'd148};
ram[45958] = {9'd55,-10'd145};
ram[45959] = {9'd58,-10'd142};
ram[45960] = {9'd62,-10'd139};
ram[45961] = {9'd65,-10'd136};
ram[45962] = {9'd68,-10'd132};
ram[45963] = {9'd71,-10'd129};
ram[45964] = {9'd74,-10'd126};
ram[45965] = {9'd77,-10'd123};
ram[45966] = {9'd80,-10'd120};
ram[45967] = {9'd84,-10'd117};
ram[45968] = {9'd87,-10'd114};
ram[45969] = {9'd90,-10'd110};
ram[45970] = {9'd93,-10'd107};
ram[45971] = {9'd96,-10'd104};
ram[45972] = {9'd99,-10'd101};
ram[45973] = {-9'd98,-10'd98};
ram[45974] = {-9'd95,-10'd95};
ram[45975] = {-9'd92,-10'd92};
ram[45976] = {-9'd88,-10'd88};
ram[45977] = {-9'd85,-10'd85};
ram[45978] = {-9'd82,-10'd82};
ram[45979] = {-9'd79,-10'd79};
ram[45980] = {-9'd76,-10'd76};
ram[45981] = {-9'd73,-10'd73};
ram[45982] = {-9'd70,-10'd70};
ram[45983] = {-9'd66,-10'd66};
ram[45984] = {-9'd63,-10'd63};
ram[45985] = {-9'd60,-10'd60};
ram[45986] = {-9'd57,-10'd57};
ram[45987] = {-9'd54,-10'd54};
ram[45988] = {-9'd51,-10'd51};
ram[45989] = {-9'd48,-10'd48};
ram[45990] = {-9'd44,-10'd44};
ram[45991] = {-9'd41,-10'd41};
ram[45992] = {-9'd38,-10'd38};
ram[45993] = {-9'd35,-10'd35};
ram[45994] = {-9'd32,-10'd32};
ram[45995] = {-9'd29,-10'd29};
ram[45996] = {-9'd26,-10'd26};
ram[45997] = {-9'd22,-10'd22};
ram[45998] = {-9'd19,-10'd19};
ram[45999] = {-9'd16,-10'd16};
ram[46000] = {-9'd13,-10'd13};
ram[46001] = {-9'd10,-10'd10};
ram[46002] = {-9'd7,-10'd7};
ram[46003] = {-9'd4,-10'd4};
ram[46004] = {9'd0,10'd0};
ram[46005] = {9'd3,10'd3};
ram[46006] = {9'd6,10'd6};
ram[46007] = {9'd9,10'd9};
ram[46008] = {9'd12,10'd12};
ram[46009] = {9'd15,10'd15};
ram[46010] = {9'd18,10'd18};
ram[46011] = {9'd21,10'd21};
ram[46012] = {9'd25,10'd25};
ram[46013] = {9'd28,10'd28};
ram[46014] = {9'd31,10'd31};
ram[46015] = {9'd34,10'd34};
ram[46016] = {9'd37,10'd37};
ram[46017] = {9'd40,10'd40};
ram[46018] = {9'd43,10'd43};
ram[46019] = {9'd47,10'd47};
ram[46020] = {9'd50,10'd50};
ram[46021] = {9'd53,10'd53};
ram[46022] = {9'd56,10'd56};
ram[46023] = {9'd59,10'd59};
ram[46024] = {9'd62,10'd62};
ram[46025] = {9'd65,10'd65};
ram[46026] = {9'd69,10'd69};
ram[46027] = {9'd72,10'd72};
ram[46028] = {9'd75,10'd75};
ram[46029] = {9'd78,10'd78};
ram[46030] = {9'd81,10'd81};
ram[46031] = {9'd84,10'd84};
ram[46032] = {9'd87,10'd87};
ram[46033] = {9'd91,10'd91};
ram[46034] = {9'd94,10'd94};
ram[46035] = {9'd97,10'd97};
ram[46036] = {-9'd100,10'd100};
ram[46037] = {-9'd97,10'd103};
ram[46038] = {-9'd94,10'd106};
ram[46039] = {-9'd91,10'd109};
ram[46040] = {-9'd88,10'd113};
ram[46041] = {-9'd85,10'd116};
ram[46042] = {-9'd81,10'd119};
ram[46043] = {-9'd78,10'd122};
ram[46044] = {-9'd75,10'd125};
ram[46045] = {-9'd72,10'd128};
ram[46046] = {-9'd69,10'd131};
ram[46047] = {-9'd66,10'd135};
ram[46048] = {-9'd63,10'd138};
ram[46049] = {-9'd59,10'd141};
ram[46050] = {-9'd56,10'd144};
ram[46051] = {-9'd53,10'd147};
ram[46052] = {-9'd50,10'd150};
ram[46053] = {-9'd47,10'd153};
ram[46054] = {-9'd44,10'd157};
ram[46055] = {-9'd41,10'd160};
ram[46056] = {-9'd37,10'd163};
ram[46057] = {-9'd34,10'd166};
ram[46058] = {-9'd31,10'd169};
ram[46059] = {-9'd28,10'd172};
ram[46060] = {-9'd25,10'd175};
ram[46061] = {-9'd22,10'd179};
ram[46062] = {-9'd19,10'd182};
ram[46063] = {-9'd15,10'd185};
ram[46064] = {-9'd12,10'd188};
ram[46065] = {-9'd9,10'd191};
ram[46066] = {-9'd6,10'd194};
ram[46067] = {-9'd3,10'd197};
ram[46068] = {9'd0,10'd201};
ram[46069] = {9'd3,10'd204};
ram[46070] = {9'd7,10'd207};
ram[46071] = {9'd10,10'd210};
ram[46072] = {9'd13,10'd213};
ram[46073] = {9'd16,10'd216};
ram[46074] = {9'd19,10'd219};
ram[46075] = {9'd22,10'd223};
ram[46076] = {9'd25,10'd226};
ram[46077] = {9'd29,10'd229};
ram[46078] = {9'd32,10'd232};
ram[46079] = {9'd35,10'd235};
ram[46080] = {9'd35,10'd235};
ram[46081] = {9'd38,10'd238};
ram[46082] = {9'd41,10'd241};
ram[46083] = {9'd44,10'd245};
ram[46084] = {9'd47,10'd248};
ram[46085] = {9'd51,10'd251};
ram[46086] = {9'd54,10'd254};
ram[46087] = {9'd57,10'd257};
ram[46088] = {9'd60,10'd260};
ram[46089] = {9'd63,10'd263};
ram[46090] = {9'd66,10'd267};
ram[46091] = {9'd69,10'd270};
ram[46092] = {9'd73,10'd273};
ram[46093] = {9'd76,10'd276};
ram[46094] = {9'd79,10'd279};
ram[46095] = {9'd82,10'd282};
ram[46096] = {9'd85,10'd285};
ram[46097] = {9'd88,10'd289};
ram[46098] = {9'd91,10'd292};
ram[46099] = {9'd95,10'd295};
ram[46100] = {9'd98,10'd298};
ram[46101] = {-9'd99,10'd301};
ram[46102] = {-9'd96,10'd304};
ram[46103] = {-9'd93,10'd307};
ram[46104] = {-9'd90,10'd311};
ram[46105] = {-9'd87,10'd314};
ram[46106] = {-9'd84,10'd317};
ram[46107] = {-9'd81,10'd320};
ram[46108] = {-9'd77,10'd323};
ram[46109] = {-9'd74,10'd326};
ram[46110] = {-9'd71,10'd329};
ram[46111] = {-9'd68,10'd333};
ram[46112] = {-9'd65,10'd336};
ram[46113] = {-9'd62,10'd339};
ram[46114] = {-9'd59,10'd342};
ram[46115] = {-9'd55,10'd345};
ram[46116] = {-9'd52,10'd348};
ram[46117] = {-9'd49,10'd351};
ram[46118] = {-9'd46,10'd354};
ram[46119] = {-9'd43,10'd358};
ram[46120] = {-9'd40,10'd361};
ram[46121] = {-9'd37,10'd364};
ram[46122] = {-9'd33,10'd367};
ram[46123] = {-9'd30,10'd370};
ram[46124] = {-9'd27,10'd373};
ram[46125] = {-9'd24,10'd376};
ram[46126] = {-9'd21,10'd380};
ram[46127] = {-9'd18,10'd383};
ram[46128] = {-9'd15,10'd386};
ram[46129] = {-9'd11,10'd389};
ram[46130] = {-9'd8,10'd392};
ram[46131] = {-9'd5,10'd395};
ram[46132] = {-9'd2,10'd398};
ram[46133] = {9'd1,-10'd399};
ram[46134] = {9'd4,-10'd396};
ram[46135] = {9'd7,-10'd393};
ram[46136] = {9'd10,-10'd390};
ram[46137] = {9'd14,-10'd387};
ram[46138] = {9'd17,-10'd384};
ram[46139] = {9'd20,-10'd381};
ram[46140] = {9'd23,-10'd377};
ram[46141] = {9'd26,-10'd374};
ram[46142] = {9'd29,-10'd371};
ram[46143] = {9'd32,-10'd368};
ram[46144] = {9'd36,-10'd365};
ram[46145] = {9'd39,-10'd362};
ram[46146] = {9'd42,-10'd359};
ram[46147] = {9'd45,-10'd355};
ram[46148] = {9'd48,-10'd352};
ram[46149] = {9'd51,-10'd349};
ram[46150] = {9'd54,-10'd346};
ram[46151] = {9'd58,-10'd343};
ram[46152] = {9'd61,-10'd340};
ram[46153] = {9'd64,-10'd337};
ram[46154] = {9'd67,-10'd334};
ram[46155] = {9'd70,-10'd330};
ram[46156] = {9'd73,-10'd327};
ram[46157] = {9'd76,-10'd324};
ram[46158] = {9'd80,-10'd321};
ram[46159] = {9'd83,-10'd318};
ram[46160] = {9'd86,-10'd315};
ram[46161] = {9'd89,-10'd312};
ram[46162] = {9'd92,-10'd308};
ram[46163] = {9'd95,-10'd305};
ram[46164] = {9'd98,-10'd302};
ram[46165] = {-9'd99,-10'd299};
ram[46166] = {-9'd96,-10'd296};
ram[46167] = {-9'd92,-10'd293};
ram[46168] = {-9'd89,-10'd290};
ram[46169] = {-9'd86,-10'd286};
ram[46170] = {-9'd83,-10'd283};
ram[46171] = {-9'd80,-10'd280};
ram[46172] = {-9'd77,-10'd277};
ram[46173] = {-9'd74,-10'd274};
ram[46174] = {-9'd70,-10'd271};
ram[46175] = {-9'd67,-10'd268};
ram[46176] = {-9'd64,-10'd264};
ram[46177] = {-9'd61,-10'd261};
ram[46178] = {-9'd58,-10'd258};
ram[46179] = {-9'd55,-10'd255};
ram[46180] = {-9'd52,-10'd252};
ram[46181] = {-9'd48,-10'd249};
ram[46182] = {-9'd45,-10'd246};
ram[46183] = {-9'd42,-10'd242};
ram[46184] = {-9'd39,-10'd239};
ram[46185] = {-9'd36,-10'd236};
ram[46186] = {-9'd33,-10'd233};
ram[46187] = {-9'd30,-10'd230};
ram[46188] = {-9'd26,-10'd227};
ram[46189] = {-9'd23,-10'd224};
ram[46190] = {-9'd20,-10'd220};
ram[46191] = {-9'd17,-10'd217};
ram[46192] = {-9'd14,-10'd214};
ram[46193] = {-9'd11,-10'd211};
ram[46194] = {-9'd8,-10'd208};
ram[46195] = {-9'd4,-10'd205};
ram[46196] = {-9'd1,-10'd202};
ram[46197] = {9'd2,-10'd198};
ram[46198] = {9'd5,-10'd195};
ram[46199] = {9'd8,-10'd192};
ram[46200] = {9'd11,-10'd189};
ram[46201] = {9'd14,-10'd186};
ram[46202] = {9'd18,-10'd183};
ram[46203] = {9'd21,-10'd180};
ram[46204] = {9'd24,-10'd176};
ram[46205] = {9'd27,-10'd173};
ram[46206] = {9'd30,-10'd170};
ram[46207] = {9'd33,-10'd167};
ram[46208] = {9'd33,-10'd167};
ram[46209] = {9'd36,-10'd164};
ram[46210] = {9'd40,-10'd161};
ram[46211] = {9'd43,-10'd158};
ram[46212] = {9'd46,-10'd154};
ram[46213] = {9'd49,-10'd151};
ram[46214] = {9'd52,-10'd148};
ram[46215] = {9'd55,-10'd145};
ram[46216] = {9'd58,-10'd142};
ram[46217] = {9'd62,-10'd139};
ram[46218] = {9'd65,-10'd136};
ram[46219] = {9'd68,-10'd132};
ram[46220] = {9'd71,-10'd129};
ram[46221] = {9'd74,-10'd126};
ram[46222] = {9'd77,-10'd123};
ram[46223] = {9'd80,-10'd120};
ram[46224] = {9'd84,-10'd117};
ram[46225] = {9'd87,-10'd114};
ram[46226] = {9'd90,-10'd110};
ram[46227] = {9'd93,-10'd107};
ram[46228] = {9'd96,-10'd104};
ram[46229] = {9'd99,-10'd101};
ram[46230] = {-9'd98,-10'd98};
ram[46231] = {-9'd95,-10'd95};
ram[46232] = {-9'd92,-10'd92};
ram[46233] = {-9'd88,-10'd88};
ram[46234] = {-9'd85,-10'd85};
ram[46235] = {-9'd82,-10'd82};
ram[46236] = {-9'd79,-10'd79};
ram[46237] = {-9'd76,-10'd76};
ram[46238] = {-9'd73,-10'd73};
ram[46239] = {-9'd70,-10'd70};
ram[46240] = {-9'd66,-10'd66};
ram[46241] = {-9'd63,-10'd63};
ram[46242] = {-9'd60,-10'd60};
ram[46243] = {-9'd57,-10'd57};
ram[46244] = {-9'd54,-10'd54};
ram[46245] = {-9'd51,-10'd51};
ram[46246] = {-9'd48,-10'd48};
ram[46247] = {-9'd44,-10'd44};
ram[46248] = {-9'd41,-10'd41};
ram[46249] = {-9'd38,-10'd38};
ram[46250] = {-9'd35,-10'd35};
ram[46251] = {-9'd32,-10'd32};
ram[46252] = {-9'd29,-10'd29};
ram[46253] = {-9'd26,-10'd26};
ram[46254] = {-9'd22,-10'd22};
ram[46255] = {-9'd19,-10'd19};
ram[46256] = {-9'd16,-10'd16};
ram[46257] = {-9'd13,-10'd13};
ram[46258] = {-9'd10,-10'd10};
ram[46259] = {-9'd7,-10'd7};
ram[46260] = {-9'd4,-10'd4};
ram[46261] = {9'd0,10'd0};
ram[46262] = {9'd3,10'd3};
ram[46263] = {9'd6,10'd6};
ram[46264] = {9'd9,10'd9};
ram[46265] = {9'd12,10'd12};
ram[46266] = {9'd15,10'd15};
ram[46267] = {9'd18,10'd18};
ram[46268] = {9'd21,10'd21};
ram[46269] = {9'd25,10'd25};
ram[46270] = {9'd28,10'd28};
ram[46271] = {9'd31,10'd31};
ram[46272] = {9'd34,10'd34};
ram[46273] = {9'd37,10'd37};
ram[46274] = {9'd40,10'd40};
ram[46275] = {9'd43,10'd43};
ram[46276] = {9'd47,10'd47};
ram[46277] = {9'd50,10'd50};
ram[46278] = {9'd53,10'd53};
ram[46279] = {9'd56,10'd56};
ram[46280] = {9'd59,10'd59};
ram[46281] = {9'd62,10'd62};
ram[46282] = {9'd65,10'd65};
ram[46283] = {9'd69,10'd69};
ram[46284] = {9'd72,10'd72};
ram[46285] = {9'd75,10'd75};
ram[46286] = {9'd78,10'd78};
ram[46287] = {9'd81,10'd81};
ram[46288] = {9'd84,10'd84};
ram[46289] = {9'd87,10'd87};
ram[46290] = {9'd91,10'd91};
ram[46291] = {9'd94,10'd94};
ram[46292] = {9'd97,10'd97};
ram[46293] = {-9'd100,10'd100};
ram[46294] = {-9'd97,10'd103};
ram[46295] = {-9'd94,10'd106};
ram[46296] = {-9'd91,10'd109};
ram[46297] = {-9'd88,10'd113};
ram[46298] = {-9'd85,10'd116};
ram[46299] = {-9'd81,10'd119};
ram[46300] = {-9'd78,10'd122};
ram[46301] = {-9'd75,10'd125};
ram[46302] = {-9'd72,10'd128};
ram[46303] = {-9'd69,10'd131};
ram[46304] = {-9'd66,10'd135};
ram[46305] = {-9'd63,10'd138};
ram[46306] = {-9'd59,10'd141};
ram[46307] = {-9'd56,10'd144};
ram[46308] = {-9'd53,10'd147};
ram[46309] = {-9'd50,10'd150};
ram[46310] = {-9'd47,10'd153};
ram[46311] = {-9'd44,10'd157};
ram[46312] = {-9'd41,10'd160};
ram[46313] = {-9'd37,10'd163};
ram[46314] = {-9'd34,10'd166};
ram[46315] = {-9'd31,10'd169};
ram[46316] = {-9'd28,10'd172};
ram[46317] = {-9'd25,10'd175};
ram[46318] = {-9'd22,10'd179};
ram[46319] = {-9'd19,10'd182};
ram[46320] = {-9'd15,10'd185};
ram[46321] = {-9'd12,10'd188};
ram[46322] = {-9'd9,10'd191};
ram[46323] = {-9'd6,10'd194};
ram[46324] = {-9'd3,10'd197};
ram[46325] = {9'd0,10'd201};
ram[46326] = {9'd3,10'd204};
ram[46327] = {9'd7,10'd207};
ram[46328] = {9'd10,10'd210};
ram[46329] = {9'd13,10'd213};
ram[46330] = {9'd16,10'd216};
ram[46331] = {9'd19,10'd219};
ram[46332] = {9'd22,10'd223};
ram[46333] = {9'd25,10'd226};
ram[46334] = {9'd29,10'd229};
ram[46335] = {9'd32,10'd232};
ram[46336] = {9'd32,10'd232};
ram[46337] = {9'd35,10'd235};
ram[46338] = {9'd38,10'd238};
ram[46339] = {9'd41,10'd241};
ram[46340] = {9'd44,10'd245};
ram[46341] = {9'd47,10'd248};
ram[46342] = {9'd51,10'd251};
ram[46343] = {9'd54,10'd254};
ram[46344] = {9'd57,10'd257};
ram[46345] = {9'd60,10'd260};
ram[46346] = {9'd63,10'd263};
ram[46347] = {9'd66,10'd267};
ram[46348] = {9'd69,10'd270};
ram[46349] = {9'd73,10'd273};
ram[46350] = {9'd76,10'd276};
ram[46351] = {9'd79,10'd279};
ram[46352] = {9'd82,10'd282};
ram[46353] = {9'd85,10'd285};
ram[46354] = {9'd88,10'd289};
ram[46355] = {9'd91,10'd292};
ram[46356] = {9'd95,10'd295};
ram[46357] = {9'd98,10'd298};
ram[46358] = {-9'd99,10'd301};
ram[46359] = {-9'd96,10'd304};
ram[46360] = {-9'd93,10'd307};
ram[46361] = {-9'd90,10'd311};
ram[46362] = {-9'd87,10'd314};
ram[46363] = {-9'd84,10'd317};
ram[46364] = {-9'd81,10'd320};
ram[46365] = {-9'd77,10'd323};
ram[46366] = {-9'd74,10'd326};
ram[46367] = {-9'd71,10'd329};
ram[46368] = {-9'd68,10'd333};
ram[46369] = {-9'd65,10'd336};
ram[46370] = {-9'd62,10'd339};
ram[46371] = {-9'd59,10'd342};
ram[46372] = {-9'd55,10'd345};
ram[46373] = {-9'd52,10'd348};
ram[46374] = {-9'd49,10'd351};
ram[46375] = {-9'd46,10'd354};
ram[46376] = {-9'd43,10'd358};
ram[46377] = {-9'd40,10'd361};
ram[46378] = {-9'd37,10'd364};
ram[46379] = {-9'd33,10'd367};
ram[46380] = {-9'd30,10'd370};
ram[46381] = {-9'd27,10'd373};
ram[46382] = {-9'd24,10'd376};
ram[46383] = {-9'd21,10'd380};
ram[46384] = {-9'd18,10'd383};
ram[46385] = {-9'd15,10'd386};
ram[46386] = {-9'd11,10'd389};
ram[46387] = {-9'd8,10'd392};
ram[46388] = {-9'd5,10'd395};
ram[46389] = {-9'd2,10'd398};
ram[46390] = {9'd1,-10'd399};
ram[46391] = {9'd4,-10'd396};
ram[46392] = {9'd7,-10'd393};
ram[46393] = {9'd10,-10'd390};
ram[46394] = {9'd14,-10'd387};
ram[46395] = {9'd17,-10'd384};
ram[46396] = {9'd20,-10'd381};
ram[46397] = {9'd23,-10'd377};
ram[46398] = {9'd26,-10'd374};
ram[46399] = {9'd29,-10'd371};
ram[46400] = {9'd32,-10'd368};
ram[46401] = {9'd36,-10'd365};
ram[46402] = {9'd39,-10'd362};
ram[46403] = {9'd42,-10'd359};
ram[46404] = {9'd45,-10'd355};
ram[46405] = {9'd48,-10'd352};
ram[46406] = {9'd51,-10'd349};
ram[46407] = {9'd54,-10'd346};
ram[46408] = {9'd58,-10'd343};
ram[46409] = {9'd61,-10'd340};
ram[46410] = {9'd64,-10'd337};
ram[46411] = {9'd67,-10'd334};
ram[46412] = {9'd70,-10'd330};
ram[46413] = {9'd73,-10'd327};
ram[46414] = {9'd76,-10'd324};
ram[46415] = {9'd80,-10'd321};
ram[46416] = {9'd83,-10'd318};
ram[46417] = {9'd86,-10'd315};
ram[46418] = {9'd89,-10'd312};
ram[46419] = {9'd92,-10'd308};
ram[46420] = {9'd95,-10'd305};
ram[46421] = {9'd98,-10'd302};
ram[46422] = {-9'd99,-10'd299};
ram[46423] = {-9'd96,-10'd296};
ram[46424] = {-9'd92,-10'd293};
ram[46425] = {-9'd89,-10'd290};
ram[46426] = {-9'd86,-10'd286};
ram[46427] = {-9'd83,-10'd283};
ram[46428] = {-9'd80,-10'd280};
ram[46429] = {-9'd77,-10'd277};
ram[46430] = {-9'd74,-10'd274};
ram[46431] = {-9'd70,-10'd271};
ram[46432] = {-9'd67,-10'd268};
ram[46433] = {-9'd64,-10'd264};
ram[46434] = {-9'd61,-10'd261};
ram[46435] = {-9'd58,-10'd258};
ram[46436] = {-9'd55,-10'd255};
ram[46437] = {-9'd52,-10'd252};
ram[46438] = {-9'd48,-10'd249};
ram[46439] = {-9'd45,-10'd246};
ram[46440] = {-9'd42,-10'd242};
ram[46441] = {-9'd39,-10'd239};
ram[46442] = {-9'd36,-10'd236};
ram[46443] = {-9'd33,-10'd233};
ram[46444] = {-9'd30,-10'd230};
ram[46445] = {-9'd26,-10'd227};
ram[46446] = {-9'd23,-10'd224};
ram[46447] = {-9'd20,-10'd220};
ram[46448] = {-9'd17,-10'd217};
ram[46449] = {-9'd14,-10'd214};
ram[46450] = {-9'd11,-10'd211};
ram[46451] = {-9'd8,-10'd208};
ram[46452] = {-9'd4,-10'd205};
ram[46453] = {-9'd1,-10'd202};
ram[46454] = {9'd2,-10'd198};
ram[46455] = {9'd5,-10'd195};
ram[46456] = {9'd8,-10'd192};
ram[46457] = {9'd11,-10'd189};
ram[46458] = {9'd14,-10'd186};
ram[46459] = {9'd18,-10'd183};
ram[46460] = {9'd21,-10'd180};
ram[46461] = {9'd24,-10'd176};
ram[46462] = {9'd27,-10'd173};
ram[46463] = {9'd30,-10'd170};
ram[46464] = {9'd30,-10'd170};
ram[46465] = {9'd33,-10'd167};
ram[46466] = {9'd36,-10'd164};
ram[46467] = {9'd40,-10'd161};
ram[46468] = {9'd43,-10'd158};
ram[46469] = {9'd46,-10'd154};
ram[46470] = {9'd49,-10'd151};
ram[46471] = {9'd52,-10'd148};
ram[46472] = {9'd55,-10'd145};
ram[46473] = {9'd58,-10'd142};
ram[46474] = {9'd62,-10'd139};
ram[46475] = {9'd65,-10'd136};
ram[46476] = {9'd68,-10'd132};
ram[46477] = {9'd71,-10'd129};
ram[46478] = {9'd74,-10'd126};
ram[46479] = {9'd77,-10'd123};
ram[46480] = {9'd80,-10'd120};
ram[46481] = {9'd84,-10'd117};
ram[46482] = {9'd87,-10'd114};
ram[46483] = {9'd90,-10'd110};
ram[46484] = {9'd93,-10'd107};
ram[46485] = {9'd96,-10'd104};
ram[46486] = {9'd99,-10'd101};
ram[46487] = {-9'd98,-10'd98};
ram[46488] = {-9'd95,-10'd95};
ram[46489] = {-9'd92,-10'd92};
ram[46490] = {-9'd88,-10'd88};
ram[46491] = {-9'd85,-10'd85};
ram[46492] = {-9'd82,-10'd82};
ram[46493] = {-9'd79,-10'd79};
ram[46494] = {-9'd76,-10'd76};
ram[46495] = {-9'd73,-10'd73};
ram[46496] = {-9'd70,-10'd70};
ram[46497] = {-9'd66,-10'd66};
ram[46498] = {-9'd63,-10'd63};
ram[46499] = {-9'd60,-10'd60};
ram[46500] = {-9'd57,-10'd57};
ram[46501] = {-9'd54,-10'd54};
ram[46502] = {-9'd51,-10'd51};
ram[46503] = {-9'd48,-10'd48};
ram[46504] = {-9'd44,-10'd44};
ram[46505] = {-9'd41,-10'd41};
ram[46506] = {-9'd38,-10'd38};
ram[46507] = {-9'd35,-10'd35};
ram[46508] = {-9'd32,-10'd32};
ram[46509] = {-9'd29,-10'd29};
ram[46510] = {-9'd26,-10'd26};
ram[46511] = {-9'd22,-10'd22};
ram[46512] = {-9'd19,-10'd19};
ram[46513] = {-9'd16,-10'd16};
ram[46514] = {-9'd13,-10'd13};
ram[46515] = {-9'd10,-10'd10};
ram[46516] = {-9'd7,-10'd7};
ram[46517] = {-9'd4,-10'd4};
ram[46518] = {9'd0,10'd0};
ram[46519] = {9'd3,10'd3};
ram[46520] = {9'd6,10'd6};
ram[46521] = {9'd9,10'd9};
ram[46522] = {9'd12,10'd12};
ram[46523] = {9'd15,10'd15};
ram[46524] = {9'd18,10'd18};
ram[46525] = {9'd21,10'd21};
ram[46526] = {9'd25,10'd25};
ram[46527] = {9'd28,10'd28};
ram[46528] = {9'd31,10'd31};
ram[46529] = {9'd34,10'd34};
ram[46530] = {9'd37,10'd37};
ram[46531] = {9'd40,10'd40};
ram[46532] = {9'd43,10'd43};
ram[46533] = {9'd47,10'd47};
ram[46534] = {9'd50,10'd50};
ram[46535] = {9'd53,10'd53};
ram[46536] = {9'd56,10'd56};
ram[46537] = {9'd59,10'd59};
ram[46538] = {9'd62,10'd62};
ram[46539] = {9'd65,10'd65};
ram[46540] = {9'd69,10'd69};
ram[46541] = {9'd72,10'd72};
ram[46542] = {9'd75,10'd75};
ram[46543] = {9'd78,10'd78};
ram[46544] = {9'd81,10'd81};
ram[46545] = {9'd84,10'd84};
ram[46546] = {9'd87,10'd87};
ram[46547] = {9'd91,10'd91};
ram[46548] = {9'd94,10'd94};
ram[46549] = {9'd97,10'd97};
ram[46550] = {-9'd100,10'd100};
ram[46551] = {-9'd97,10'd103};
ram[46552] = {-9'd94,10'd106};
ram[46553] = {-9'd91,10'd109};
ram[46554] = {-9'd88,10'd113};
ram[46555] = {-9'd85,10'd116};
ram[46556] = {-9'd81,10'd119};
ram[46557] = {-9'd78,10'd122};
ram[46558] = {-9'd75,10'd125};
ram[46559] = {-9'd72,10'd128};
ram[46560] = {-9'd69,10'd131};
ram[46561] = {-9'd66,10'd135};
ram[46562] = {-9'd63,10'd138};
ram[46563] = {-9'd59,10'd141};
ram[46564] = {-9'd56,10'd144};
ram[46565] = {-9'd53,10'd147};
ram[46566] = {-9'd50,10'd150};
ram[46567] = {-9'd47,10'd153};
ram[46568] = {-9'd44,10'd157};
ram[46569] = {-9'd41,10'd160};
ram[46570] = {-9'd37,10'd163};
ram[46571] = {-9'd34,10'd166};
ram[46572] = {-9'd31,10'd169};
ram[46573] = {-9'd28,10'd172};
ram[46574] = {-9'd25,10'd175};
ram[46575] = {-9'd22,10'd179};
ram[46576] = {-9'd19,10'd182};
ram[46577] = {-9'd15,10'd185};
ram[46578] = {-9'd12,10'd188};
ram[46579] = {-9'd9,10'd191};
ram[46580] = {-9'd6,10'd194};
ram[46581] = {-9'd3,10'd197};
ram[46582] = {9'd0,10'd201};
ram[46583] = {9'd3,10'd204};
ram[46584] = {9'd7,10'd207};
ram[46585] = {9'd10,10'd210};
ram[46586] = {9'd13,10'd213};
ram[46587] = {9'd16,10'd216};
ram[46588] = {9'd19,10'd219};
ram[46589] = {9'd22,10'd223};
ram[46590] = {9'd25,10'd226};
ram[46591] = {9'd29,10'd229};
ram[46592] = {9'd29,10'd229};
ram[46593] = {9'd32,10'd232};
ram[46594] = {9'd35,10'd235};
ram[46595] = {9'd38,10'd238};
ram[46596] = {9'd41,10'd241};
ram[46597] = {9'd44,10'd245};
ram[46598] = {9'd47,10'd248};
ram[46599] = {9'd51,10'd251};
ram[46600] = {9'd54,10'd254};
ram[46601] = {9'd57,10'd257};
ram[46602] = {9'd60,10'd260};
ram[46603] = {9'd63,10'd263};
ram[46604] = {9'd66,10'd267};
ram[46605] = {9'd69,10'd270};
ram[46606] = {9'd73,10'd273};
ram[46607] = {9'd76,10'd276};
ram[46608] = {9'd79,10'd279};
ram[46609] = {9'd82,10'd282};
ram[46610] = {9'd85,10'd285};
ram[46611] = {9'd88,10'd289};
ram[46612] = {9'd91,10'd292};
ram[46613] = {9'd95,10'd295};
ram[46614] = {9'd98,10'd298};
ram[46615] = {-9'd99,10'd301};
ram[46616] = {-9'd96,10'd304};
ram[46617] = {-9'd93,10'd307};
ram[46618] = {-9'd90,10'd311};
ram[46619] = {-9'd87,10'd314};
ram[46620] = {-9'd84,10'd317};
ram[46621] = {-9'd81,10'd320};
ram[46622] = {-9'd77,10'd323};
ram[46623] = {-9'd74,10'd326};
ram[46624] = {-9'd71,10'd329};
ram[46625] = {-9'd68,10'd333};
ram[46626] = {-9'd65,10'd336};
ram[46627] = {-9'd62,10'd339};
ram[46628] = {-9'd59,10'd342};
ram[46629] = {-9'd55,10'd345};
ram[46630] = {-9'd52,10'd348};
ram[46631] = {-9'd49,10'd351};
ram[46632] = {-9'd46,10'd354};
ram[46633] = {-9'd43,10'd358};
ram[46634] = {-9'd40,10'd361};
ram[46635] = {-9'd37,10'd364};
ram[46636] = {-9'd33,10'd367};
ram[46637] = {-9'd30,10'd370};
ram[46638] = {-9'd27,10'd373};
ram[46639] = {-9'd24,10'd376};
ram[46640] = {-9'd21,10'd380};
ram[46641] = {-9'd18,10'd383};
ram[46642] = {-9'd15,10'd386};
ram[46643] = {-9'd11,10'd389};
ram[46644] = {-9'd8,10'd392};
ram[46645] = {-9'd5,10'd395};
ram[46646] = {-9'd2,10'd398};
ram[46647] = {9'd1,-10'd399};
ram[46648] = {9'd4,-10'd396};
ram[46649] = {9'd7,-10'd393};
ram[46650] = {9'd10,-10'd390};
ram[46651] = {9'd14,-10'd387};
ram[46652] = {9'd17,-10'd384};
ram[46653] = {9'd20,-10'd381};
ram[46654] = {9'd23,-10'd377};
ram[46655] = {9'd26,-10'd374};
ram[46656] = {9'd29,-10'd371};
ram[46657] = {9'd32,-10'd368};
ram[46658] = {9'd36,-10'd365};
ram[46659] = {9'd39,-10'd362};
ram[46660] = {9'd42,-10'd359};
ram[46661] = {9'd45,-10'd355};
ram[46662] = {9'd48,-10'd352};
ram[46663] = {9'd51,-10'd349};
ram[46664] = {9'd54,-10'd346};
ram[46665] = {9'd58,-10'd343};
ram[46666] = {9'd61,-10'd340};
ram[46667] = {9'd64,-10'd337};
ram[46668] = {9'd67,-10'd334};
ram[46669] = {9'd70,-10'd330};
ram[46670] = {9'd73,-10'd327};
ram[46671] = {9'd76,-10'd324};
ram[46672] = {9'd80,-10'd321};
ram[46673] = {9'd83,-10'd318};
ram[46674] = {9'd86,-10'd315};
ram[46675] = {9'd89,-10'd312};
ram[46676] = {9'd92,-10'd308};
ram[46677] = {9'd95,-10'd305};
ram[46678] = {9'd98,-10'd302};
ram[46679] = {-9'd99,-10'd299};
ram[46680] = {-9'd96,-10'd296};
ram[46681] = {-9'd92,-10'd293};
ram[46682] = {-9'd89,-10'd290};
ram[46683] = {-9'd86,-10'd286};
ram[46684] = {-9'd83,-10'd283};
ram[46685] = {-9'd80,-10'd280};
ram[46686] = {-9'd77,-10'd277};
ram[46687] = {-9'd74,-10'd274};
ram[46688] = {-9'd70,-10'd271};
ram[46689] = {-9'd67,-10'd268};
ram[46690] = {-9'd64,-10'd264};
ram[46691] = {-9'd61,-10'd261};
ram[46692] = {-9'd58,-10'd258};
ram[46693] = {-9'd55,-10'd255};
ram[46694] = {-9'd52,-10'd252};
ram[46695] = {-9'd48,-10'd249};
ram[46696] = {-9'd45,-10'd246};
ram[46697] = {-9'd42,-10'd242};
ram[46698] = {-9'd39,-10'd239};
ram[46699] = {-9'd36,-10'd236};
ram[46700] = {-9'd33,-10'd233};
ram[46701] = {-9'd30,-10'd230};
ram[46702] = {-9'd26,-10'd227};
ram[46703] = {-9'd23,-10'd224};
ram[46704] = {-9'd20,-10'd220};
ram[46705] = {-9'd17,-10'd217};
ram[46706] = {-9'd14,-10'd214};
ram[46707] = {-9'd11,-10'd211};
ram[46708] = {-9'd8,-10'd208};
ram[46709] = {-9'd4,-10'd205};
ram[46710] = {-9'd1,-10'd202};
ram[46711] = {9'd2,-10'd198};
ram[46712] = {9'd5,-10'd195};
ram[46713] = {9'd8,-10'd192};
ram[46714] = {9'd11,-10'd189};
ram[46715] = {9'd14,-10'd186};
ram[46716] = {9'd18,-10'd183};
ram[46717] = {9'd21,-10'd180};
ram[46718] = {9'd24,-10'd176};
ram[46719] = {9'd27,-10'd173};
ram[46720] = {9'd27,-10'd173};
ram[46721] = {9'd30,-10'd170};
ram[46722] = {9'd33,-10'd167};
ram[46723] = {9'd36,-10'd164};
ram[46724] = {9'd40,-10'd161};
ram[46725] = {9'd43,-10'd158};
ram[46726] = {9'd46,-10'd154};
ram[46727] = {9'd49,-10'd151};
ram[46728] = {9'd52,-10'd148};
ram[46729] = {9'd55,-10'd145};
ram[46730] = {9'd58,-10'd142};
ram[46731] = {9'd62,-10'd139};
ram[46732] = {9'd65,-10'd136};
ram[46733] = {9'd68,-10'd132};
ram[46734] = {9'd71,-10'd129};
ram[46735] = {9'd74,-10'd126};
ram[46736] = {9'd77,-10'd123};
ram[46737] = {9'd80,-10'd120};
ram[46738] = {9'd84,-10'd117};
ram[46739] = {9'd87,-10'd114};
ram[46740] = {9'd90,-10'd110};
ram[46741] = {9'd93,-10'd107};
ram[46742] = {9'd96,-10'd104};
ram[46743] = {9'd99,-10'd101};
ram[46744] = {-9'd98,-10'd98};
ram[46745] = {-9'd95,-10'd95};
ram[46746] = {-9'd92,-10'd92};
ram[46747] = {-9'd88,-10'd88};
ram[46748] = {-9'd85,-10'd85};
ram[46749] = {-9'd82,-10'd82};
ram[46750] = {-9'd79,-10'd79};
ram[46751] = {-9'd76,-10'd76};
ram[46752] = {-9'd73,-10'd73};
ram[46753] = {-9'd70,-10'd70};
ram[46754] = {-9'd66,-10'd66};
ram[46755] = {-9'd63,-10'd63};
ram[46756] = {-9'd60,-10'd60};
ram[46757] = {-9'd57,-10'd57};
ram[46758] = {-9'd54,-10'd54};
ram[46759] = {-9'd51,-10'd51};
ram[46760] = {-9'd48,-10'd48};
ram[46761] = {-9'd44,-10'd44};
ram[46762] = {-9'd41,-10'd41};
ram[46763] = {-9'd38,-10'd38};
ram[46764] = {-9'd35,-10'd35};
ram[46765] = {-9'd32,-10'd32};
ram[46766] = {-9'd29,-10'd29};
ram[46767] = {-9'd26,-10'd26};
ram[46768] = {-9'd22,-10'd22};
ram[46769] = {-9'd19,-10'd19};
ram[46770] = {-9'd16,-10'd16};
ram[46771] = {-9'd13,-10'd13};
ram[46772] = {-9'd10,-10'd10};
ram[46773] = {-9'd7,-10'd7};
ram[46774] = {-9'd4,-10'd4};
ram[46775] = {9'd0,10'd0};
ram[46776] = {9'd3,10'd3};
ram[46777] = {9'd6,10'd6};
ram[46778] = {9'd9,10'd9};
ram[46779] = {9'd12,10'd12};
ram[46780] = {9'd15,10'd15};
ram[46781] = {9'd18,10'd18};
ram[46782] = {9'd21,10'd21};
ram[46783] = {9'd25,10'd25};
ram[46784] = {9'd28,10'd28};
ram[46785] = {9'd31,10'd31};
ram[46786] = {9'd34,10'd34};
ram[46787] = {9'd37,10'd37};
ram[46788] = {9'd40,10'd40};
ram[46789] = {9'd43,10'd43};
ram[46790] = {9'd47,10'd47};
ram[46791] = {9'd50,10'd50};
ram[46792] = {9'd53,10'd53};
ram[46793] = {9'd56,10'd56};
ram[46794] = {9'd59,10'd59};
ram[46795] = {9'd62,10'd62};
ram[46796] = {9'd65,10'd65};
ram[46797] = {9'd69,10'd69};
ram[46798] = {9'd72,10'd72};
ram[46799] = {9'd75,10'd75};
ram[46800] = {9'd78,10'd78};
ram[46801] = {9'd81,10'd81};
ram[46802] = {9'd84,10'd84};
ram[46803] = {9'd87,10'd87};
ram[46804] = {9'd91,10'd91};
ram[46805] = {9'd94,10'd94};
ram[46806] = {9'd97,10'd97};
ram[46807] = {-9'd100,10'd100};
ram[46808] = {-9'd97,10'd103};
ram[46809] = {-9'd94,10'd106};
ram[46810] = {-9'd91,10'd109};
ram[46811] = {-9'd88,10'd113};
ram[46812] = {-9'd85,10'd116};
ram[46813] = {-9'd81,10'd119};
ram[46814] = {-9'd78,10'd122};
ram[46815] = {-9'd75,10'd125};
ram[46816] = {-9'd72,10'd128};
ram[46817] = {-9'd69,10'd131};
ram[46818] = {-9'd66,10'd135};
ram[46819] = {-9'd63,10'd138};
ram[46820] = {-9'd59,10'd141};
ram[46821] = {-9'd56,10'd144};
ram[46822] = {-9'd53,10'd147};
ram[46823] = {-9'd50,10'd150};
ram[46824] = {-9'd47,10'd153};
ram[46825] = {-9'd44,10'd157};
ram[46826] = {-9'd41,10'd160};
ram[46827] = {-9'd37,10'd163};
ram[46828] = {-9'd34,10'd166};
ram[46829] = {-9'd31,10'd169};
ram[46830] = {-9'd28,10'd172};
ram[46831] = {-9'd25,10'd175};
ram[46832] = {-9'd22,10'd179};
ram[46833] = {-9'd19,10'd182};
ram[46834] = {-9'd15,10'd185};
ram[46835] = {-9'd12,10'd188};
ram[46836] = {-9'd9,10'd191};
ram[46837] = {-9'd6,10'd194};
ram[46838] = {-9'd3,10'd197};
ram[46839] = {9'd0,10'd201};
ram[46840] = {9'd3,10'd204};
ram[46841] = {9'd7,10'd207};
ram[46842] = {9'd10,10'd210};
ram[46843] = {9'd13,10'd213};
ram[46844] = {9'd16,10'd216};
ram[46845] = {9'd19,10'd219};
ram[46846] = {9'd22,10'd223};
ram[46847] = {9'd25,10'd226};
ram[46848] = {9'd25,10'd226};
ram[46849] = {9'd29,10'd229};
ram[46850] = {9'd32,10'd232};
ram[46851] = {9'd35,10'd235};
ram[46852] = {9'd38,10'd238};
ram[46853] = {9'd41,10'd241};
ram[46854] = {9'd44,10'd245};
ram[46855] = {9'd47,10'd248};
ram[46856] = {9'd51,10'd251};
ram[46857] = {9'd54,10'd254};
ram[46858] = {9'd57,10'd257};
ram[46859] = {9'd60,10'd260};
ram[46860] = {9'd63,10'd263};
ram[46861] = {9'd66,10'd267};
ram[46862] = {9'd69,10'd270};
ram[46863] = {9'd73,10'd273};
ram[46864] = {9'd76,10'd276};
ram[46865] = {9'd79,10'd279};
ram[46866] = {9'd82,10'd282};
ram[46867] = {9'd85,10'd285};
ram[46868] = {9'd88,10'd289};
ram[46869] = {9'd91,10'd292};
ram[46870] = {9'd95,10'd295};
ram[46871] = {9'd98,10'd298};
ram[46872] = {-9'd99,10'd301};
ram[46873] = {-9'd96,10'd304};
ram[46874] = {-9'd93,10'd307};
ram[46875] = {-9'd90,10'd311};
ram[46876] = {-9'd87,10'd314};
ram[46877] = {-9'd84,10'd317};
ram[46878] = {-9'd81,10'd320};
ram[46879] = {-9'd77,10'd323};
ram[46880] = {-9'd74,10'd326};
ram[46881] = {-9'd71,10'd329};
ram[46882] = {-9'd68,10'd333};
ram[46883] = {-9'd65,10'd336};
ram[46884] = {-9'd62,10'd339};
ram[46885] = {-9'd59,10'd342};
ram[46886] = {-9'd55,10'd345};
ram[46887] = {-9'd52,10'd348};
ram[46888] = {-9'd49,10'd351};
ram[46889] = {-9'd46,10'd354};
ram[46890] = {-9'd43,10'd358};
ram[46891] = {-9'd40,10'd361};
ram[46892] = {-9'd37,10'd364};
ram[46893] = {-9'd33,10'd367};
ram[46894] = {-9'd30,10'd370};
ram[46895] = {-9'd27,10'd373};
ram[46896] = {-9'd24,10'd376};
ram[46897] = {-9'd21,10'd380};
ram[46898] = {-9'd18,10'd383};
ram[46899] = {-9'd15,10'd386};
ram[46900] = {-9'd11,10'd389};
ram[46901] = {-9'd8,10'd392};
ram[46902] = {-9'd5,10'd395};
ram[46903] = {-9'd2,10'd398};
ram[46904] = {9'd1,-10'd399};
ram[46905] = {9'd4,-10'd396};
ram[46906] = {9'd7,-10'd393};
ram[46907] = {9'd10,-10'd390};
ram[46908] = {9'd14,-10'd387};
ram[46909] = {9'd17,-10'd384};
ram[46910] = {9'd20,-10'd381};
ram[46911] = {9'd23,-10'd377};
ram[46912] = {9'd26,-10'd374};
ram[46913] = {9'd29,-10'd371};
ram[46914] = {9'd32,-10'd368};
ram[46915] = {9'd36,-10'd365};
ram[46916] = {9'd39,-10'd362};
ram[46917] = {9'd42,-10'd359};
ram[46918] = {9'd45,-10'd355};
ram[46919] = {9'd48,-10'd352};
ram[46920] = {9'd51,-10'd349};
ram[46921] = {9'd54,-10'd346};
ram[46922] = {9'd58,-10'd343};
ram[46923] = {9'd61,-10'd340};
ram[46924] = {9'd64,-10'd337};
ram[46925] = {9'd67,-10'd334};
ram[46926] = {9'd70,-10'd330};
ram[46927] = {9'd73,-10'd327};
ram[46928] = {9'd76,-10'd324};
ram[46929] = {9'd80,-10'd321};
ram[46930] = {9'd83,-10'd318};
ram[46931] = {9'd86,-10'd315};
ram[46932] = {9'd89,-10'd312};
ram[46933] = {9'd92,-10'd308};
ram[46934] = {9'd95,-10'd305};
ram[46935] = {9'd98,-10'd302};
ram[46936] = {-9'd99,-10'd299};
ram[46937] = {-9'd96,-10'd296};
ram[46938] = {-9'd92,-10'd293};
ram[46939] = {-9'd89,-10'd290};
ram[46940] = {-9'd86,-10'd286};
ram[46941] = {-9'd83,-10'd283};
ram[46942] = {-9'd80,-10'd280};
ram[46943] = {-9'd77,-10'd277};
ram[46944] = {-9'd74,-10'd274};
ram[46945] = {-9'd70,-10'd271};
ram[46946] = {-9'd67,-10'd268};
ram[46947] = {-9'd64,-10'd264};
ram[46948] = {-9'd61,-10'd261};
ram[46949] = {-9'd58,-10'd258};
ram[46950] = {-9'd55,-10'd255};
ram[46951] = {-9'd52,-10'd252};
ram[46952] = {-9'd48,-10'd249};
ram[46953] = {-9'd45,-10'd246};
ram[46954] = {-9'd42,-10'd242};
ram[46955] = {-9'd39,-10'd239};
ram[46956] = {-9'd36,-10'd236};
ram[46957] = {-9'd33,-10'd233};
ram[46958] = {-9'd30,-10'd230};
ram[46959] = {-9'd26,-10'd227};
ram[46960] = {-9'd23,-10'd224};
ram[46961] = {-9'd20,-10'd220};
ram[46962] = {-9'd17,-10'd217};
ram[46963] = {-9'd14,-10'd214};
ram[46964] = {-9'd11,-10'd211};
ram[46965] = {-9'd8,-10'd208};
ram[46966] = {-9'd4,-10'd205};
ram[46967] = {-9'd1,-10'd202};
ram[46968] = {9'd2,-10'd198};
ram[46969] = {9'd5,-10'd195};
ram[46970] = {9'd8,-10'd192};
ram[46971] = {9'd11,-10'd189};
ram[46972] = {9'd14,-10'd186};
ram[46973] = {9'd18,-10'd183};
ram[46974] = {9'd21,-10'd180};
ram[46975] = {9'd24,-10'd176};
ram[46976] = {9'd24,-10'd176};
ram[46977] = {9'd27,-10'd173};
ram[46978] = {9'd30,-10'd170};
ram[46979] = {9'd33,-10'd167};
ram[46980] = {9'd36,-10'd164};
ram[46981] = {9'd40,-10'd161};
ram[46982] = {9'd43,-10'd158};
ram[46983] = {9'd46,-10'd154};
ram[46984] = {9'd49,-10'd151};
ram[46985] = {9'd52,-10'd148};
ram[46986] = {9'd55,-10'd145};
ram[46987] = {9'd58,-10'd142};
ram[46988] = {9'd62,-10'd139};
ram[46989] = {9'd65,-10'd136};
ram[46990] = {9'd68,-10'd132};
ram[46991] = {9'd71,-10'd129};
ram[46992] = {9'd74,-10'd126};
ram[46993] = {9'd77,-10'd123};
ram[46994] = {9'd80,-10'd120};
ram[46995] = {9'd84,-10'd117};
ram[46996] = {9'd87,-10'd114};
ram[46997] = {9'd90,-10'd110};
ram[46998] = {9'd93,-10'd107};
ram[46999] = {9'd96,-10'd104};
ram[47000] = {9'd99,-10'd101};
ram[47001] = {-9'd98,-10'd98};
ram[47002] = {-9'd95,-10'd95};
ram[47003] = {-9'd92,-10'd92};
ram[47004] = {-9'd88,-10'd88};
ram[47005] = {-9'd85,-10'd85};
ram[47006] = {-9'd82,-10'd82};
ram[47007] = {-9'd79,-10'd79};
ram[47008] = {-9'd76,-10'd76};
ram[47009] = {-9'd73,-10'd73};
ram[47010] = {-9'd70,-10'd70};
ram[47011] = {-9'd66,-10'd66};
ram[47012] = {-9'd63,-10'd63};
ram[47013] = {-9'd60,-10'd60};
ram[47014] = {-9'd57,-10'd57};
ram[47015] = {-9'd54,-10'd54};
ram[47016] = {-9'd51,-10'd51};
ram[47017] = {-9'd48,-10'd48};
ram[47018] = {-9'd44,-10'd44};
ram[47019] = {-9'd41,-10'd41};
ram[47020] = {-9'd38,-10'd38};
ram[47021] = {-9'd35,-10'd35};
ram[47022] = {-9'd32,-10'd32};
ram[47023] = {-9'd29,-10'd29};
ram[47024] = {-9'd26,-10'd26};
ram[47025] = {-9'd22,-10'd22};
ram[47026] = {-9'd19,-10'd19};
ram[47027] = {-9'd16,-10'd16};
ram[47028] = {-9'd13,-10'd13};
ram[47029] = {-9'd10,-10'd10};
ram[47030] = {-9'd7,-10'd7};
ram[47031] = {-9'd4,-10'd4};
ram[47032] = {9'd0,10'd0};
ram[47033] = {9'd3,10'd3};
ram[47034] = {9'd6,10'd6};
ram[47035] = {9'd9,10'd9};
ram[47036] = {9'd12,10'd12};
ram[47037] = {9'd15,10'd15};
ram[47038] = {9'd18,10'd18};
ram[47039] = {9'd21,10'd21};
ram[47040] = {9'd25,10'd25};
ram[47041] = {9'd28,10'd28};
ram[47042] = {9'd31,10'd31};
ram[47043] = {9'd34,10'd34};
ram[47044] = {9'd37,10'd37};
ram[47045] = {9'd40,10'd40};
ram[47046] = {9'd43,10'd43};
ram[47047] = {9'd47,10'd47};
ram[47048] = {9'd50,10'd50};
ram[47049] = {9'd53,10'd53};
ram[47050] = {9'd56,10'd56};
ram[47051] = {9'd59,10'd59};
ram[47052] = {9'd62,10'd62};
ram[47053] = {9'd65,10'd65};
ram[47054] = {9'd69,10'd69};
ram[47055] = {9'd72,10'd72};
ram[47056] = {9'd75,10'd75};
ram[47057] = {9'd78,10'd78};
ram[47058] = {9'd81,10'd81};
ram[47059] = {9'd84,10'd84};
ram[47060] = {9'd87,10'd87};
ram[47061] = {9'd91,10'd91};
ram[47062] = {9'd94,10'd94};
ram[47063] = {9'd97,10'd97};
ram[47064] = {-9'd100,10'd100};
ram[47065] = {-9'd97,10'd103};
ram[47066] = {-9'd94,10'd106};
ram[47067] = {-9'd91,10'd109};
ram[47068] = {-9'd88,10'd113};
ram[47069] = {-9'd85,10'd116};
ram[47070] = {-9'd81,10'd119};
ram[47071] = {-9'd78,10'd122};
ram[47072] = {-9'd75,10'd125};
ram[47073] = {-9'd72,10'd128};
ram[47074] = {-9'd69,10'd131};
ram[47075] = {-9'd66,10'd135};
ram[47076] = {-9'd63,10'd138};
ram[47077] = {-9'd59,10'd141};
ram[47078] = {-9'd56,10'd144};
ram[47079] = {-9'd53,10'd147};
ram[47080] = {-9'd50,10'd150};
ram[47081] = {-9'd47,10'd153};
ram[47082] = {-9'd44,10'd157};
ram[47083] = {-9'd41,10'd160};
ram[47084] = {-9'd37,10'd163};
ram[47085] = {-9'd34,10'd166};
ram[47086] = {-9'd31,10'd169};
ram[47087] = {-9'd28,10'd172};
ram[47088] = {-9'd25,10'd175};
ram[47089] = {-9'd22,10'd179};
ram[47090] = {-9'd19,10'd182};
ram[47091] = {-9'd15,10'd185};
ram[47092] = {-9'd12,10'd188};
ram[47093] = {-9'd9,10'd191};
ram[47094] = {-9'd6,10'd194};
ram[47095] = {-9'd3,10'd197};
ram[47096] = {9'd0,10'd201};
ram[47097] = {9'd3,10'd204};
ram[47098] = {9'd7,10'd207};
ram[47099] = {9'd10,10'd210};
ram[47100] = {9'd13,10'd213};
ram[47101] = {9'd16,10'd216};
ram[47102] = {9'd19,10'd219};
ram[47103] = {9'd22,10'd223};
ram[47104] = {9'd22,10'd223};
ram[47105] = {9'd25,10'd226};
ram[47106] = {9'd29,10'd229};
ram[47107] = {9'd32,10'd232};
ram[47108] = {9'd35,10'd235};
ram[47109] = {9'd38,10'd238};
ram[47110] = {9'd41,10'd241};
ram[47111] = {9'd44,10'd245};
ram[47112] = {9'd47,10'd248};
ram[47113] = {9'd51,10'd251};
ram[47114] = {9'd54,10'd254};
ram[47115] = {9'd57,10'd257};
ram[47116] = {9'd60,10'd260};
ram[47117] = {9'd63,10'd263};
ram[47118] = {9'd66,10'd267};
ram[47119] = {9'd69,10'd270};
ram[47120] = {9'd73,10'd273};
ram[47121] = {9'd76,10'd276};
ram[47122] = {9'd79,10'd279};
ram[47123] = {9'd82,10'd282};
ram[47124] = {9'd85,10'd285};
ram[47125] = {9'd88,10'd289};
ram[47126] = {9'd91,10'd292};
ram[47127] = {9'd95,10'd295};
ram[47128] = {9'd98,10'd298};
ram[47129] = {-9'd99,10'd301};
ram[47130] = {-9'd96,10'd304};
ram[47131] = {-9'd93,10'd307};
ram[47132] = {-9'd90,10'd311};
ram[47133] = {-9'd87,10'd314};
ram[47134] = {-9'd84,10'd317};
ram[47135] = {-9'd81,10'd320};
ram[47136] = {-9'd77,10'd323};
ram[47137] = {-9'd74,10'd326};
ram[47138] = {-9'd71,10'd329};
ram[47139] = {-9'd68,10'd333};
ram[47140] = {-9'd65,10'd336};
ram[47141] = {-9'd62,10'd339};
ram[47142] = {-9'd59,10'd342};
ram[47143] = {-9'd55,10'd345};
ram[47144] = {-9'd52,10'd348};
ram[47145] = {-9'd49,10'd351};
ram[47146] = {-9'd46,10'd354};
ram[47147] = {-9'd43,10'd358};
ram[47148] = {-9'd40,10'd361};
ram[47149] = {-9'd37,10'd364};
ram[47150] = {-9'd33,10'd367};
ram[47151] = {-9'd30,10'd370};
ram[47152] = {-9'd27,10'd373};
ram[47153] = {-9'd24,10'd376};
ram[47154] = {-9'd21,10'd380};
ram[47155] = {-9'd18,10'd383};
ram[47156] = {-9'd15,10'd386};
ram[47157] = {-9'd11,10'd389};
ram[47158] = {-9'd8,10'd392};
ram[47159] = {-9'd5,10'd395};
ram[47160] = {-9'd2,10'd398};
ram[47161] = {9'd1,-10'd399};
ram[47162] = {9'd4,-10'd396};
ram[47163] = {9'd7,-10'd393};
ram[47164] = {9'd10,-10'd390};
ram[47165] = {9'd14,-10'd387};
ram[47166] = {9'd17,-10'd384};
ram[47167] = {9'd20,-10'd381};
ram[47168] = {9'd23,-10'd377};
ram[47169] = {9'd26,-10'd374};
ram[47170] = {9'd29,-10'd371};
ram[47171] = {9'd32,-10'd368};
ram[47172] = {9'd36,-10'd365};
ram[47173] = {9'd39,-10'd362};
ram[47174] = {9'd42,-10'd359};
ram[47175] = {9'd45,-10'd355};
ram[47176] = {9'd48,-10'd352};
ram[47177] = {9'd51,-10'd349};
ram[47178] = {9'd54,-10'd346};
ram[47179] = {9'd58,-10'd343};
ram[47180] = {9'd61,-10'd340};
ram[47181] = {9'd64,-10'd337};
ram[47182] = {9'd67,-10'd334};
ram[47183] = {9'd70,-10'd330};
ram[47184] = {9'd73,-10'd327};
ram[47185] = {9'd76,-10'd324};
ram[47186] = {9'd80,-10'd321};
ram[47187] = {9'd83,-10'd318};
ram[47188] = {9'd86,-10'd315};
ram[47189] = {9'd89,-10'd312};
ram[47190] = {9'd92,-10'd308};
ram[47191] = {9'd95,-10'd305};
ram[47192] = {9'd98,-10'd302};
ram[47193] = {-9'd99,-10'd299};
ram[47194] = {-9'd96,-10'd296};
ram[47195] = {-9'd92,-10'd293};
ram[47196] = {-9'd89,-10'd290};
ram[47197] = {-9'd86,-10'd286};
ram[47198] = {-9'd83,-10'd283};
ram[47199] = {-9'd80,-10'd280};
ram[47200] = {-9'd77,-10'd277};
ram[47201] = {-9'd74,-10'd274};
ram[47202] = {-9'd70,-10'd271};
ram[47203] = {-9'd67,-10'd268};
ram[47204] = {-9'd64,-10'd264};
ram[47205] = {-9'd61,-10'd261};
ram[47206] = {-9'd58,-10'd258};
ram[47207] = {-9'd55,-10'd255};
ram[47208] = {-9'd52,-10'd252};
ram[47209] = {-9'd48,-10'd249};
ram[47210] = {-9'd45,-10'd246};
ram[47211] = {-9'd42,-10'd242};
ram[47212] = {-9'd39,-10'd239};
ram[47213] = {-9'd36,-10'd236};
ram[47214] = {-9'd33,-10'd233};
ram[47215] = {-9'd30,-10'd230};
ram[47216] = {-9'd26,-10'd227};
ram[47217] = {-9'd23,-10'd224};
ram[47218] = {-9'd20,-10'd220};
ram[47219] = {-9'd17,-10'd217};
ram[47220] = {-9'd14,-10'd214};
ram[47221] = {-9'd11,-10'd211};
ram[47222] = {-9'd8,-10'd208};
ram[47223] = {-9'd4,-10'd205};
ram[47224] = {-9'd1,-10'd202};
ram[47225] = {9'd2,-10'd198};
ram[47226] = {9'd5,-10'd195};
ram[47227] = {9'd8,-10'd192};
ram[47228] = {9'd11,-10'd189};
ram[47229] = {9'd14,-10'd186};
ram[47230] = {9'd18,-10'd183};
ram[47231] = {9'd21,-10'd180};
ram[47232] = {9'd21,-10'd180};
ram[47233] = {9'd24,-10'd176};
ram[47234] = {9'd27,-10'd173};
ram[47235] = {9'd30,-10'd170};
ram[47236] = {9'd33,-10'd167};
ram[47237] = {9'd36,-10'd164};
ram[47238] = {9'd40,-10'd161};
ram[47239] = {9'd43,-10'd158};
ram[47240] = {9'd46,-10'd154};
ram[47241] = {9'd49,-10'd151};
ram[47242] = {9'd52,-10'd148};
ram[47243] = {9'd55,-10'd145};
ram[47244] = {9'd58,-10'd142};
ram[47245] = {9'd62,-10'd139};
ram[47246] = {9'd65,-10'd136};
ram[47247] = {9'd68,-10'd132};
ram[47248] = {9'd71,-10'd129};
ram[47249] = {9'd74,-10'd126};
ram[47250] = {9'd77,-10'd123};
ram[47251] = {9'd80,-10'd120};
ram[47252] = {9'd84,-10'd117};
ram[47253] = {9'd87,-10'd114};
ram[47254] = {9'd90,-10'd110};
ram[47255] = {9'd93,-10'd107};
ram[47256] = {9'd96,-10'd104};
ram[47257] = {9'd99,-10'd101};
ram[47258] = {-9'd98,-10'd98};
ram[47259] = {-9'd95,-10'd95};
ram[47260] = {-9'd92,-10'd92};
ram[47261] = {-9'd88,-10'd88};
ram[47262] = {-9'd85,-10'd85};
ram[47263] = {-9'd82,-10'd82};
ram[47264] = {-9'd79,-10'd79};
ram[47265] = {-9'd76,-10'd76};
ram[47266] = {-9'd73,-10'd73};
ram[47267] = {-9'd70,-10'd70};
ram[47268] = {-9'd66,-10'd66};
ram[47269] = {-9'd63,-10'd63};
ram[47270] = {-9'd60,-10'd60};
ram[47271] = {-9'd57,-10'd57};
ram[47272] = {-9'd54,-10'd54};
ram[47273] = {-9'd51,-10'd51};
ram[47274] = {-9'd48,-10'd48};
ram[47275] = {-9'd44,-10'd44};
ram[47276] = {-9'd41,-10'd41};
ram[47277] = {-9'd38,-10'd38};
ram[47278] = {-9'd35,-10'd35};
ram[47279] = {-9'd32,-10'd32};
ram[47280] = {-9'd29,-10'd29};
ram[47281] = {-9'd26,-10'd26};
ram[47282] = {-9'd22,-10'd22};
ram[47283] = {-9'd19,-10'd19};
ram[47284] = {-9'd16,-10'd16};
ram[47285] = {-9'd13,-10'd13};
ram[47286] = {-9'd10,-10'd10};
ram[47287] = {-9'd7,-10'd7};
ram[47288] = {-9'd4,-10'd4};
ram[47289] = {9'd0,10'd0};
ram[47290] = {9'd3,10'd3};
ram[47291] = {9'd6,10'd6};
ram[47292] = {9'd9,10'd9};
ram[47293] = {9'd12,10'd12};
ram[47294] = {9'd15,10'd15};
ram[47295] = {9'd18,10'd18};
ram[47296] = {9'd21,10'd21};
ram[47297] = {9'd25,10'd25};
ram[47298] = {9'd28,10'd28};
ram[47299] = {9'd31,10'd31};
ram[47300] = {9'd34,10'd34};
ram[47301] = {9'd37,10'd37};
ram[47302] = {9'd40,10'd40};
ram[47303] = {9'd43,10'd43};
ram[47304] = {9'd47,10'd47};
ram[47305] = {9'd50,10'd50};
ram[47306] = {9'd53,10'd53};
ram[47307] = {9'd56,10'd56};
ram[47308] = {9'd59,10'd59};
ram[47309] = {9'd62,10'd62};
ram[47310] = {9'd65,10'd65};
ram[47311] = {9'd69,10'd69};
ram[47312] = {9'd72,10'd72};
ram[47313] = {9'd75,10'd75};
ram[47314] = {9'd78,10'd78};
ram[47315] = {9'd81,10'd81};
ram[47316] = {9'd84,10'd84};
ram[47317] = {9'd87,10'd87};
ram[47318] = {9'd91,10'd91};
ram[47319] = {9'd94,10'd94};
ram[47320] = {9'd97,10'd97};
ram[47321] = {-9'd100,10'd100};
ram[47322] = {-9'd97,10'd103};
ram[47323] = {-9'd94,10'd106};
ram[47324] = {-9'd91,10'd109};
ram[47325] = {-9'd88,10'd113};
ram[47326] = {-9'd85,10'd116};
ram[47327] = {-9'd81,10'd119};
ram[47328] = {-9'd78,10'd122};
ram[47329] = {-9'd75,10'd125};
ram[47330] = {-9'd72,10'd128};
ram[47331] = {-9'd69,10'd131};
ram[47332] = {-9'd66,10'd135};
ram[47333] = {-9'd63,10'd138};
ram[47334] = {-9'd59,10'd141};
ram[47335] = {-9'd56,10'd144};
ram[47336] = {-9'd53,10'd147};
ram[47337] = {-9'd50,10'd150};
ram[47338] = {-9'd47,10'd153};
ram[47339] = {-9'd44,10'd157};
ram[47340] = {-9'd41,10'd160};
ram[47341] = {-9'd37,10'd163};
ram[47342] = {-9'd34,10'd166};
ram[47343] = {-9'd31,10'd169};
ram[47344] = {-9'd28,10'd172};
ram[47345] = {-9'd25,10'd175};
ram[47346] = {-9'd22,10'd179};
ram[47347] = {-9'd19,10'd182};
ram[47348] = {-9'd15,10'd185};
ram[47349] = {-9'd12,10'd188};
ram[47350] = {-9'd9,10'd191};
ram[47351] = {-9'd6,10'd194};
ram[47352] = {-9'd3,10'd197};
ram[47353] = {9'd0,10'd201};
ram[47354] = {9'd3,10'd204};
ram[47355] = {9'd7,10'd207};
ram[47356] = {9'd10,10'd210};
ram[47357] = {9'd13,10'd213};
ram[47358] = {9'd16,10'd216};
ram[47359] = {9'd19,10'd219};
ram[47360] = {9'd19,10'd219};
ram[47361] = {9'd22,10'd223};
ram[47362] = {9'd25,10'd226};
ram[47363] = {9'd29,10'd229};
ram[47364] = {9'd32,10'd232};
ram[47365] = {9'd35,10'd235};
ram[47366] = {9'd38,10'd238};
ram[47367] = {9'd41,10'd241};
ram[47368] = {9'd44,10'd245};
ram[47369] = {9'd47,10'd248};
ram[47370] = {9'd51,10'd251};
ram[47371] = {9'd54,10'd254};
ram[47372] = {9'd57,10'd257};
ram[47373] = {9'd60,10'd260};
ram[47374] = {9'd63,10'd263};
ram[47375] = {9'd66,10'd267};
ram[47376] = {9'd69,10'd270};
ram[47377] = {9'd73,10'd273};
ram[47378] = {9'd76,10'd276};
ram[47379] = {9'd79,10'd279};
ram[47380] = {9'd82,10'd282};
ram[47381] = {9'd85,10'd285};
ram[47382] = {9'd88,10'd289};
ram[47383] = {9'd91,10'd292};
ram[47384] = {9'd95,10'd295};
ram[47385] = {9'd98,10'd298};
ram[47386] = {-9'd99,10'd301};
ram[47387] = {-9'd96,10'd304};
ram[47388] = {-9'd93,10'd307};
ram[47389] = {-9'd90,10'd311};
ram[47390] = {-9'd87,10'd314};
ram[47391] = {-9'd84,10'd317};
ram[47392] = {-9'd81,10'd320};
ram[47393] = {-9'd77,10'd323};
ram[47394] = {-9'd74,10'd326};
ram[47395] = {-9'd71,10'd329};
ram[47396] = {-9'd68,10'd333};
ram[47397] = {-9'd65,10'd336};
ram[47398] = {-9'd62,10'd339};
ram[47399] = {-9'd59,10'd342};
ram[47400] = {-9'd55,10'd345};
ram[47401] = {-9'd52,10'd348};
ram[47402] = {-9'd49,10'd351};
ram[47403] = {-9'd46,10'd354};
ram[47404] = {-9'd43,10'd358};
ram[47405] = {-9'd40,10'd361};
ram[47406] = {-9'd37,10'd364};
ram[47407] = {-9'd33,10'd367};
ram[47408] = {-9'd30,10'd370};
ram[47409] = {-9'd27,10'd373};
ram[47410] = {-9'd24,10'd376};
ram[47411] = {-9'd21,10'd380};
ram[47412] = {-9'd18,10'd383};
ram[47413] = {-9'd15,10'd386};
ram[47414] = {-9'd11,10'd389};
ram[47415] = {-9'd8,10'd392};
ram[47416] = {-9'd5,10'd395};
ram[47417] = {-9'd2,10'd398};
ram[47418] = {9'd1,-10'd399};
ram[47419] = {9'd4,-10'd396};
ram[47420] = {9'd7,-10'd393};
ram[47421] = {9'd10,-10'd390};
ram[47422] = {9'd14,-10'd387};
ram[47423] = {9'd17,-10'd384};
ram[47424] = {9'd20,-10'd381};
ram[47425] = {9'd23,-10'd377};
ram[47426] = {9'd26,-10'd374};
ram[47427] = {9'd29,-10'd371};
ram[47428] = {9'd32,-10'd368};
ram[47429] = {9'd36,-10'd365};
ram[47430] = {9'd39,-10'd362};
ram[47431] = {9'd42,-10'd359};
ram[47432] = {9'd45,-10'd355};
ram[47433] = {9'd48,-10'd352};
ram[47434] = {9'd51,-10'd349};
ram[47435] = {9'd54,-10'd346};
ram[47436] = {9'd58,-10'd343};
ram[47437] = {9'd61,-10'd340};
ram[47438] = {9'd64,-10'd337};
ram[47439] = {9'd67,-10'd334};
ram[47440] = {9'd70,-10'd330};
ram[47441] = {9'd73,-10'd327};
ram[47442] = {9'd76,-10'd324};
ram[47443] = {9'd80,-10'd321};
ram[47444] = {9'd83,-10'd318};
ram[47445] = {9'd86,-10'd315};
ram[47446] = {9'd89,-10'd312};
ram[47447] = {9'd92,-10'd308};
ram[47448] = {9'd95,-10'd305};
ram[47449] = {9'd98,-10'd302};
ram[47450] = {-9'd99,-10'd299};
ram[47451] = {-9'd96,-10'd296};
ram[47452] = {-9'd92,-10'd293};
ram[47453] = {-9'd89,-10'd290};
ram[47454] = {-9'd86,-10'd286};
ram[47455] = {-9'd83,-10'd283};
ram[47456] = {-9'd80,-10'd280};
ram[47457] = {-9'd77,-10'd277};
ram[47458] = {-9'd74,-10'd274};
ram[47459] = {-9'd70,-10'd271};
ram[47460] = {-9'd67,-10'd268};
ram[47461] = {-9'd64,-10'd264};
ram[47462] = {-9'd61,-10'd261};
ram[47463] = {-9'd58,-10'd258};
ram[47464] = {-9'd55,-10'd255};
ram[47465] = {-9'd52,-10'd252};
ram[47466] = {-9'd48,-10'd249};
ram[47467] = {-9'd45,-10'd246};
ram[47468] = {-9'd42,-10'd242};
ram[47469] = {-9'd39,-10'd239};
ram[47470] = {-9'd36,-10'd236};
ram[47471] = {-9'd33,-10'd233};
ram[47472] = {-9'd30,-10'd230};
ram[47473] = {-9'd26,-10'd227};
ram[47474] = {-9'd23,-10'd224};
ram[47475] = {-9'd20,-10'd220};
ram[47476] = {-9'd17,-10'd217};
ram[47477] = {-9'd14,-10'd214};
ram[47478] = {-9'd11,-10'd211};
ram[47479] = {-9'd8,-10'd208};
ram[47480] = {-9'd4,-10'd205};
ram[47481] = {-9'd1,-10'd202};
ram[47482] = {9'd2,-10'd198};
ram[47483] = {9'd5,-10'd195};
ram[47484] = {9'd8,-10'd192};
ram[47485] = {9'd11,-10'd189};
ram[47486] = {9'd14,-10'd186};
ram[47487] = {9'd18,-10'd183};
ram[47488] = {9'd18,-10'd183};
ram[47489] = {9'd21,-10'd180};
ram[47490] = {9'd24,-10'd176};
ram[47491] = {9'd27,-10'd173};
ram[47492] = {9'd30,-10'd170};
ram[47493] = {9'd33,-10'd167};
ram[47494] = {9'd36,-10'd164};
ram[47495] = {9'd40,-10'd161};
ram[47496] = {9'd43,-10'd158};
ram[47497] = {9'd46,-10'd154};
ram[47498] = {9'd49,-10'd151};
ram[47499] = {9'd52,-10'd148};
ram[47500] = {9'd55,-10'd145};
ram[47501] = {9'd58,-10'd142};
ram[47502] = {9'd62,-10'd139};
ram[47503] = {9'd65,-10'd136};
ram[47504] = {9'd68,-10'd132};
ram[47505] = {9'd71,-10'd129};
ram[47506] = {9'd74,-10'd126};
ram[47507] = {9'd77,-10'd123};
ram[47508] = {9'd80,-10'd120};
ram[47509] = {9'd84,-10'd117};
ram[47510] = {9'd87,-10'd114};
ram[47511] = {9'd90,-10'd110};
ram[47512] = {9'd93,-10'd107};
ram[47513] = {9'd96,-10'd104};
ram[47514] = {9'd99,-10'd101};
ram[47515] = {-9'd98,-10'd98};
ram[47516] = {-9'd95,-10'd95};
ram[47517] = {-9'd92,-10'd92};
ram[47518] = {-9'd88,-10'd88};
ram[47519] = {-9'd85,-10'd85};
ram[47520] = {-9'd82,-10'd82};
ram[47521] = {-9'd79,-10'd79};
ram[47522] = {-9'd76,-10'd76};
ram[47523] = {-9'd73,-10'd73};
ram[47524] = {-9'd70,-10'd70};
ram[47525] = {-9'd66,-10'd66};
ram[47526] = {-9'd63,-10'd63};
ram[47527] = {-9'd60,-10'd60};
ram[47528] = {-9'd57,-10'd57};
ram[47529] = {-9'd54,-10'd54};
ram[47530] = {-9'd51,-10'd51};
ram[47531] = {-9'd48,-10'd48};
ram[47532] = {-9'd44,-10'd44};
ram[47533] = {-9'd41,-10'd41};
ram[47534] = {-9'd38,-10'd38};
ram[47535] = {-9'd35,-10'd35};
ram[47536] = {-9'd32,-10'd32};
ram[47537] = {-9'd29,-10'd29};
ram[47538] = {-9'd26,-10'd26};
ram[47539] = {-9'd22,-10'd22};
ram[47540] = {-9'd19,-10'd19};
ram[47541] = {-9'd16,-10'd16};
ram[47542] = {-9'd13,-10'd13};
ram[47543] = {-9'd10,-10'd10};
ram[47544] = {-9'd7,-10'd7};
ram[47545] = {-9'd4,-10'd4};
ram[47546] = {9'd0,10'd0};
ram[47547] = {9'd3,10'd3};
ram[47548] = {9'd6,10'd6};
ram[47549] = {9'd9,10'd9};
ram[47550] = {9'd12,10'd12};
ram[47551] = {9'd15,10'd15};
ram[47552] = {9'd18,10'd18};
ram[47553] = {9'd21,10'd21};
ram[47554] = {9'd25,10'd25};
ram[47555] = {9'd28,10'd28};
ram[47556] = {9'd31,10'd31};
ram[47557] = {9'd34,10'd34};
ram[47558] = {9'd37,10'd37};
ram[47559] = {9'd40,10'd40};
ram[47560] = {9'd43,10'd43};
ram[47561] = {9'd47,10'd47};
ram[47562] = {9'd50,10'd50};
ram[47563] = {9'd53,10'd53};
ram[47564] = {9'd56,10'd56};
ram[47565] = {9'd59,10'd59};
ram[47566] = {9'd62,10'd62};
ram[47567] = {9'd65,10'd65};
ram[47568] = {9'd69,10'd69};
ram[47569] = {9'd72,10'd72};
ram[47570] = {9'd75,10'd75};
ram[47571] = {9'd78,10'd78};
ram[47572] = {9'd81,10'd81};
ram[47573] = {9'd84,10'd84};
ram[47574] = {9'd87,10'd87};
ram[47575] = {9'd91,10'd91};
ram[47576] = {9'd94,10'd94};
ram[47577] = {9'd97,10'd97};
ram[47578] = {-9'd100,10'd100};
ram[47579] = {-9'd97,10'd103};
ram[47580] = {-9'd94,10'd106};
ram[47581] = {-9'd91,10'd109};
ram[47582] = {-9'd88,10'd113};
ram[47583] = {-9'd85,10'd116};
ram[47584] = {-9'd81,10'd119};
ram[47585] = {-9'd78,10'd122};
ram[47586] = {-9'd75,10'd125};
ram[47587] = {-9'd72,10'd128};
ram[47588] = {-9'd69,10'd131};
ram[47589] = {-9'd66,10'd135};
ram[47590] = {-9'd63,10'd138};
ram[47591] = {-9'd59,10'd141};
ram[47592] = {-9'd56,10'd144};
ram[47593] = {-9'd53,10'd147};
ram[47594] = {-9'd50,10'd150};
ram[47595] = {-9'd47,10'd153};
ram[47596] = {-9'd44,10'd157};
ram[47597] = {-9'd41,10'd160};
ram[47598] = {-9'd37,10'd163};
ram[47599] = {-9'd34,10'd166};
ram[47600] = {-9'd31,10'd169};
ram[47601] = {-9'd28,10'd172};
ram[47602] = {-9'd25,10'd175};
ram[47603] = {-9'd22,10'd179};
ram[47604] = {-9'd19,10'd182};
ram[47605] = {-9'd15,10'd185};
ram[47606] = {-9'd12,10'd188};
ram[47607] = {-9'd9,10'd191};
ram[47608] = {-9'd6,10'd194};
ram[47609] = {-9'd3,10'd197};
ram[47610] = {9'd0,10'd201};
ram[47611] = {9'd3,10'd204};
ram[47612] = {9'd7,10'd207};
ram[47613] = {9'd10,10'd210};
ram[47614] = {9'd13,10'd213};
ram[47615] = {9'd16,10'd216};
ram[47616] = {9'd16,10'd216};
ram[47617] = {9'd19,10'd219};
ram[47618] = {9'd22,10'd223};
ram[47619] = {9'd25,10'd226};
ram[47620] = {9'd29,10'd229};
ram[47621] = {9'd32,10'd232};
ram[47622] = {9'd35,10'd235};
ram[47623] = {9'd38,10'd238};
ram[47624] = {9'd41,10'd241};
ram[47625] = {9'd44,10'd245};
ram[47626] = {9'd47,10'd248};
ram[47627] = {9'd51,10'd251};
ram[47628] = {9'd54,10'd254};
ram[47629] = {9'd57,10'd257};
ram[47630] = {9'd60,10'd260};
ram[47631] = {9'd63,10'd263};
ram[47632] = {9'd66,10'd267};
ram[47633] = {9'd69,10'd270};
ram[47634] = {9'd73,10'd273};
ram[47635] = {9'd76,10'd276};
ram[47636] = {9'd79,10'd279};
ram[47637] = {9'd82,10'd282};
ram[47638] = {9'd85,10'd285};
ram[47639] = {9'd88,10'd289};
ram[47640] = {9'd91,10'd292};
ram[47641] = {9'd95,10'd295};
ram[47642] = {9'd98,10'd298};
ram[47643] = {-9'd99,10'd301};
ram[47644] = {-9'd96,10'd304};
ram[47645] = {-9'd93,10'd307};
ram[47646] = {-9'd90,10'd311};
ram[47647] = {-9'd87,10'd314};
ram[47648] = {-9'd84,10'd317};
ram[47649] = {-9'd81,10'd320};
ram[47650] = {-9'd77,10'd323};
ram[47651] = {-9'd74,10'd326};
ram[47652] = {-9'd71,10'd329};
ram[47653] = {-9'd68,10'd333};
ram[47654] = {-9'd65,10'd336};
ram[47655] = {-9'd62,10'd339};
ram[47656] = {-9'd59,10'd342};
ram[47657] = {-9'd55,10'd345};
ram[47658] = {-9'd52,10'd348};
ram[47659] = {-9'd49,10'd351};
ram[47660] = {-9'd46,10'd354};
ram[47661] = {-9'd43,10'd358};
ram[47662] = {-9'd40,10'd361};
ram[47663] = {-9'd37,10'd364};
ram[47664] = {-9'd33,10'd367};
ram[47665] = {-9'd30,10'd370};
ram[47666] = {-9'd27,10'd373};
ram[47667] = {-9'd24,10'd376};
ram[47668] = {-9'd21,10'd380};
ram[47669] = {-9'd18,10'd383};
ram[47670] = {-9'd15,10'd386};
ram[47671] = {-9'd11,10'd389};
ram[47672] = {-9'd8,10'd392};
ram[47673] = {-9'd5,10'd395};
ram[47674] = {-9'd2,10'd398};
ram[47675] = {9'd1,-10'd399};
ram[47676] = {9'd4,-10'd396};
ram[47677] = {9'd7,-10'd393};
ram[47678] = {9'd10,-10'd390};
ram[47679] = {9'd14,-10'd387};
ram[47680] = {9'd17,-10'd384};
ram[47681] = {9'd20,-10'd381};
ram[47682] = {9'd23,-10'd377};
ram[47683] = {9'd26,-10'd374};
ram[47684] = {9'd29,-10'd371};
ram[47685] = {9'd32,-10'd368};
ram[47686] = {9'd36,-10'd365};
ram[47687] = {9'd39,-10'd362};
ram[47688] = {9'd42,-10'd359};
ram[47689] = {9'd45,-10'd355};
ram[47690] = {9'd48,-10'd352};
ram[47691] = {9'd51,-10'd349};
ram[47692] = {9'd54,-10'd346};
ram[47693] = {9'd58,-10'd343};
ram[47694] = {9'd61,-10'd340};
ram[47695] = {9'd64,-10'd337};
ram[47696] = {9'd67,-10'd334};
ram[47697] = {9'd70,-10'd330};
ram[47698] = {9'd73,-10'd327};
ram[47699] = {9'd76,-10'd324};
ram[47700] = {9'd80,-10'd321};
ram[47701] = {9'd83,-10'd318};
ram[47702] = {9'd86,-10'd315};
ram[47703] = {9'd89,-10'd312};
ram[47704] = {9'd92,-10'd308};
ram[47705] = {9'd95,-10'd305};
ram[47706] = {9'd98,-10'd302};
ram[47707] = {-9'd99,-10'd299};
ram[47708] = {-9'd96,-10'd296};
ram[47709] = {-9'd92,-10'd293};
ram[47710] = {-9'd89,-10'd290};
ram[47711] = {-9'd86,-10'd286};
ram[47712] = {-9'd83,-10'd283};
ram[47713] = {-9'd80,-10'd280};
ram[47714] = {-9'd77,-10'd277};
ram[47715] = {-9'd74,-10'd274};
ram[47716] = {-9'd70,-10'd271};
ram[47717] = {-9'd67,-10'd268};
ram[47718] = {-9'd64,-10'd264};
ram[47719] = {-9'd61,-10'd261};
ram[47720] = {-9'd58,-10'd258};
ram[47721] = {-9'd55,-10'd255};
ram[47722] = {-9'd52,-10'd252};
ram[47723] = {-9'd48,-10'd249};
ram[47724] = {-9'd45,-10'd246};
ram[47725] = {-9'd42,-10'd242};
ram[47726] = {-9'd39,-10'd239};
ram[47727] = {-9'd36,-10'd236};
ram[47728] = {-9'd33,-10'd233};
ram[47729] = {-9'd30,-10'd230};
ram[47730] = {-9'd26,-10'd227};
ram[47731] = {-9'd23,-10'd224};
ram[47732] = {-9'd20,-10'd220};
ram[47733] = {-9'd17,-10'd217};
ram[47734] = {-9'd14,-10'd214};
ram[47735] = {-9'd11,-10'd211};
ram[47736] = {-9'd8,-10'd208};
ram[47737] = {-9'd4,-10'd205};
ram[47738] = {-9'd1,-10'd202};
ram[47739] = {9'd2,-10'd198};
ram[47740] = {9'd5,-10'd195};
ram[47741] = {9'd8,-10'd192};
ram[47742] = {9'd11,-10'd189};
ram[47743] = {9'd14,-10'd186};
ram[47744] = {9'd14,-10'd186};
ram[47745] = {9'd18,-10'd183};
ram[47746] = {9'd21,-10'd180};
ram[47747] = {9'd24,-10'd176};
ram[47748] = {9'd27,-10'd173};
ram[47749] = {9'd30,-10'd170};
ram[47750] = {9'd33,-10'd167};
ram[47751] = {9'd36,-10'd164};
ram[47752] = {9'd40,-10'd161};
ram[47753] = {9'd43,-10'd158};
ram[47754] = {9'd46,-10'd154};
ram[47755] = {9'd49,-10'd151};
ram[47756] = {9'd52,-10'd148};
ram[47757] = {9'd55,-10'd145};
ram[47758] = {9'd58,-10'd142};
ram[47759] = {9'd62,-10'd139};
ram[47760] = {9'd65,-10'd136};
ram[47761] = {9'd68,-10'd132};
ram[47762] = {9'd71,-10'd129};
ram[47763] = {9'd74,-10'd126};
ram[47764] = {9'd77,-10'd123};
ram[47765] = {9'd80,-10'd120};
ram[47766] = {9'd84,-10'd117};
ram[47767] = {9'd87,-10'd114};
ram[47768] = {9'd90,-10'd110};
ram[47769] = {9'd93,-10'd107};
ram[47770] = {9'd96,-10'd104};
ram[47771] = {9'd99,-10'd101};
ram[47772] = {-9'd98,-10'd98};
ram[47773] = {-9'd95,-10'd95};
ram[47774] = {-9'd92,-10'd92};
ram[47775] = {-9'd88,-10'd88};
ram[47776] = {-9'd85,-10'd85};
ram[47777] = {-9'd82,-10'd82};
ram[47778] = {-9'd79,-10'd79};
ram[47779] = {-9'd76,-10'd76};
ram[47780] = {-9'd73,-10'd73};
ram[47781] = {-9'd70,-10'd70};
ram[47782] = {-9'd66,-10'd66};
ram[47783] = {-9'd63,-10'd63};
ram[47784] = {-9'd60,-10'd60};
ram[47785] = {-9'd57,-10'd57};
ram[47786] = {-9'd54,-10'd54};
ram[47787] = {-9'd51,-10'd51};
ram[47788] = {-9'd48,-10'd48};
ram[47789] = {-9'd44,-10'd44};
ram[47790] = {-9'd41,-10'd41};
ram[47791] = {-9'd38,-10'd38};
ram[47792] = {-9'd35,-10'd35};
ram[47793] = {-9'd32,-10'd32};
ram[47794] = {-9'd29,-10'd29};
ram[47795] = {-9'd26,-10'd26};
ram[47796] = {-9'd22,-10'd22};
ram[47797] = {-9'd19,-10'd19};
ram[47798] = {-9'd16,-10'd16};
ram[47799] = {-9'd13,-10'd13};
ram[47800] = {-9'd10,-10'd10};
ram[47801] = {-9'd7,-10'd7};
ram[47802] = {-9'd4,-10'd4};
ram[47803] = {9'd0,10'd0};
ram[47804] = {9'd3,10'd3};
ram[47805] = {9'd6,10'd6};
ram[47806] = {9'd9,10'd9};
ram[47807] = {9'd12,10'd12};
ram[47808] = {9'd15,10'd15};
ram[47809] = {9'd18,10'd18};
ram[47810] = {9'd21,10'd21};
ram[47811] = {9'd25,10'd25};
ram[47812] = {9'd28,10'd28};
ram[47813] = {9'd31,10'd31};
ram[47814] = {9'd34,10'd34};
ram[47815] = {9'd37,10'd37};
ram[47816] = {9'd40,10'd40};
ram[47817] = {9'd43,10'd43};
ram[47818] = {9'd47,10'd47};
ram[47819] = {9'd50,10'd50};
ram[47820] = {9'd53,10'd53};
ram[47821] = {9'd56,10'd56};
ram[47822] = {9'd59,10'd59};
ram[47823] = {9'd62,10'd62};
ram[47824] = {9'd65,10'd65};
ram[47825] = {9'd69,10'd69};
ram[47826] = {9'd72,10'd72};
ram[47827] = {9'd75,10'd75};
ram[47828] = {9'd78,10'd78};
ram[47829] = {9'd81,10'd81};
ram[47830] = {9'd84,10'd84};
ram[47831] = {9'd87,10'd87};
ram[47832] = {9'd91,10'd91};
ram[47833] = {9'd94,10'd94};
ram[47834] = {9'd97,10'd97};
ram[47835] = {-9'd100,10'd100};
ram[47836] = {-9'd97,10'd103};
ram[47837] = {-9'd94,10'd106};
ram[47838] = {-9'd91,10'd109};
ram[47839] = {-9'd88,10'd113};
ram[47840] = {-9'd85,10'd116};
ram[47841] = {-9'd81,10'd119};
ram[47842] = {-9'd78,10'd122};
ram[47843] = {-9'd75,10'd125};
ram[47844] = {-9'd72,10'd128};
ram[47845] = {-9'd69,10'd131};
ram[47846] = {-9'd66,10'd135};
ram[47847] = {-9'd63,10'd138};
ram[47848] = {-9'd59,10'd141};
ram[47849] = {-9'd56,10'd144};
ram[47850] = {-9'd53,10'd147};
ram[47851] = {-9'd50,10'd150};
ram[47852] = {-9'd47,10'd153};
ram[47853] = {-9'd44,10'd157};
ram[47854] = {-9'd41,10'd160};
ram[47855] = {-9'd37,10'd163};
ram[47856] = {-9'd34,10'd166};
ram[47857] = {-9'd31,10'd169};
ram[47858] = {-9'd28,10'd172};
ram[47859] = {-9'd25,10'd175};
ram[47860] = {-9'd22,10'd179};
ram[47861] = {-9'd19,10'd182};
ram[47862] = {-9'd15,10'd185};
ram[47863] = {-9'd12,10'd188};
ram[47864] = {-9'd9,10'd191};
ram[47865] = {-9'd6,10'd194};
ram[47866] = {-9'd3,10'd197};
ram[47867] = {9'd0,10'd201};
ram[47868] = {9'd3,10'd204};
ram[47869] = {9'd7,10'd207};
ram[47870] = {9'd10,10'd210};
ram[47871] = {9'd13,10'd213};
ram[47872] = {9'd13,10'd213};
ram[47873] = {9'd16,10'd216};
ram[47874] = {9'd19,10'd219};
ram[47875] = {9'd22,10'd223};
ram[47876] = {9'd25,10'd226};
ram[47877] = {9'd29,10'd229};
ram[47878] = {9'd32,10'd232};
ram[47879] = {9'd35,10'd235};
ram[47880] = {9'd38,10'd238};
ram[47881] = {9'd41,10'd241};
ram[47882] = {9'd44,10'd245};
ram[47883] = {9'd47,10'd248};
ram[47884] = {9'd51,10'd251};
ram[47885] = {9'd54,10'd254};
ram[47886] = {9'd57,10'd257};
ram[47887] = {9'd60,10'd260};
ram[47888] = {9'd63,10'd263};
ram[47889] = {9'd66,10'd267};
ram[47890] = {9'd69,10'd270};
ram[47891] = {9'd73,10'd273};
ram[47892] = {9'd76,10'd276};
ram[47893] = {9'd79,10'd279};
ram[47894] = {9'd82,10'd282};
ram[47895] = {9'd85,10'd285};
ram[47896] = {9'd88,10'd289};
ram[47897] = {9'd91,10'd292};
ram[47898] = {9'd95,10'd295};
ram[47899] = {9'd98,10'd298};
ram[47900] = {-9'd99,10'd301};
ram[47901] = {-9'd96,10'd304};
ram[47902] = {-9'd93,10'd307};
ram[47903] = {-9'd90,10'd311};
ram[47904] = {-9'd87,10'd314};
ram[47905] = {-9'd84,10'd317};
ram[47906] = {-9'd81,10'd320};
ram[47907] = {-9'd77,10'd323};
ram[47908] = {-9'd74,10'd326};
ram[47909] = {-9'd71,10'd329};
ram[47910] = {-9'd68,10'd333};
ram[47911] = {-9'd65,10'd336};
ram[47912] = {-9'd62,10'd339};
ram[47913] = {-9'd59,10'd342};
ram[47914] = {-9'd55,10'd345};
ram[47915] = {-9'd52,10'd348};
ram[47916] = {-9'd49,10'd351};
ram[47917] = {-9'd46,10'd354};
ram[47918] = {-9'd43,10'd358};
ram[47919] = {-9'd40,10'd361};
ram[47920] = {-9'd37,10'd364};
ram[47921] = {-9'd33,10'd367};
ram[47922] = {-9'd30,10'd370};
ram[47923] = {-9'd27,10'd373};
ram[47924] = {-9'd24,10'd376};
ram[47925] = {-9'd21,10'd380};
ram[47926] = {-9'd18,10'd383};
ram[47927] = {-9'd15,10'd386};
ram[47928] = {-9'd11,10'd389};
ram[47929] = {-9'd8,10'd392};
ram[47930] = {-9'd5,10'd395};
ram[47931] = {-9'd2,10'd398};
ram[47932] = {9'd1,-10'd399};
ram[47933] = {9'd4,-10'd396};
ram[47934] = {9'd7,-10'd393};
ram[47935] = {9'd10,-10'd390};
ram[47936] = {9'd14,-10'd387};
ram[47937] = {9'd17,-10'd384};
ram[47938] = {9'd20,-10'd381};
ram[47939] = {9'd23,-10'd377};
ram[47940] = {9'd26,-10'd374};
ram[47941] = {9'd29,-10'd371};
ram[47942] = {9'd32,-10'd368};
ram[47943] = {9'd36,-10'd365};
ram[47944] = {9'd39,-10'd362};
ram[47945] = {9'd42,-10'd359};
ram[47946] = {9'd45,-10'd355};
ram[47947] = {9'd48,-10'd352};
ram[47948] = {9'd51,-10'd349};
ram[47949] = {9'd54,-10'd346};
ram[47950] = {9'd58,-10'd343};
ram[47951] = {9'd61,-10'd340};
ram[47952] = {9'd64,-10'd337};
ram[47953] = {9'd67,-10'd334};
ram[47954] = {9'd70,-10'd330};
ram[47955] = {9'd73,-10'd327};
ram[47956] = {9'd76,-10'd324};
ram[47957] = {9'd80,-10'd321};
ram[47958] = {9'd83,-10'd318};
ram[47959] = {9'd86,-10'd315};
ram[47960] = {9'd89,-10'd312};
ram[47961] = {9'd92,-10'd308};
ram[47962] = {9'd95,-10'd305};
ram[47963] = {9'd98,-10'd302};
ram[47964] = {-9'd99,-10'd299};
ram[47965] = {-9'd96,-10'd296};
ram[47966] = {-9'd92,-10'd293};
ram[47967] = {-9'd89,-10'd290};
ram[47968] = {-9'd86,-10'd286};
ram[47969] = {-9'd83,-10'd283};
ram[47970] = {-9'd80,-10'd280};
ram[47971] = {-9'd77,-10'd277};
ram[47972] = {-9'd74,-10'd274};
ram[47973] = {-9'd70,-10'd271};
ram[47974] = {-9'd67,-10'd268};
ram[47975] = {-9'd64,-10'd264};
ram[47976] = {-9'd61,-10'd261};
ram[47977] = {-9'd58,-10'd258};
ram[47978] = {-9'd55,-10'd255};
ram[47979] = {-9'd52,-10'd252};
ram[47980] = {-9'd48,-10'd249};
ram[47981] = {-9'd45,-10'd246};
ram[47982] = {-9'd42,-10'd242};
ram[47983] = {-9'd39,-10'd239};
ram[47984] = {-9'd36,-10'd236};
ram[47985] = {-9'd33,-10'd233};
ram[47986] = {-9'd30,-10'd230};
ram[47987] = {-9'd26,-10'd227};
ram[47988] = {-9'd23,-10'd224};
ram[47989] = {-9'd20,-10'd220};
ram[47990] = {-9'd17,-10'd217};
ram[47991] = {-9'd14,-10'd214};
ram[47992] = {-9'd11,-10'd211};
ram[47993] = {-9'd8,-10'd208};
ram[47994] = {-9'd4,-10'd205};
ram[47995] = {-9'd1,-10'd202};
ram[47996] = {9'd2,-10'd198};
ram[47997] = {9'd5,-10'd195};
ram[47998] = {9'd8,-10'd192};
ram[47999] = {9'd11,-10'd189};
ram[48000] = {9'd11,-10'd189};
ram[48001] = {9'd14,-10'd186};
ram[48002] = {9'd18,-10'd183};
ram[48003] = {9'd21,-10'd180};
ram[48004] = {9'd24,-10'd176};
ram[48005] = {9'd27,-10'd173};
ram[48006] = {9'd30,-10'd170};
ram[48007] = {9'd33,-10'd167};
ram[48008] = {9'd36,-10'd164};
ram[48009] = {9'd40,-10'd161};
ram[48010] = {9'd43,-10'd158};
ram[48011] = {9'd46,-10'd154};
ram[48012] = {9'd49,-10'd151};
ram[48013] = {9'd52,-10'd148};
ram[48014] = {9'd55,-10'd145};
ram[48015] = {9'd58,-10'd142};
ram[48016] = {9'd62,-10'd139};
ram[48017] = {9'd65,-10'd136};
ram[48018] = {9'd68,-10'd132};
ram[48019] = {9'd71,-10'd129};
ram[48020] = {9'd74,-10'd126};
ram[48021] = {9'd77,-10'd123};
ram[48022] = {9'd80,-10'd120};
ram[48023] = {9'd84,-10'd117};
ram[48024] = {9'd87,-10'd114};
ram[48025] = {9'd90,-10'd110};
ram[48026] = {9'd93,-10'd107};
ram[48027] = {9'd96,-10'd104};
ram[48028] = {9'd99,-10'd101};
ram[48029] = {-9'd98,-10'd98};
ram[48030] = {-9'd95,-10'd95};
ram[48031] = {-9'd92,-10'd92};
ram[48032] = {-9'd88,-10'd88};
ram[48033] = {-9'd85,-10'd85};
ram[48034] = {-9'd82,-10'd82};
ram[48035] = {-9'd79,-10'd79};
ram[48036] = {-9'd76,-10'd76};
ram[48037] = {-9'd73,-10'd73};
ram[48038] = {-9'd70,-10'd70};
ram[48039] = {-9'd66,-10'd66};
ram[48040] = {-9'd63,-10'd63};
ram[48041] = {-9'd60,-10'd60};
ram[48042] = {-9'd57,-10'd57};
ram[48043] = {-9'd54,-10'd54};
ram[48044] = {-9'd51,-10'd51};
ram[48045] = {-9'd48,-10'd48};
ram[48046] = {-9'd44,-10'd44};
ram[48047] = {-9'd41,-10'd41};
ram[48048] = {-9'd38,-10'd38};
ram[48049] = {-9'd35,-10'd35};
ram[48050] = {-9'd32,-10'd32};
ram[48051] = {-9'd29,-10'd29};
ram[48052] = {-9'd26,-10'd26};
ram[48053] = {-9'd22,-10'd22};
ram[48054] = {-9'd19,-10'd19};
ram[48055] = {-9'd16,-10'd16};
ram[48056] = {-9'd13,-10'd13};
ram[48057] = {-9'd10,-10'd10};
ram[48058] = {-9'd7,-10'd7};
ram[48059] = {-9'd4,-10'd4};
ram[48060] = {9'd0,10'd0};
ram[48061] = {9'd3,10'd3};
ram[48062] = {9'd6,10'd6};
ram[48063] = {9'd9,10'd9};
ram[48064] = {9'd12,10'd12};
ram[48065] = {9'd15,10'd15};
ram[48066] = {9'd18,10'd18};
ram[48067] = {9'd21,10'd21};
ram[48068] = {9'd25,10'd25};
ram[48069] = {9'd28,10'd28};
ram[48070] = {9'd31,10'd31};
ram[48071] = {9'd34,10'd34};
ram[48072] = {9'd37,10'd37};
ram[48073] = {9'd40,10'd40};
ram[48074] = {9'd43,10'd43};
ram[48075] = {9'd47,10'd47};
ram[48076] = {9'd50,10'd50};
ram[48077] = {9'd53,10'd53};
ram[48078] = {9'd56,10'd56};
ram[48079] = {9'd59,10'd59};
ram[48080] = {9'd62,10'd62};
ram[48081] = {9'd65,10'd65};
ram[48082] = {9'd69,10'd69};
ram[48083] = {9'd72,10'd72};
ram[48084] = {9'd75,10'd75};
ram[48085] = {9'd78,10'd78};
ram[48086] = {9'd81,10'd81};
ram[48087] = {9'd84,10'd84};
ram[48088] = {9'd87,10'd87};
ram[48089] = {9'd91,10'd91};
ram[48090] = {9'd94,10'd94};
ram[48091] = {9'd97,10'd97};
ram[48092] = {-9'd100,10'd100};
ram[48093] = {-9'd97,10'd103};
ram[48094] = {-9'd94,10'd106};
ram[48095] = {-9'd91,10'd109};
ram[48096] = {-9'd88,10'd113};
ram[48097] = {-9'd85,10'd116};
ram[48098] = {-9'd81,10'd119};
ram[48099] = {-9'd78,10'd122};
ram[48100] = {-9'd75,10'd125};
ram[48101] = {-9'd72,10'd128};
ram[48102] = {-9'd69,10'd131};
ram[48103] = {-9'd66,10'd135};
ram[48104] = {-9'd63,10'd138};
ram[48105] = {-9'd59,10'd141};
ram[48106] = {-9'd56,10'd144};
ram[48107] = {-9'd53,10'd147};
ram[48108] = {-9'd50,10'd150};
ram[48109] = {-9'd47,10'd153};
ram[48110] = {-9'd44,10'd157};
ram[48111] = {-9'd41,10'd160};
ram[48112] = {-9'd37,10'd163};
ram[48113] = {-9'd34,10'd166};
ram[48114] = {-9'd31,10'd169};
ram[48115] = {-9'd28,10'd172};
ram[48116] = {-9'd25,10'd175};
ram[48117] = {-9'd22,10'd179};
ram[48118] = {-9'd19,10'd182};
ram[48119] = {-9'd15,10'd185};
ram[48120] = {-9'd12,10'd188};
ram[48121] = {-9'd9,10'd191};
ram[48122] = {-9'd6,10'd194};
ram[48123] = {-9'd3,10'd197};
ram[48124] = {9'd0,10'd201};
ram[48125] = {9'd3,10'd204};
ram[48126] = {9'd7,10'd207};
ram[48127] = {9'd10,10'd210};
ram[48128] = {9'd10,10'd210};
ram[48129] = {9'd13,10'd213};
ram[48130] = {9'd16,10'd216};
ram[48131] = {9'd19,10'd219};
ram[48132] = {9'd22,10'd223};
ram[48133] = {9'd25,10'd226};
ram[48134] = {9'd29,10'd229};
ram[48135] = {9'd32,10'd232};
ram[48136] = {9'd35,10'd235};
ram[48137] = {9'd38,10'd238};
ram[48138] = {9'd41,10'd241};
ram[48139] = {9'd44,10'd245};
ram[48140] = {9'd47,10'd248};
ram[48141] = {9'd51,10'd251};
ram[48142] = {9'd54,10'd254};
ram[48143] = {9'd57,10'd257};
ram[48144] = {9'd60,10'd260};
ram[48145] = {9'd63,10'd263};
ram[48146] = {9'd66,10'd267};
ram[48147] = {9'd69,10'd270};
ram[48148] = {9'd73,10'd273};
ram[48149] = {9'd76,10'd276};
ram[48150] = {9'd79,10'd279};
ram[48151] = {9'd82,10'd282};
ram[48152] = {9'd85,10'd285};
ram[48153] = {9'd88,10'd289};
ram[48154] = {9'd91,10'd292};
ram[48155] = {9'd95,10'd295};
ram[48156] = {9'd98,10'd298};
ram[48157] = {-9'd99,10'd301};
ram[48158] = {-9'd96,10'd304};
ram[48159] = {-9'd93,10'd307};
ram[48160] = {-9'd90,10'd311};
ram[48161] = {-9'd87,10'd314};
ram[48162] = {-9'd84,10'd317};
ram[48163] = {-9'd81,10'd320};
ram[48164] = {-9'd77,10'd323};
ram[48165] = {-9'd74,10'd326};
ram[48166] = {-9'd71,10'd329};
ram[48167] = {-9'd68,10'd333};
ram[48168] = {-9'd65,10'd336};
ram[48169] = {-9'd62,10'd339};
ram[48170] = {-9'd59,10'd342};
ram[48171] = {-9'd55,10'd345};
ram[48172] = {-9'd52,10'd348};
ram[48173] = {-9'd49,10'd351};
ram[48174] = {-9'd46,10'd354};
ram[48175] = {-9'd43,10'd358};
ram[48176] = {-9'd40,10'd361};
ram[48177] = {-9'd37,10'd364};
ram[48178] = {-9'd33,10'd367};
ram[48179] = {-9'd30,10'd370};
ram[48180] = {-9'd27,10'd373};
ram[48181] = {-9'd24,10'd376};
ram[48182] = {-9'd21,10'd380};
ram[48183] = {-9'd18,10'd383};
ram[48184] = {-9'd15,10'd386};
ram[48185] = {-9'd11,10'd389};
ram[48186] = {-9'd8,10'd392};
ram[48187] = {-9'd5,10'd395};
ram[48188] = {-9'd2,10'd398};
ram[48189] = {9'd1,-10'd399};
ram[48190] = {9'd4,-10'd396};
ram[48191] = {9'd7,-10'd393};
ram[48192] = {9'd10,-10'd390};
ram[48193] = {9'd14,-10'd387};
ram[48194] = {9'd17,-10'd384};
ram[48195] = {9'd20,-10'd381};
ram[48196] = {9'd23,-10'd377};
ram[48197] = {9'd26,-10'd374};
ram[48198] = {9'd29,-10'd371};
ram[48199] = {9'd32,-10'd368};
ram[48200] = {9'd36,-10'd365};
ram[48201] = {9'd39,-10'd362};
ram[48202] = {9'd42,-10'd359};
ram[48203] = {9'd45,-10'd355};
ram[48204] = {9'd48,-10'd352};
ram[48205] = {9'd51,-10'd349};
ram[48206] = {9'd54,-10'd346};
ram[48207] = {9'd58,-10'd343};
ram[48208] = {9'd61,-10'd340};
ram[48209] = {9'd64,-10'd337};
ram[48210] = {9'd67,-10'd334};
ram[48211] = {9'd70,-10'd330};
ram[48212] = {9'd73,-10'd327};
ram[48213] = {9'd76,-10'd324};
ram[48214] = {9'd80,-10'd321};
ram[48215] = {9'd83,-10'd318};
ram[48216] = {9'd86,-10'd315};
ram[48217] = {9'd89,-10'd312};
ram[48218] = {9'd92,-10'd308};
ram[48219] = {9'd95,-10'd305};
ram[48220] = {9'd98,-10'd302};
ram[48221] = {-9'd99,-10'd299};
ram[48222] = {-9'd96,-10'd296};
ram[48223] = {-9'd92,-10'd293};
ram[48224] = {-9'd89,-10'd290};
ram[48225] = {-9'd86,-10'd286};
ram[48226] = {-9'd83,-10'd283};
ram[48227] = {-9'd80,-10'd280};
ram[48228] = {-9'd77,-10'd277};
ram[48229] = {-9'd74,-10'd274};
ram[48230] = {-9'd70,-10'd271};
ram[48231] = {-9'd67,-10'd268};
ram[48232] = {-9'd64,-10'd264};
ram[48233] = {-9'd61,-10'd261};
ram[48234] = {-9'd58,-10'd258};
ram[48235] = {-9'd55,-10'd255};
ram[48236] = {-9'd52,-10'd252};
ram[48237] = {-9'd48,-10'd249};
ram[48238] = {-9'd45,-10'd246};
ram[48239] = {-9'd42,-10'd242};
ram[48240] = {-9'd39,-10'd239};
ram[48241] = {-9'd36,-10'd236};
ram[48242] = {-9'd33,-10'd233};
ram[48243] = {-9'd30,-10'd230};
ram[48244] = {-9'd26,-10'd227};
ram[48245] = {-9'd23,-10'd224};
ram[48246] = {-9'd20,-10'd220};
ram[48247] = {-9'd17,-10'd217};
ram[48248] = {-9'd14,-10'd214};
ram[48249] = {-9'd11,-10'd211};
ram[48250] = {-9'd8,-10'd208};
ram[48251] = {-9'd4,-10'd205};
ram[48252] = {-9'd1,-10'd202};
ram[48253] = {9'd2,-10'd198};
ram[48254] = {9'd5,-10'd195};
ram[48255] = {9'd8,-10'd192};
ram[48256] = {9'd8,-10'd192};
ram[48257] = {9'd11,-10'd189};
ram[48258] = {9'd14,-10'd186};
ram[48259] = {9'd18,-10'd183};
ram[48260] = {9'd21,-10'd180};
ram[48261] = {9'd24,-10'd176};
ram[48262] = {9'd27,-10'd173};
ram[48263] = {9'd30,-10'd170};
ram[48264] = {9'd33,-10'd167};
ram[48265] = {9'd36,-10'd164};
ram[48266] = {9'd40,-10'd161};
ram[48267] = {9'd43,-10'd158};
ram[48268] = {9'd46,-10'd154};
ram[48269] = {9'd49,-10'd151};
ram[48270] = {9'd52,-10'd148};
ram[48271] = {9'd55,-10'd145};
ram[48272] = {9'd58,-10'd142};
ram[48273] = {9'd62,-10'd139};
ram[48274] = {9'd65,-10'd136};
ram[48275] = {9'd68,-10'd132};
ram[48276] = {9'd71,-10'd129};
ram[48277] = {9'd74,-10'd126};
ram[48278] = {9'd77,-10'd123};
ram[48279] = {9'd80,-10'd120};
ram[48280] = {9'd84,-10'd117};
ram[48281] = {9'd87,-10'd114};
ram[48282] = {9'd90,-10'd110};
ram[48283] = {9'd93,-10'd107};
ram[48284] = {9'd96,-10'd104};
ram[48285] = {9'd99,-10'd101};
ram[48286] = {-9'd98,-10'd98};
ram[48287] = {-9'd95,-10'd95};
ram[48288] = {-9'd92,-10'd92};
ram[48289] = {-9'd88,-10'd88};
ram[48290] = {-9'd85,-10'd85};
ram[48291] = {-9'd82,-10'd82};
ram[48292] = {-9'd79,-10'd79};
ram[48293] = {-9'd76,-10'd76};
ram[48294] = {-9'd73,-10'd73};
ram[48295] = {-9'd70,-10'd70};
ram[48296] = {-9'd66,-10'd66};
ram[48297] = {-9'd63,-10'd63};
ram[48298] = {-9'd60,-10'd60};
ram[48299] = {-9'd57,-10'd57};
ram[48300] = {-9'd54,-10'd54};
ram[48301] = {-9'd51,-10'd51};
ram[48302] = {-9'd48,-10'd48};
ram[48303] = {-9'd44,-10'd44};
ram[48304] = {-9'd41,-10'd41};
ram[48305] = {-9'd38,-10'd38};
ram[48306] = {-9'd35,-10'd35};
ram[48307] = {-9'd32,-10'd32};
ram[48308] = {-9'd29,-10'd29};
ram[48309] = {-9'd26,-10'd26};
ram[48310] = {-9'd22,-10'd22};
ram[48311] = {-9'd19,-10'd19};
ram[48312] = {-9'd16,-10'd16};
ram[48313] = {-9'd13,-10'd13};
ram[48314] = {-9'd10,-10'd10};
ram[48315] = {-9'd7,-10'd7};
ram[48316] = {-9'd4,-10'd4};
ram[48317] = {9'd0,10'd0};
ram[48318] = {9'd3,10'd3};
ram[48319] = {9'd6,10'd6};
ram[48320] = {9'd9,10'd9};
ram[48321] = {9'd12,10'd12};
ram[48322] = {9'd15,10'd15};
ram[48323] = {9'd18,10'd18};
ram[48324] = {9'd21,10'd21};
ram[48325] = {9'd25,10'd25};
ram[48326] = {9'd28,10'd28};
ram[48327] = {9'd31,10'd31};
ram[48328] = {9'd34,10'd34};
ram[48329] = {9'd37,10'd37};
ram[48330] = {9'd40,10'd40};
ram[48331] = {9'd43,10'd43};
ram[48332] = {9'd47,10'd47};
ram[48333] = {9'd50,10'd50};
ram[48334] = {9'd53,10'd53};
ram[48335] = {9'd56,10'd56};
ram[48336] = {9'd59,10'd59};
ram[48337] = {9'd62,10'd62};
ram[48338] = {9'd65,10'd65};
ram[48339] = {9'd69,10'd69};
ram[48340] = {9'd72,10'd72};
ram[48341] = {9'd75,10'd75};
ram[48342] = {9'd78,10'd78};
ram[48343] = {9'd81,10'd81};
ram[48344] = {9'd84,10'd84};
ram[48345] = {9'd87,10'd87};
ram[48346] = {9'd91,10'd91};
ram[48347] = {9'd94,10'd94};
ram[48348] = {9'd97,10'd97};
ram[48349] = {-9'd100,10'd100};
ram[48350] = {-9'd97,10'd103};
ram[48351] = {-9'd94,10'd106};
ram[48352] = {-9'd91,10'd109};
ram[48353] = {-9'd88,10'd113};
ram[48354] = {-9'd85,10'd116};
ram[48355] = {-9'd81,10'd119};
ram[48356] = {-9'd78,10'd122};
ram[48357] = {-9'd75,10'd125};
ram[48358] = {-9'd72,10'd128};
ram[48359] = {-9'd69,10'd131};
ram[48360] = {-9'd66,10'd135};
ram[48361] = {-9'd63,10'd138};
ram[48362] = {-9'd59,10'd141};
ram[48363] = {-9'd56,10'd144};
ram[48364] = {-9'd53,10'd147};
ram[48365] = {-9'd50,10'd150};
ram[48366] = {-9'd47,10'd153};
ram[48367] = {-9'd44,10'd157};
ram[48368] = {-9'd41,10'd160};
ram[48369] = {-9'd37,10'd163};
ram[48370] = {-9'd34,10'd166};
ram[48371] = {-9'd31,10'd169};
ram[48372] = {-9'd28,10'd172};
ram[48373] = {-9'd25,10'd175};
ram[48374] = {-9'd22,10'd179};
ram[48375] = {-9'd19,10'd182};
ram[48376] = {-9'd15,10'd185};
ram[48377] = {-9'd12,10'd188};
ram[48378] = {-9'd9,10'd191};
ram[48379] = {-9'd6,10'd194};
ram[48380] = {-9'd3,10'd197};
ram[48381] = {9'd0,10'd201};
ram[48382] = {9'd3,10'd204};
ram[48383] = {9'd7,10'd207};
ram[48384] = {9'd7,10'd207};
ram[48385] = {9'd10,10'd210};
ram[48386] = {9'd13,10'd213};
ram[48387] = {9'd16,10'd216};
ram[48388] = {9'd19,10'd219};
ram[48389] = {9'd22,10'd223};
ram[48390] = {9'd25,10'd226};
ram[48391] = {9'd29,10'd229};
ram[48392] = {9'd32,10'd232};
ram[48393] = {9'd35,10'd235};
ram[48394] = {9'd38,10'd238};
ram[48395] = {9'd41,10'd241};
ram[48396] = {9'd44,10'd245};
ram[48397] = {9'd47,10'd248};
ram[48398] = {9'd51,10'd251};
ram[48399] = {9'd54,10'd254};
ram[48400] = {9'd57,10'd257};
ram[48401] = {9'd60,10'd260};
ram[48402] = {9'd63,10'd263};
ram[48403] = {9'd66,10'd267};
ram[48404] = {9'd69,10'd270};
ram[48405] = {9'd73,10'd273};
ram[48406] = {9'd76,10'd276};
ram[48407] = {9'd79,10'd279};
ram[48408] = {9'd82,10'd282};
ram[48409] = {9'd85,10'd285};
ram[48410] = {9'd88,10'd289};
ram[48411] = {9'd91,10'd292};
ram[48412] = {9'd95,10'd295};
ram[48413] = {9'd98,10'd298};
ram[48414] = {-9'd99,10'd301};
ram[48415] = {-9'd96,10'd304};
ram[48416] = {-9'd93,10'd307};
ram[48417] = {-9'd90,10'd311};
ram[48418] = {-9'd87,10'd314};
ram[48419] = {-9'd84,10'd317};
ram[48420] = {-9'd81,10'd320};
ram[48421] = {-9'd77,10'd323};
ram[48422] = {-9'd74,10'd326};
ram[48423] = {-9'd71,10'd329};
ram[48424] = {-9'd68,10'd333};
ram[48425] = {-9'd65,10'd336};
ram[48426] = {-9'd62,10'd339};
ram[48427] = {-9'd59,10'd342};
ram[48428] = {-9'd55,10'd345};
ram[48429] = {-9'd52,10'd348};
ram[48430] = {-9'd49,10'd351};
ram[48431] = {-9'd46,10'd354};
ram[48432] = {-9'd43,10'd358};
ram[48433] = {-9'd40,10'd361};
ram[48434] = {-9'd37,10'd364};
ram[48435] = {-9'd33,10'd367};
ram[48436] = {-9'd30,10'd370};
ram[48437] = {-9'd27,10'd373};
ram[48438] = {-9'd24,10'd376};
ram[48439] = {-9'd21,10'd380};
ram[48440] = {-9'd18,10'd383};
ram[48441] = {-9'd15,10'd386};
ram[48442] = {-9'd11,10'd389};
ram[48443] = {-9'd8,10'd392};
ram[48444] = {-9'd5,10'd395};
ram[48445] = {-9'd2,10'd398};
ram[48446] = {9'd1,-10'd399};
ram[48447] = {9'd4,-10'd396};
ram[48448] = {9'd7,-10'd393};
ram[48449] = {9'd10,-10'd390};
ram[48450] = {9'd14,-10'd387};
ram[48451] = {9'd17,-10'd384};
ram[48452] = {9'd20,-10'd381};
ram[48453] = {9'd23,-10'd377};
ram[48454] = {9'd26,-10'd374};
ram[48455] = {9'd29,-10'd371};
ram[48456] = {9'd32,-10'd368};
ram[48457] = {9'd36,-10'd365};
ram[48458] = {9'd39,-10'd362};
ram[48459] = {9'd42,-10'd359};
ram[48460] = {9'd45,-10'd355};
ram[48461] = {9'd48,-10'd352};
ram[48462] = {9'd51,-10'd349};
ram[48463] = {9'd54,-10'd346};
ram[48464] = {9'd58,-10'd343};
ram[48465] = {9'd61,-10'd340};
ram[48466] = {9'd64,-10'd337};
ram[48467] = {9'd67,-10'd334};
ram[48468] = {9'd70,-10'd330};
ram[48469] = {9'd73,-10'd327};
ram[48470] = {9'd76,-10'd324};
ram[48471] = {9'd80,-10'd321};
ram[48472] = {9'd83,-10'd318};
ram[48473] = {9'd86,-10'd315};
ram[48474] = {9'd89,-10'd312};
ram[48475] = {9'd92,-10'd308};
ram[48476] = {9'd95,-10'd305};
ram[48477] = {9'd98,-10'd302};
ram[48478] = {-9'd99,-10'd299};
ram[48479] = {-9'd96,-10'd296};
ram[48480] = {-9'd92,-10'd293};
ram[48481] = {-9'd89,-10'd290};
ram[48482] = {-9'd86,-10'd286};
ram[48483] = {-9'd83,-10'd283};
ram[48484] = {-9'd80,-10'd280};
ram[48485] = {-9'd77,-10'd277};
ram[48486] = {-9'd74,-10'd274};
ram[48487] = {-9'd70,-10'd271};
ram[48488] = {-9'd67,-10'd268};
ram[48489] = {-9'd64,-10'd264};
ram[48490] = {-9'd61,-10'd261};
ram[48491] = {-9'd58,-10'd258};
ram[48492] = {-9'd55,-10'd255};
ram[48493] = {-9'd52,-10'd252};
ram[48494] = {-9'd48,-10'd249};
ram[48495] = {-9'd45,-10'd246};
ram[48496] = {-9'd42,-10'd242};
ram[48497] = {-9'd39,-10'd239};
ram[48498] = {-9'd36,-10'd236};
ram[48499] = {-9'd33,-10'd233};
ram[48500] = {-9'd30,-10'd230};
ram[48501] = {-9'd26,-10'd227};
ram[48502] = {-9'd23,-10'd224};
ram[48503] = {-9'd20,-10'd220};
ram[48504] = {-9'd17,-10'd217};
ram[48505] = {-9'd14,-10'd214};
ram[48506] = {-9'd11,-10'd211};
ram[48507] = {-9'd8,-10'd208};
ram[48508] = {-9'd4,-10'd205};
ram[48509] = {-9'd1,-10'd202};
ram[48510] = {9'd2,-10'd198};
ram[48511] = {9'd5,-10'd195};
ram[48512] = {9'd5,-10'd195};
ram[48513] = {9'd8,-10'd192};
ram[48514] = {9'd11,-10'd189};
ram[48515] = {9'd14,-10'd186};
ram[48516] = {9'd18,-10'd183};
ram[48517] = {9'd21,-10'd180};
ram[48518] = {9'd24,-10'd176};
ram[48519] = {9'd27,-10'd173};
ram[48520] = {9'd30,-10'd170};
ram[48521] = {9'd33,-10'd167};
ram[48522] = {9'd36,-10'd164};
ram[48523] = {9'd40,-10'd161};
ram[48524] = {9'd43,-10'd158};
ram[48525] = {9'd46,-10'd154};
ram[48526] = {9'd49,-10'd151};
ram[48527] = {9'd52,-10'd148};
ram[48528] = {9'd55,-10'd145};
ram[48529] = {9'd58,-10'd142};
ram[48530] = {9'd62,-10'd139};
ram[48531] = {9'd65,-10'd136};
ram[48532] = {9'd68,-10'd132};
ram[48533] = {9'd71,-10'd129};
ram[48534] = {9'd74,-10'd126};
ram[48535] = {9'd77,-10'd123};
ram[48536] = {9'd80,-10'd120};
ram[48537] = {9'd84,-10'd117};
ram[48538] = {9'd87,-10'd114};
ram[48539] = {9'd90,-10'd110};
ram[48540] = {9'd93,-10'd107};
ram[48541] = {9'd96,-10'd104};
ram[48542] = {9'd99,-10'd101};
ram[48543] = {-9'd98,-10'd98};
ram[48544] = {-9'd95,-10'd95};
ram[48545] = {-9'd92,-10'd92};
ram[48546] = {-9'd88,-10'd88};
ram[48547] = {-9'd85,-10'd85};
ram[48548] = {-9'd82,-10'd82};
ram[48549] = {-9'd79,-10'd79};
ram[48550] = {-9'd76,-10'd76};
ram[48551] = {-9'd73,-10'd73};
ram[48552] = {-9'd70,-10'd70};
ram[48553] = {-9'd66,-10'd66};
ram[48554] = {-9'd63,-10'd63};
ram[48555] = {-9'd60,-10'd60};
ram[48556] = {-9'd57,-10'd57};
ram[48557] = {-9'd54,-10'd54};
ram[48558] = {-9'd51,-10'd51};
ram[48559] = {-9'd48,-10'd48};
ram[48560] = {-9'd44,-10'd44};
ram[48561] = {-9'd41,-10'd41};
ram[48562] = {-9'd38,-10'd38};
ram[48563] = {-9'd35,-10'd35};
ram[48564] = {-9'd32,-10'd32};
ram[48565] = {-9'd29,-10'd29};
ram[48566] = {-9'd26,-10'd26};
ram[48567] = {-9'd22,-10'd22};
ram[48568] = {-9'd19,-10'd19};
ram[48569] = {-9'd16,-10'd16};
ram[48570] = {-9'd13,-10'd13};
ram[48571] = {-9'd10,-10'd10};
ram[48572] = {-9'd7,-10'd7};
ram[48573] = {-9'd4,-10'd4};
ram[48574] = {9'd0,10'd0};
ram[48575] = {9'd3,10'd3};
ram[48576] = {9'd6,10'd6};
ram[48577] = {9'd9,10'd9};
ram[48578] = {9'd12,10'd12};
ram[48579] = {9'd15,10'd15};
ram[48580] = {9'd18,10'd18};
ram[48581] = {9'd21,10'd21};
ram[48582] = {9'd25,10'd25};
ram[48583] = {9'd28,10'd28};
ram[48584] = {9'd31,10'd31};
ram[48585] = {9'd34,10'd34};
ram[48586] = {9'd37,10'd37};
ram[48587] = {9'd40,10'd40};
ram[48588] = {9'd43,10'd43};
ram[48589] = {9'd47,10'd47};
ram[48590] = {9'd50,10'd50};
ram[48591] = {9'd53,10'd53};
ram[48592] = {9'd56,10'd56};
ram[48593] = {9'd59,10'd59};
ram[48594] = {9'd62,10'd62};
ram[48595] = {9'd65,10'd65};
ram[48596] = {9'd69,10'd69};
ram[48597] = {9'd72,10'd72};
ram[48598] = {9'd75,10'd75};
ram[48599] = {9'd78,10'd78};
ram[48600] = {9'd81,10'd81};
ram[48601] = {9'd84,10'd84};
ram[48602] = {9'd87,10'd87};
ram[48603] = {9'd91,10'd91};
ram[48604] = {9'd94,10'd94};
ram[48605] = {9'd97,10'd97};
ram[48606] = {-9'd100,10'd100};
ram[48607] = {-9'd97,10'd103};
ram[48608] = {-9'd94,10'd106};
ram[48609] = {-9'd91,10'd109};
ram[48610] = {-9'd88,10'd113};
ram[48611] = {-9'd85,10'd116};
ram[48612] = {-9'd81,10'd119};
ram[48613] = {-9'd78,10'd122};
ram[48614] = {-9'd75,10'd125};
ram[48615] = {-9'd72,10'd128};
ram[48616] = {-9'd69,10'd131};
ram[48617] = {-9'd66,10'd135};
ram[48618] = {-9'd63,10'd138};
ram[48619] = {-9'd59,10'd141};
ram[48620] = {-9'd56,10'd144};
ram[48621] = {-9'd53,10'd147};
ram[48622] = {-9'd50,10'd150};
ram[48623] = {-9'd47,10'd153};
ram[48624] = {-9'd44,10'd157};
ram[48625] = {-9'd41,10'd160};
ram[48626] = {-9'd37,10'd163};
ram[48627] = {-9'd34,10'd166};
ram[48628] = {-9'd31,10'd169};
ram[48629] = {-9'd28,10'd172};
ram[48630] = {-9'd25,10'd175};
ram[48631] = {-9'd22,10'd179};
ram[48632] = {-9'd19,10'd182};
ram[48633] = {-9'd15,10'd185};
ram[48634] = {-9'd12,10'd188};
ram[48635] = {-9'd9,10'd191};
ram[48636] = {-9'd6,10'd194};
ram[48637] = {-9'd3,10'd197};
ram[48638] = {9'd0,10'd201};
ram[48639] = {9'd3,10'd204};
ram[48640] = {9'd3,10'd204};
ram[48641] = {9'd7,10'd207};
ram[48642] = {9'd10,10'd210};
ram[48643] = {9'd13,10'd213};
ram[48644] = {9'd16,10'd216};
ram[48645] = {9'd19,10'd219};
ram[48646] = {9'd22,10'd223};
ram[48647] = {9'd25,10'd226};
ram[48648] = {9'd29,10'd229};
ram[48649] = {9'd32,10'd232};
ram[48650] = {9'd35,10'd235};
ram[48651] = {9'd38,10'd238};
ram[48652] = {9'd41,10'd241};
ram[48653] = {9'd44,10'd245};
ram[48654] = {9'd47,10'd248};
ram[48655] = {9'd51,10'd251};
ram[48656] = {9'd54,10'd254};
ram[48657] = {9'd57,10'd257};
ram[48658] = {9'd60,10'd260};
ram[48659] = {9'd63,10'd263};
ram[48660] = {9'd66,10'd267};
ram[48661] = {9'd69,10'd270};
ram[48662] = {9'd73,10'd273};
ram[48663] = {9'd76,10'd276};
ram[48664] = {9'd79,10'd279};
ram[48665] = {9'd82,10'd282};
ram[48666] = {9'd85,10'd285};
ram[48667] = {9'd88,10'd289};
ram[48668] = {9'd91,10'd292};
ram[48669] = {9'd95,10'd295};
ram[48670] = {9'd98,10'd298};
ram[48671] = {-9'd99,10'd301};
ram[48672] = {-9'd96,10'd304};
ram[48673] = {-9'd93,10'd307};
ram[48674] = {-9'd90,10'd311};
ram[48675] = {-9'd87,10'd314};
ram[48676] = {-9'd84,10'd317};
ram[48677] = {-9'd81,10'd320};
ram[48678] = {-9'd77,10'd323};
ram[48679] = {-9'd74,10'd326};
ram[48680] = {-9'd71,10'd329};
ram[48681] = {-9'd68,10'd333};
ram[48682] = {-9'd65,10'd336};
ram[48683] = {-9'd62,10'd339};
ram[48684] = {-9'd59,10'd342};
ram[48685] = {-9'd55,10'd345};
ram[48686] = {-9'd52,10'd348};
ram[48687] = {-9'd49,10'd351};
ram[48688] = {-9'd46,10'd354};
ram[48689] = {-9'd43,10'd358};
ram[48690] = {-9'd40,10'd361};
ram[48691] = {-9'd37,10'd364};
ram[48692] = {-9'd33,10'd367};
ram[48693] = {-9'd30,10'd370};
ram[48694] = {-9'd27,10'd373};
ram[48695] = {-9'd24,10'd376};
ram[48696] = {-9'd21,10'd380};
ram[48697] = {-9'd18,10'd383};
ram[48698] = {-9'd15,10'd386};
ram[48699] = {-9'd11,10'd389};
ram[48700] = {-9'd8,10'd392};
ram[48701] = {-9'd5,10'd395};
ram[48702] = {-9'd2,10'd398};
ram[48703] = {9'd1,-10'd399};
ram[48704] = {9'd4,-10'd396};
ram[48705] = {9'd7,-10'd393};
ram[48706] = {9'd10,-10'd390};
ram[48707] = {9'd14,-10'd387};
ram[48708] = {9'd17,-10'd384};
ram[48709] = {9'd20,-10'd381};
ram[48710] = {9'd23,-10'd377};
ram[48711] = {9'd26,-10'd374};
ram[48712] = {9'd29,-10'd371};
ram[48713] = {9'd32,-10'd368};
ram[48714] = {9'd36,-10'd365};
ram[48715] = {9'd39,-10'd362};
ram[48716] = {9'd42,-10'd359};
ram[48717] = {9'd45,-10'd355};
ram[48718] = {9'd48,-10'd352};
ram[48719] = {9'd51,-10'd349};
ram[48720] = {9'd54,-10'd346};
ram[48721] = {9'd58,-10'd343};
ram[48722] = {9'd61,-10'd340};
ram[48723] = {9'd64,-10'd337};
ram[48724] = {9'd67,-10'd334};
ram[48725] = {9'd70,-10'd330};
ram[48726] = {9'd73,-10'd327};
ram[48727] = {9'd76,-10'd324};
ram[48728] = {9'd80,-10'd321};
ram[48729] = {9'd83,-10'd318};
ram[48730] = {9'd86,-10'd315};
ram[48731] = {9'd89,-10'd312};
ram[48732] = {9'd92,-10'd308};
ram[48733] = {9'd95,-10'd305};
ram[48734] = {9'd98,-10'd302};
ram[48735] = {-9'd99,-10'd299};
ram[48736] = {-9'd96,-10'd296};
ram[48737] = {-9'd92,-10'd293};
ram[48738] = {-9'd89,-10'd290};
ram[48739] = {-9'd86,-10'd286};
ram[48740] = {-9'd83,-10'd283};
ram[48741] = {-9'd80,-10'd280};
ram[48742] = {-9'd77,-10'd277};
ram[48743] = {-9'd74,-10'd274};
ram[48744] = {-9'd70,-10'd271};
ram[48745] = {-9'd67,-10'd268};
ram[48746] = {-9'd64,-10'd264};
ram[48747] = {-9'd61,-10'd261};
ram[48748] = {-9'd58,-10'd258};
ram[48749] = {-9'd55,-10'd255};
ram[48750] = {-9'd52,-10'd252};
ram[48751] = {-9'd48,-10'd249};
ram[48752] = {-9'd45,-10'd246};
ram[48753] = {-9'd42,-10'd242};
ram[48754] = {-9'd39,-10'd239};
ram[48755] = {-9'd36,-10'd236};
ram[48756] = {-9'd33,-10'd233};
ram[48757] = {-9'd30,-10'd230};
ram[48758] = {-9'd26,-10'd227};
ram[48759] = {-9'd23,-10'd224};
ram[48760] = {-9'd20,-10'd220};
ram[48761] = {-9'd17,-10'd217};
ram[48762] = {-9'd14,-10'd214};
ram[48763] = {-9'd11,-10'd211};
ram[48764] = {-9'd8,-10'd208};
ram[48765] = {-9'd4,-10'd205};
ram[48766] = {-9'd1,-10'd202};
ram[48767] = {9'd2,-10'd198};
ram[48768] = {9'd2,-10'd198};
ram[48769] = {9'd5,-10'd195};
ram[48770] = {9'd8,-10'd192};
ram[48771] = {9'd11,-10'd189};
ram[48772] = {9'd14,-10'd186};
ram[48773] = {9'd18,-10'd183};
ram[48774] = {9'd21,-10'd180};
ram[48775] = {9'd24,-10'd176};
ram[48776] = {9'd27,-10'd173};
ram[48777] = {9'd30,-10'd170};
ram[48778] = {9'd33,-10'd167};
ram[48779] = {9'd36,-10'd164};
ram[48780] = {9'd40,-10'd161};
ram[48781] = {9'd43,-10'd158};
ram[48782] = {9'd46,-10'd154};
ram[48783] = {9'd49,-10'd151};
ram[48784] = {9'd52,-10'd148};
ram[48785] = {9'd55,-10'd145};
ram[48786] = {9'd58,-10'd142};
ram[48787] = {9'd62,-10'd139};
ram[48788] = {9'd65,-10'd136};
ram[48789] = {9'd68,-10'd132};
ram[48790] = {9'd71,-10'd129};
ram[48791] = {9'd74,-10'd126};
ram[48792] = {9'd77,-10'd123};
ram[48793] = {9'd80,-10'd120};
ram[48794] = {9'd84,-10'd117};
ram[48795] = {9'd87,-10'd114};
ram[48796] = {9'd90,-10'd110};
ram[48797] = {9'd93,-10'd107};
ram[48798] = {9'd96,-10'd104};
ram[48799] = {9'd99,-10'd101};
ram[48800] = {-9'd98,-10'd98};
ram[48801] = {-9'd95,-10'd95};
ram[48802] = {-9'd92,-10'd92};
ram[48803] = {-9'd88,-10'd88};
ram[48804] = {-9'd85,-10'd85};
ram[48805] = {-9'd82,-10'd82};
ram[48806] = {-9'd79,-10'd79};
ram[48807] = {-9'd76,-10'd76};
ram[48808] = {-9'd73,-10'd73};
ram[48809] = {-9'd70,-10'd70};
ram[48810] = {-9'd66,-10'd66};
ram[48811] = {-9'd63,-10'd63};
ram[48812] = {-9'd60,-10'd60};
ram[48813] = {-9'd57,-10'd57};
ram[48814] = {-9'd54,-10'd54};
ram[48815] = {-9'd51,-10'd51};
ram[48816] = {-9'd48,-10'd48};
ram[48817] = {-9'd44,-10'd44};
ram[48818] = {-9'd41,-10'd41};
ram[48819] = {-9'd38,-10'd38};
ram[48820] = {-9'd35,-10'd35};
ram[48821] = {-9'd32,-10'd32};
ram[48822] = {-9'd29,-10'd29};
ram[48823] = {-9'd26,-10'd26};
ram[48824] = {-9'd22,-10'd22};
ram[48825] = {-9'd19,-10'd19};
ram[48826] = {-9'd16,-10'd16};
ram[48827] = {-9'd13,-10'd13};
ram[48828] = {-9'd10,-10'd10};
ram[48829] = {-9'd7,-10'd7};
ram[48830] = {-9'd4,-10'd4};
ram[48831] = {9'd0,10'd0};
ram[48832] = {9'd3,10'd3};
ram[48833] = {9'd6,10'd6};
ram[48834] = {9'd9,10'd9};
ram[48835] = {9'd12,10'd12};
ram[48836] = {9'd15,10'd15};
ram[48837] = {9'd18,10'd18};
ram[48838] = {9'd21,10'd21};
ram[48839] = {9'd25,10'd25};
ram[48840] = {9'd28,10'd28};
ram[48841] = {9'd31,10'd31};
ram[48842] = {9'd34,10'd34};
ram[48843] = {9'd37,10'd37};
ram[48844] = {9'd40,10'd40};
ram[48845] = {9'd43,10'd43};
ram[48846] = {9'd47,10'd47};
ram[48847] = {9'd50,10'd50};
ram[48848] = {9'd53,10'd53};
ram[48849] = {9'd56,10'd56};
ram[48850] = {9'd59,10'd59};
ram[48851] = {9'd62,10'd62};
ram[48852] = {9'd65,10'd65};
ram[48853] = {9'd69,10'd69};
ram[48854] = {9'd72,10'd72};
ram[48855] = {9'd75,10'd75};
ram[48856] = {9'd78,10'd78};
ram[48857] = {9'd81,10'd81};
ram[48858] = {9'd84,10'd84};
ram[48859] = {9'd87,10'd87};
ram[48860] = {9'd91,10'd91};
ram[48861] = {9'd94,10'd94};
ram[48862] = {9'd97,10'd97};
ram[48863] = {-9'd100,10'd100};
ram[48864] = {-9'd97,10'd103};
ram[48865] = {-9'd94,10'd106};
ram[48866] = {-9'd91,10'd109};
ram[48867] = {-9'd88,10'd113};
ram[48868] = {-9'd85,10'd116};
ram[48869] = {-9'd81,10'd119};
ram[48870] = {-9'd78,10'd122};
ram[48871] = {-9'd75,10'd125};
ram[48872] = {-9'd72,10'd128};
ram[48873] = {-9'd69,10'd131};
ram[48874] = {-9'd66,10'd135};
ram[48875] = {-9'd63,10'd138};
ram[48876] = {-9'd59,10'd141};
ram[48877] = {-9'd56,10'd144};
ram[48878] = {-9'd53,10'd147};
ram[48879] = {-9'd50,10'd150};
ram[48880] = {-9'd47,10'd153};
ram[48881] = {-9'd44,10'd157};
ram[48882] = {-9'd41,10'd160};
ram[48883] = {-9'd37,10'd163};
ram[48884] = {-9'd34,10'd166};
ram[48885] = {-9'd31,10'd169};
ram[48886] = {-9'd28,10'd172};
ram[48887] = {-9'd25,10'd175};
ram[48888] = {-9'd22,10'd179};
ram[48889] = {-9'd19,10'd182};
ram[48890] = {-9'd15,10'd185};
ram[48891] = {-9'd12,10'd188};
ram[48892] = {-9'd9,10'd191};
ram[48893] = {-9'd6,10'd194};
ram[48894] = {-9'd3,10'd197};
ram[48895] = {9'd0,10'd201};
ram[48896] = {9'd0,10'd201};
ram[48897] = {9'd3,10'd204};
ram[48898] = {9'd7,10'd207};
ram[48899] = {9'd10,10'd210};
ram[48900] = {9'd13,10'd213};
ram[48901] = {9'd16,10'd216};
ram[48902] = {9'd19,10'd219};
ram[48903] = {9'd22,10'd223};
ram[48904] = {9'd25,10'd226};
ram[48905] = {9'd29,10'd229};
ram[48906] = {9'd32,10'd232};
ram[48907] = {9'd35,10'd235};
ram[48908] = {9'd38,10'd238};
ram[48909] = {9'd41,10'd241};
ram[48910] = {9'd44,10'd245};
ram[48911] = {9'd47,10'd248};
ram[48912] = {9'd51,10'd251};
ram[48913] = {9'd54,10'd254};
ram[48914] = {9'd57,10'd257};
ram[48915] = {9'd60,10'd260};
ram[48916] = {9'd63,10'd263};
ram[48917] = {9'd66,10'd267};
ram[48918] = {9'd69,10'd270};
ram[48919] = {9'd73,10'd273};
ram[48920] = {9'd76,10'd276};
ram[48921] = {9'd79,10'd279};
ram[48922] = {9'd82,10'd282};
ram[48923] = {9'd85,10'd285};
ram[48924] = {9'd88,10'd289};
ram[48925] = {9'd91,10'd292};
ram[48926] = {9'd95,10'd295};
ram[48927] = {9'd98,10'd298};
ram[48928] = {-9'd99,10'd301};
ram[48929] = {-9'd96,10'd304};
ram[48930] = {-9'd93,10'd307};
ram[48931] = {-9'd90,10'd311};
ram[48932] = {-9'd87,10'd314};
ram[48933] = {-9'd84,10'd317};
ram[48934] = {-9'd81,10'd320};
ram[48935] = {-9'd77,10'd323};
ram[48936] = {-9'd74,10'd326};
ram[48937] = {-9'd71,10'd329};
ram[48938] = {-9'd68,10'd333};
ram[48939] = {-9'd65,10'd336};
ram[48940] = {-9'd62,10'd339};
ram[48941] = {-9'd59,10'd342};
ram[48942] = {-9'd55,10'd345};
ram[48943] = {-9'd52,10'd348};
ram[48944] = {-9'd49,10'd351};
ram[48945] = {-9'd46,10'd354};
ram[48946] = {-9'd43,10'd358};
ram[48947] = {-9'd40,10'd361};
ram[48948] = {-9'd37,10'd364};
ram[48949] = {-9'd33,10'd367};
ram[48950] = {-9'd30,10'd370};
ram[48951] = {-9'd27,10'd373};
ram[48952] = {-9'd24,10'd376};
ram[48953] = {-9'd21,10'd380};
ram[48954] = {-9'd18,10'd383};
ram[48955] = {-9'd15,10'd386};
ram[48956] = {-9'd11,10'd389};
ram[48957] = {-9'd8,10'd392};
ram[48958] = {-9'd5,10'd395};
ram[48959] = {-9'd2,10'd398};
ram[48960] = {9'd1,-10'd399};
ram[48961] = {9'd4,-10'd396};
ram[48962] = {9'd7,-10'd393};
ram[48963] = {9'd10,-10'd390};
ram[48964] = {9'd14,-10'd387};
ram[48965] = {9'd17,-10'd384};
ram[48966] = {9'd20,-10'd381};
ram[48967] = {9'd23,-10'd377};
ram[48968] = {9'd26,-10'd374};
ram[48969] = {9'd29,-10'd371};
ram[48970] = {9'd32,-10'd368};
ram[48971] = {9'd36,-10'd365};
ram[48972] = {9'd39,-10'd362};
ram[48973] = {9'd42,-10'd359};
ram[48974] = {9'd45,-10'd355};
ram[48975] = {9'd48,-10'd352};
ram[48976] = {9'd51,-10'd349};
ram[48977] = {9'd54,-10'd346};
ram[48978] = {9'd58,-10'd343};
ram[48979] = {9'd61,-10'd340};
ram[48980] = {9'd64,-10'd337};
ram[48981] = {9'd67,-10'd334};
ram[48982] = {9'd70,-10'd330};
ram[48983] = {9'd73,-10'd327};
ram[48984] = {9'd76,-10'd324};
ram[48985] = {9'd80,-10'd321};
ram[48986] = {9'd83,-10'd318};
ram[48987] = {9'd86,-10'd315};
ram[48988] = {9'd89,-10'd312};
ram[48989] = {9'd92,-10'd308};
ram[48990] = {9'd95,-10'd305};
ram[48991] = {9'd98,-10'd302};
ram[48992] = {-9'd99,-10'd299};
ram[48993] = {-9'd96,-10'd296};
ram[48994] = {-9'd92,-10'd293};
ram[48995] = {-9'd89,-10'd290};
ram[48996] = {-9'd86,-10'd286};
ram[48997] = {-9'd83,-10'd283};
ram[48998] = {-9'd80,-10'd280};
ram[48999] = {-9'd77,-10'd277};
ram[49000] = {-9'd74,-10'd274};
ram[49001] = {-9'd70,-10'd271};
ram[49002] = {-9'd67,-10'd268};
ram[49003] = {-9'd64,-10'd264};
ram[49004] = {-9'd61,-10'd261};
ram[49005] = {-9'd58,-10'd258};
ram[49006] = {-9'd55,-10'd255};
ram[49007] = {-9'd52,-10'd252};
ram[49008] = {-9'd48,-10'd249};
ram[49009] = {-9'd45,-10'd246};
ram[49010] = {-9'd42,-10'd242};
ram[49011] = {-9'd39,-10'd239};
ram[49012] = {-9'd36,-10'd236};
ram[49013] = {-9'd33,-10'd233};
ram[49014] = {-9'd30,-10'd230};
ram[49015] = {-9'd26,-10'd227};
ram[49016] = {-9'd23,-10'd224};
ram[49017] = {-9'd20,-10'd220};
ram[49018] = {-9'd17,-10'd217};
ram[49019] = {-9'd14,-10'd214};
ram[49020] = {-9'd11,-10'd211};
ram[49021] = {-9'd8,-10'd208};
ram[49022] = {-9'd4,-10'd205};
ram[49023] = {-9'd1,-10'd202};
ram[49024] = {-9'd1,-10'd202};
ram[49025] = {9'd2,-10'd198};
ram[49026] = {9'd5,-10'd195};
ram[49027] = {9'd8,-10'd192};
ram[49028] = {9'd11,-10'd189};
ram[49029] = {9'd14,-10'd186};
ram[49030] = {9'd18,-10'd183};
ram[49031] = {9'd21,-10'd180};
ram[49032] = {9'd24,-10'd176};
ram[49033] = {9'd27,-10'd173};
ram[49034] = {9'd30,-10'd170};
ram[49035] = {9'd33,-10'd167};
ram[49036] = {9'd36,-10'd164};
ram[49037] = {9'd40,-10'd161};
ram[49038] = {9'd43,-10'd158};
ram[49039] = {9'd46,-10'd154};
ram[49040] = {9'd49,-10'd151};
ram[49041] = {9'd52,-10'd148};
ram[49042] = {9'd55,-10'd145};
ram[49043] = {9'd58,-10'd142};
ram[49044] = {9'd62,-10'd139};
ram[49045] = {9'd65,-10'd136};
ram[49046] = {9'd68,-10'd132};
ram[49047] = {9'd71,-10'd129};
ram[49048] = {9'd74,-10'd126};
ram[49049] = {9'd77,-10'd123};
ram[49050] = {9'd80,-10'd120};
ram[49051] = {9'd84,-10'd117};
ram[49052] = {9'd87,-10'd114};
ram[49053] = {9'd90,-10'd110};
ram[49054] = {9'd93,-10'd107};
ram[49055] = {9'd96,-10'd104};
ram[49056] = {9'd99,-10'd101};
ram[49057] = {-9'd98,-10'd98};
ram[49058] = {-9'd95,-10'd95};
ram[49059] = {-9'd92,-10'd92};
ram[49060] = {-9'd88,-10'd88};
ram[49061] = {-9'd85,-10'd85};
ram[49062] = {-9'd82,-10'd82};
ram[49063] = {-9'd79,-10'd79};
ram[49064] = {-9'd76,-10'd76};
ram[49065] = {-9'd73,-10'd73};
ram[49066] = {-9'd70,-10'd70};
ram[49067] = {-9'd66,-10'd66};
ram[49068] = {-9'd63,-10'd63};
ram[49069] = {-9'd60,-10'd60};
ram[49070] = {-9'd57,-10'd57};
ram[49071] = {-9'd54,-10'd54};
ram[49072] = {-9'd51,-10'd51};
ram[49073] = {-9'd48,-10'd48};
ram[49074] = {-9'd44,-10'd44};
ram[49075] = {-9'd41,-10'd41};
ram[49076] = {-9'd38,-10'd38};
ram[49077] = {-9'd35,-10'd35};
ram[49078] = {-9'd32,-10'd32};
ram[49079] = {-9'd29,-10'd29};
ram[49080] = {-9'd26,-10'd26};
ram[49081] = {-9'd22,-10'd22};
ram[49082] = {-9'd19,-10'd19};
ram[49083] = {-9'd16,-10'd16};
ram[49084] = {-9'd13,-10'd13};
ram[49085] = {-9'd10,-10'd10};
ram[49086] = {-9'd7,-10'd7};
ram[49087] = {-9'd4,-10'd4};
ram[49088] = {9'd0,10'd0};
ram[49089] = {9'd3,10'd3};
ram[49090] = {9'd6,10'd6};
ram[49091] = {9'd9,10'd9};
ram[49092] = {9'd12,10'd12};
ram[49093] = {9'd15,10'd15};
ram[49094] = {9'd18,10'd18};
ram[49095] = {9'd21,10'd21};
ram[49096] = {9'd25,10'd25};
ram[49097] = {9'd28,10'd28};
ram[49098] = {9'd31,10'd31};
ram[49099] = {9'd34,10'd34};
ram[49100] = {9'd37,10'd37};
ram[49101] = {9'd40,10'd40};
ram[49102] = {9'd43,10'd43};
ram[49103] = {9'd47,10'd47};
ram[49104] = {9'd50,10'd50};
ram[49105] = {9'd53,10'd53};
ram[49106] = {9'd56,10'd56};
ram[49107] = {9'd59,10'd59};
ram[49108] = {9'd62,10'd62};
ram[49109] = {9'd65,10'd65};
ram[49110] = {9'd69,10'd69};
ram[49111] = {9'd72,10'd72};
ram[49112] = {9'd75,10'd75};
ram[49113] = {9'd78,10'd78};
ram[49114] = {9'd81,10'd81};
ram[49115] = {9'd84,10'd84};
ram[49116] = {9'd87,10'd87};
ram[49117] = {9'd91,10'd91};
ram[49118] = {9'd94,10'd94};
ram[49119] = {9'd97,10'd97};
ram[49120] = {-9'd100,10'd100};
ram[49121] = {-9'd97,10'd103};
ram[49122] = {-9'd94,10'd106};
ram[49123] = {-9'd91,10'd109};
ram[49124] = {-9'd88,10'd113};
ram[49125] = {-9'd85,10'd116};
ram[49126] = {-9'd81,10'd119};
ram[49127] = {-9'd78,10'd122};
ram[49128] = {-9'd75,10'd125};
ram[49129] = {-9'd72,10'd128};
ram[49130] = {-9'd69,10'd131};
ram[49131] = {-9'd66,10'd135};
ram[49132] = {-9'd63,10'd138};
ram[49133] = {-9'd59,10'd141};
ram[49134] = {-9'd56,10'd144};
ram[49135] = {-9'd53,10'd147};
ram[49136] = {-9'd50,10'd150};
ram[49137] = {-9'd47,10'd153};
ram[49138] = {-9'd44,10'd157};
ram[49139] = {-9'd41,10'd160};
ram[49140] = {-9'd37,10'd163};
ram[49141] = {-9'd34,10'd166};
ram[49142] = {-9'd31,10'd169};
ram[49143] = {-9'd28,10'd172};
ram[49144] = {-9'd25,10'd175};
ram[49145] = {-9'd22,10'd179};
ram[49146] = {-9'd19,10'd182};
ram[49147] = {-9'd15,10'd185};
ram[49148] = {-9'd12,10'd188};
ram[49149] = {-9'd9,10'd191};
ram[49150] = {-9'd6,10'd194};
ram[49151] = {-9'd3,10'd197};
ram[49152] = {-9'd3,10'd197};
ram[49153] = {9'd0,10'd201};
ram[49154] = {9'd3,10'd204};
ram[49155] = {9'd7,10'd207};
ram[49156] = {9'd10,10'd210};
ram[49157] = {9'd13,10'd213};
ram[49158] = {9'd16,10'd216};
ram[49159] = {9'd19,10'd219};
ram[49160] = {9'd22,10'd223};
ram[49161] = {9'd25,10'd226};
ram[49162] = {9'd29,10'd229};
ram[49163] = {9'd32,10'd232};
ram[49164] = {9'd35,10'd235};
ram[49165] = {9'd38,10'd238};
ram[49166] = {9'd41,10'd241};
ram[49167] = {9'd44,10'd245};
ram[49168] = {9'd47,10'd248};
ram[49169] = {9'd51,10'd251};
ram[49170] = {9'd54,10'd254};
ram[49171] = {9'd57,10'd257};
ram[49172] = {9'd60,10'd260};
ram[49173] = {9'd63,10'd263};
ram[49174] = {9'd66,10'd267};
ram[49175] = {9'd69,10'd270};
ram[49176] = {9'd73,10'd273};
ram[49177] = {9'd76,10'd276};
ram[49178] = {9'd79,10'd279};
ram[49179] = {9'd82,10'd282};
ram[49180] = {9'd85,10'd285};
ram[49181] = {9'd88,10'd289};
ram[49182] = {9'd91,10'd292};
ram[49183] = {9'd95,10'd295};
ram[49184] = {9'd98,10'd298};
ram[49185] = {-9'd99,10'd301};
ram[49186] = {-9'd96,10'd304};
ram[49187] = {-9'd93,10'd307};
ram[49188] = {-9'd90,10'd311};
ram[49189] = {-9'd87,10'd314};
ram[49190] = {-9'd84,10'd317};
ram[49191] = {-9'd81,10'd320};
ram[49192] = {-9'd77,10'd323};
ram[49193] = {-9'd74,10'd326};
ram[49194] = {-9'd71,10'd329};
ram[49195] = {-9'd68,10'd333};
ram[49196] = {-9'd65,10'd336};
ram[49197] = {-9'd62,10'd339};
ram[49198] = {-9'd59,10'd342};
ram[49199] = {-9'd55,10'd345};
ram[49200] = {-9'd52,10'd348};
ram[49201] = {-9'd49,10'd351};
ram[49202] = {-9'd46,10'd354};
ram[49203] = {-9'd43,10'd358};
ram[49204] = {-9'd40,10'd361};
ram[49205] = {-9'd37,10'd364};
ram[49206] = {-9'd33,10'd367};
ram[49207] = {-9'd30,10'd370};
ram[49208] = {-9'd27,10'd373};
ram[49209] = {-9'd24,10'd376};
ram[49210] = {-9'd21,10'd380};
ram[49211] = {-9'd18,10'd383};
ram[49212] = {-9'd15,10'd386};
ram[49213] = {-9'd11,10'd389};
ram[49214] = {-9'd8,10'd392};
ram[49215] = {-9'd5,10'd395};
ram[49216] = {-9'd2,10'd398};
ram[49217] = {9'd1,-10'd399};
ram[49218] = {9'd4,-10'd396};
ram[49219] = {9'd7,-10'd393};
ram[49220] = {9'd10,-10'd390};
ram[49221] = {9'd14,-10'd387};
ram[49222] = {9'd17,-10'd384};
ram[49223] = {9'd20,-10'd381};
ram[49224] = {9'd23,-10'd377};
ram[49225] = {9'd26,-10'd374};
ram[49226] = {9'd29,-10'd371};
ram[49227] = {9'd32,-10'd368};
ram[49228] = {9'd36,-10'd365};
ram[49229] = {9'd39,-10'd362};
ram[49230] = {9'd42,-10'd359};
ram[49231] = {9'd45,-10'd355};
ram[49232] = {9'd48,-10'd352};
ram[49233] = {9'd51,-10'd349};
ram[49234] = {9'd54,-10'd346};
ram[49235] = {9'd58,-10'd343};
ram[49236] = {9'd61,-10'd340};
ram[49237] = {9'd64,-10'd337};
ram[49238] = {9'd67,-10'd334};
ram[49239] = {9'd70,-10'd330};
ram[49240] = {9'd73,-10'd327};
ram[49241] = {9'd76,-10'd324};
ram[49242] = {9'd80,-10'd321};
ram[49243] = {9'd83,-10'd318};
ram[49244] = {9'd86,-10'd315};
ram[49245] = {9'd89,-10'd312};
ram[49246] = {9'd92,-10'd308};
ram[49247] = {9'd95,-10'd305};
ram[49248] = {9'd98,-10'd302};
ram[49249] = {-9'd99,-10'd299};
ram[49250] = {-9'd96,-10'd296};
ram[49251] = {-9'd92,-10'd293};
ram[49252] = {-9'd89,-10'd290};
ram[49253] = {-9'd86,-10'd286};
ram[49254] = {-9'd83,-10'd283};
ram[49255] = {-9'd80,-10'd280};
ram[49256] = {-9'd77,-10'd277};
ram[49257] = {-9'd74,-10'd274};
ram[49258] = {-9'd70,-10'd271};
ram[49259] = {-9'd67,-10'd268};
ram[49260] = {-9'd64,-10'd264};
ram[49261] = {-9'd61,-10'd261};
ram[49262] = {-9'd58,-10'd258};
ram[49263] = {-9'd55,-10'd255};
ram[49264] = {-9'd52,-10'd252};
ram[49265] = {-9'd48,-10'd249};
ram[49266] = {-9'd45,-10'd246};
ram[49267] = {-9'd42,-10'd242};
ram[49268] = {-9'd39,-10'd239};
ram[49269] = {-9'd36,-10'd236};
ram[49270] = {-9'd33,-10'd233};
ram[49271] = {-9'd30,-10'd230};
ram[49272] = {-9'd26,-10'd227};
ram[49273] = {-9'd23,-10'd224};
ram[49274] = {-9'd20,-10'd220};
ram[49275] = {-9'd17,-10'd217};
ram[49276] = {-9'd14,-10'd214};
ram[49277] = {-9'd11,-10'd211};
ram[49278] = {-9'd8,-10'd208};
ram[49279] = {-9'd4,-10'd205};
ram[49280] = {-9'd4,-10'd205};
ram[49281] = {-9'd1,-10'd202};
ram[49282] = {9'd2,-10'd198};
ram[49283] = {9'd5,-10'd195};
ram[49284] = {9'd8,-10'd192};
ram[49285] = {9'd11,-10'd189};
ram[49286] = {9'd14,-10'd186};
ram[49287] = {9'd18,-10'd183};
ram[49288] = {9'd21,-10'd180};
ram[49289] = {9'd24,-10'd176};
ram[49290] = {9'd27,-10'd173};
ram[49291] = {9'd30,-10'd170};
ram[49292] = {9'd33,-10'd167};
ram[49293] = {9'd36,-10'd164};
ram[49294] = {9'd40,-10'd161};
ram[49295] = {9'd43,-10'd158};
ram[49296] = {9'd46,-10'd154};
ram[49297] = {9'd49,-10'd151};
ram[49298] = {9'd52,-10'd148};
ram[49299] = {9'd55,-10'd145};
ram[49300] = {9'd58,-10'd142};
ram[49301] = {9'd62,-10'd139};
ram[49302] = {9'd65,-10'd136};
ram[49303] = {9'd68,-10'd132};
ram[49304] = {9'd71,-10'd129};
ram[49305] = {9'd74,-10'd126};
ram[49306] = {9'd77,-10'd123};
ram[49307] = {9'd80,-10'd120};
ram[49308] = {9'd84,-10'd117};
ram[49309] = {9'd87,-10'd114};
ram[49310] = {9'd90,-10'd110};
ram[49311] = {9'd93,-10'd107};
ram[49312] = {9'd96,-10'd104};
ram[49313] = {9'd99,-10'd101};
ram[49314] = {-9'd98,-10'd98};
ram[49315] = {-9'd95,-10'd95};
ram[49316] = {-9'd92,-10'd92};
ram[49317] = {-9'd88,-10'd88};
ram[49318] = {-9'd85,-10'd85};
ram[49319] = {-9'd82,-10'd82};
ram[49320] = {-9'd79,-10'd79};
ram[49321] = {-9'd76,-10'd76};
ram[49322] = {-9'd73,-10'd73};
ram[49323] = {-9'd70,-10'd70};
ram[49324] = {-9'd66,-10'd66};
ram[49325] = {-9'd63,-10'd63};
ram[49326] = {-9'd60,-10'd60};
ram[49327] = {-9'd57,-10'd57};
ram[49328] = {-9'd54,-10'd54};
ram[49329] = {-9'd51,-10'd51};
ram[49330] = {-9'd48,-10'd48};
ram[49331] = {-9'd44,-10'd44};
ram[49332] = {-9'd41,-10'd41};
ram[49333] = {-9'd38,-10'd38};
ram[49334] = {-9'd35,-10'd35};
ram[49335] = {-9'd32,-10'd32};
ram[49336] = {-9'd29,-10'd29};
ram[49337] = {-9'd26,-10'd26};
ram[49338] = {-9'd22,-10'd22};
ram[49339] = {-9'd19,-10'd19};
ram[49340] = {-9'd16,-10'd16};
ram[49341] = {-9'd13,-10'd13};
ram[49342] = {-9'd10,-10'd10};
ram[49343] = {-9'd7,-10'd7};
ram[49344] = {-9'd4,-10'd4};
ram[49345] = {9'd0,10'd0};
ram[49346] = {9'd3,10'd3};
ram[49347] = {9'd6,10'd6};
ram[49348] = {9'd9,10'd9};
ram[49349] = {9'd12,10'd12};
ram[49350] = {9'd15,10'd15};
ram[49351] = {9'd18,10'd18};
ram[49352] = {9'd21,10'd21};
ram[49353] = {9'd25,10'd25};
ram[49354] = {9'd28,10'd28};
ram[49355] = {9'd31,10'd31};
ram[49356] = {9'd34,10'd34};
ram[49357] = {9'd37,10'd37};
ram[49358] = {9'd40,10'd40};
ram[49359] = {9'd43,10'd43};
ram[49360] = {9'd47,10'd47};
ram[49361] = {9'd50,10'd50};
ram[49362] = {9'd53,10'd53};
ram[49363] = {9'd56,10'd56};
ram[49364] = {9'd59,10'd59};
ram[49365] = {9'd62,10'd62};
ram[49366] = {9'd65,10'd65};
ram[49367] = {9'd69,10'd69};
ram[49368] = {9'd72,10'd72};
ram[49369] = {9'd75,10'd75};
ram[49370] = {9'd78,10'd78};
ram[49371] = {9'd81,10'd81};
ram[49372] = {9'd84,10'd84};
ram[49373] = {9'd87,10'd87};
ram[49374] = {9'd91,10'd91};
ram[49375] = {9'd94,10'd94};
ram[49376] = {9'd97,10'd97};
ram[49377] = {-9'd100,10'd100};
ram[49378] = {-9'd97,10'd103};
ram[49379] = {-9'd94,10'd106};
ram[49380] = {-9'd91,10'd109};
ram[49381] = {-9'd88,10'd113};
ram[49382] = {-9'd85,10'd116};
ram[49383] = {-9'd81,10'd119};
ram[49384] = {-9'd78,10'd122};
ram[49385] = {-9'd75,10'd125};
ram[49386] = {-9'd72,10'd128};
ram[49387] = {-9'd69,10'd131};
ram[49388] = {-9'd66,10'd135};
ram[49389] = {-9'd63,10'd138};
ram[49390] = {-9'd59,10'd141};
ram[49391] = {-9'd56,10'd144};
ram[49392] = {-9'd53,10'd147};
ram[49393] = {-9'd50,10'd150};
ram[49394] = {-9'd47,10'd153};
ram[49395] = {-9'd44,10'd157};
ram[49396] = {-9'd41,10'd160};
ram[49397] = {-9'd37,10'd163};
ram[49398] = {-9'd34,10'd166};
ram[49399] = {-9'd31,10'd169};
ram[49400] = {-9'd28,10'd172};
ram[49401] = {-9'd25,10'd175};
ram[49402] = {-9'd22,10'd179};
ram[49403] = {-9'd19,10'd182};
ram[49404] = {-9'd15,10'd185};
ram[49405] = {-9'd12,10'd188};
ram[49406] = {-9'd9,10'd191};
ram[49407] = {-9'd6,10'd194};
ram[49408] = {-9'd6,10'd194};
ram[49409] = {-9'd3,10'd197};
ram[49410] = {9'd0,10'd201};
ram[49411] = {9'd3,10'd204};
ram[49412] = {9'd7,10'd207};
ram[49413] = {9'd10,10'd210};
ram[49414] = {9'd13,10'd213};
ram[49415] = {9'd16,10'd216};
ram[49416] = {9'd19,10'd219};
ram[49417] = {9'd22,10'd223};
ram[49418] = {9'd25,10'd226};
ram[49419] = {9'd29,10'd229};
ram[49420] = {9'd32,10'd232};
ram[49421] = {9'd35,10'd235};
ram[49422] = {9'd38,10'd238};
ram[49423] = {9'd41,10'd241};
ram[49424] = {9'd44,10'd245};
ram[49425] = {9'd47,10'd248};
ram[49426] = {9'd51,10'd251};
ram[49427] = {9'd54,10'd254};
ram[49428] = {9'd57,10'd257};
ram[49429] = {9'd60,10'd260};
ram[49430] = {9'd63,10'd263};
ram[49431] = {9'd66,10'd267};
ram[49432] = {9'd69,10'd270};
ram[49433] = {9'd73,10'd273};
ram[49434] = {9'd76,10'd276};
ram[49435] = {9'd79,10'd279};
ram[49436] = {9'd82,10'd282};
ram[49437] = {9'd85,10'd285};
ram[49438] = {9'd88,10'd289};
ram[49439] = {9'd91,10'd292};
ram[49440] = {9'd95,10'd295};
ram[49441] = {9'd98,10'd298};
ram[49442] = {-9'd99,10'd301};
ram[49443] = {-9'd96,10'd304};
ram[49444] = {-9'd93,10'd307};
ram[49445] = {-9'd90,10'd311};
ram[49446] = {-9'd87,10'd314};
ram[49447] = {-9'd84,10'd317};
ram[49448] = {-9'd81,10'd320};
ram[49449] = {-9'd77,10'd323};
ram[49450] = {-9'd74,10'd326};
ram[49451] = {-9'd71,10'd329};
ram[49452] = {-9'd68,10'd333};
ram[49453] = {-9'd65,10'd336};
ram[49454] = {-9'd62,10'd339};
ram[49455] = {-9'd59,10'd342};
ram[49456] = {-9'd55,10'd345};
ram[49457] = {-9'd52,10'd348};
ram[49458] = {-9'd49,10'd351};
ram[49459] = {-9'd46,10'd354};
ram[49460] = {-9'd43,10'd358};
ram[49461] = {-9'd40,10'd361};
ram[49462] = {-9'd37,10'd364};
ram[49463] = {-9'd33,10'd367};
ram[49464] = {-9'd30,10'd370};
ram[49465] = {-9'd27,10'd373};
ram[49466] = {-9'd24,10'd376};
ram[49467] = {-9'd21,10'd380};
ram[49468] = {-9'd18,10'd383};
ram[49469] = {-9'd15,10'd386};
ram[49470] = {-9'd11,10'd389};
ram[49471] = {-9'd8,10'd392};
ram[49472] = {-9'd5,10'd395};
ram[49473] = {-9'd2,10'd398};
ram[49474] = {9'd1,-10'd399};
ram[49475] = {9'd4,-10'd396};
ram[49476] = {9'd7,-10'd393};
ram[49477] = {9'd10,-10'd390};
ram[49478] = {9'd14,-10'd387};
ram[49479] = {9'd17,-10'd384};
ram[49480] = {9'd20,-10'd381};
ram[49481] = {9'd23,-10'd377};
ram[49482] = {9'd26,-10'd374};
ram[49483] = {9'd29,-10'd371};
ram[49484] = {9'd32,-10'd368};
ram[49485] = {9'd36,-10'd365};
ram[49486] = {9'd39,-10'd362};
ram[49487] = {9'd42,-10'd359};
ram[49488] = {9'd45,-10'd355};
ram[49489] = {9'd48,-10'd352};
ram[49490] = {9'd51,-10'd349};
ram[49491] = {9'd54,-10'd346};
ram[49492] = {9'd58,-10'd343};
ram[49493] = {9'd61,-10'd340};
ram[49494] = {9'd64,-10'd337};
ram[49495] = {9'd67,-10'd334};
ram[49496] = {9'd70,-10'd330};
ram[49497] = {9'd73,-10'd327};
ram[49498] = {9'd76,-10'd324};
ram[49499] = {9'd80,-10'd321};
ram[49500] = {9'd83,-10'd318};
ram[49501] = {9'd86,-10'd315};
ram[49502] = {9'd89,-10'd312};
ram[49503] = {9'd92,-10'd308};
ram[49504] = {9'd95,-10'd305};
ram[49505] = {9'd98,-10'd302};
ram[49506] = {-9'd99,-10'd299};
ram[49507] = {-9'd96,-10'd296};
ram[49508] = {-9'd92,-10'd293};
ram[49509] = {-9'd89,-10'd290};
ram[49510] = {-9'd86,-10'd286};
ram[49511] = {-9'd83,-10'd283};
ram[49512] = {-9'd80,-10'd280};
ram[49513] = {-9'd77,-10'd277};
ram[49514] = {-9'd74,-10'd274};
ram[49515] = {-9'd70,-10'd271};
ram[49516] = {-9'd67,-10'd268};
ram[49517] = {-9'd64,-10'd264};
ram[49518] = {-9'd61,-10'd261};
ram[49519] = {-9'd58,-10'd258};
ram[49520] = {-9'd55,-10'd255};
ram[49521] = {-9'd52,-10'd252};
ram[49522] = {-9'd48,-10'd249};
ram[49523] = {-9'd45,-10'd246};
ram[49524] = {-9'd42,-10'd242};
ram[49525] = {-9'd39,-10'd239};
ram[49526] = {-9'd36,-10'd236};
ram[49527] = {-9'd33,-10'd233};
ram[49528] = {-9'd30,-10'd230};
ram[49529] = {-9'd26,-10'd227};
ram[49530] = {-9'd23,-10'd224};
ram[49531] = {-9'd20,-10'd220};
ram[49532] = {-9'd17,-10'd217};
ram[49533] = {-9'd14,-10'd214};
ram[49534] = {-9'd11,-10'd211};
ram[49535] = {-9'd8,-10'd208};
ram[49536] = {-9'd8,-10'd208};
ram[49537] = {-9'd4,-10'd205};
ram[49538] = {-9'd1,-10'd202};
ram[49539] = {9'd2,-10'd198};
ram[49540] = {9'd5,-10'd195};
ram[49541] = {9'd8,-10'd192};
ram[49542] = {9'd11,-10'd189};
ram[49543] = {9'd14,-10'd186};
ram[49544] = {9'd18,-10'd183};
ram[49545] = {9'd21,-10'd180};
ram[49546] = {9'd24,-10'd176};
ram[49547] = {9'd27,-10'd173};
ram[49548] = {9'd30,-10'd170};
ram[49549] = {9'd33,-10'd167};
ram[49550] = {9'd36,-10'd164};
ram[49551] = {9'd40,-10'd161};
ram[49552] = {9'd43,-10'd158};
ram[49553] = {9'd46,-10'd154};
ram[49554] = {9'd49,-10'd151};
ram[49555] = {9'd52,-10'd148};
ram[49556] = {9'd55,-10'd145};
ram[49557] = {9'd58,-10'd142};
ram[49558] = {9'd62,-10'd139};
ram[49559] = {9'd65,-10'd136};
ram[49560] = {9'd68,-10'd132};
ram[49561] = {9'd71,-10'd129};
ram[49562] = {9'd74,-10'd126};
ram[49563] = {9'd77,-10'd123};
ram[49564] = {9'd80,-10'd120};
ram[49565] = {9'd84,-10'd117};
ram[49566] = {9'd87,-10'd114};
ram[49567] = {9'd90,-10'd110};
ram[49568] = {9'd93,-10'd107};
ram[49569] = {9'd96,-10'd104};
ram[49570] = {9'd99,-10'd101};
ram[49571] = {-9'd98,-10'd98};
ram[49572] = {-9'd95,-10'd95};
ram[49573] = {-9'd92,-10'd92};
ram[49574] = {-9'd88,-10'd88};
ram[49575] = {-9'd85,-10'd85};
ram[49576] = {-9'd82,-10'd82};
ram[49577] = {-9'd79,-10'd79};
ram[49578] = {-9'd76,-10'd76};
ram[49579] = {-9'd73,-10'd73};
ram[49580] = {-9'd70,-10'd70};
ram[49581] = {-9'd66,-10'd66};
ram[49582] = {-9'd63,-10'd63};
ram[49583] = {-9'd60,-10'd60};
ram[49584] = {-9'd57,-10'd57};
ram[49585] = {-9'd54,-10'd54};
ram[49586] = {-9'd51,-10'd51};
ram[49587] = {-9'd48,-10'd48};
ram[49588] = {-9'd44,-10'd44};
ram[49589] = {-9'd41,-10'd41};
ram[49590] = {-9'd38,-10'd38};
ram[49591] = {-9'd35,-10'd35};
ram[49592] = {-9'd32,-10'd32};
ram[49593] = {-9'd29,-10'd29};
ram[49594] = {-9'd26,-10'd26};
ram[49595] = {-9'd22,-10'd22};
ram[49596] = {-9'd19,-10'd19};
ram[49597] = {-9'd16,-10'd16};
ram[49598] = {-9'd13,-10'd13};
ram[49599] = {-9'd10,-10'd10};
ram[49600] = {-9'd7,-10'd7};
ram[49601] = {-9'd4,-10'd4};
ram[49602] = {9'd0,10'd0};
ram[49603] = {9'd3,10'd3};
ram[49604] = {9'd6,10'd6};
ram[49605] = {9'd9,10'd9};
ram[49606] = {9'd12,10'd12};
ram[49607] = {9'd15,10'd15};
ram[49608] = {9'd18,10'd18};
ram[49609] = {9'd21,10'd21};
ram[49610] = {9'd25,10'd25};
ram[49611] = {9'd28,10'd28};
ram[49612] = {9'd31,10'd31};
ram[49613] = {9'd34,10'd34};
ram[49614] = {9'd37,10'd37};
ram[49615] = {9'd40,10'd40};
ram[49616] = {9'd43,10'd43};
ram[49617] = {9'd47,10'd47};
ram[49618] = {9'd50,10'd50};
ram[49619] = {9'd53,10'd53};
ram[49620] = {9'd56,10'd56};
ram[49621] = {9'd59,10'd59};
ram[49622] = {9'd62,10'd62};
ram[49623] = {9'd65,10'd65};
ram[49624] = {9'd69,10'd69};
ram[49625] = {9'd72,10'd72};
ram[49626] = {9'd75,10'd75};
ram[49627] = {9'd78,10'd78};
ram[49628] = {9'd81,10'd81};
ram[49629] = {9'd84,10'd84};
ram[49630] = {9'd87,10'd87};
ram[49631] = {9'd91,10'd91};
ram[49632] = {9'd94,10'd94};
ram[49633] = {9'd97,10'd97};
ram[49634] = {-9'd100,10'd100};
ram[49635] = {-9'd97,10'd103};
ram[49636] = {-9'd94,10'd106};
ram[49637] = {-9'd91,10'd109};
ram[49638] = {-9'd88,10'd113};
ram[49639] = {-9'd85,10'd116};
ram[49640] = {-9'd81,10'd119};
ram[49641] = {-9'd78,10'd122};
ram[49642] = {-9'd75,10'd125};
ram[49643] = {-9'd72,10'd128};
ram[49644] = {-9'd69,10'd131};
ram[49645] = {-9'd66,10'd135};
ram[49646] = {-9'd63,10'd138};
ram[49647] = {-9'd59,10'd141};
ram[49648] = {-9'd56,10'd144};
ram[49649] = {-9'd53,10'd147};
ram[49650] = {-9'd50,10'd150};
ram[49651] = {-9'd47,10'd153};
ram[49652] = {-9'd44,10'd157};
ram[49653] = {-9'd41,10'd160};
ram[49654] = {-9'd37,10'd163};
ram[49655] = {-9'd34,10'd166};
ram[49656] = {-9'd31,10'd169};
ram[49657] = {-9'd28,10'd172};
ram[49658] = {-9'd25,10'd175};
ram[49659] = {-9'd22,10'd179};
ram[49660] = {-9'd19,10'd182};
ram[49661] = {-9'd15,10'd185};
ram[49662] = {-9'd12,10'd188};
ram[49663] = {-9'd9,10'd191};
ram[49664] = {-9'd9,10'd191};
ram[49665] = {-9'd6,10'd194};
ram[49666] = {-9'd3,10'd197};
ram[49667] = {9'd0,10'd201};
ram[49668] = {9'd3,10'd204};
ram[49669] = {9'd7,10'd207};
ram[49670] = {9'd10,10'd210};
ram[49671] = {9'd13,10'd213};
ram[49672] = {9'd16,10'd216};
ram[49673] = {9'd19,10'd219};
ram[49674] = {9'd22,10'd223};
ram[49675] = {9'd25,10'd226};
ram[49676] = {9'd29,10'd229};
ram[49677] = {9'd32,10'd232};
ram[49678] = {9'd35,10'd235};
ram[49679] = {9'd38,10'd238};
ram[49680] = {9'd41,10'd241};
ram[49681] = {9'd44,10'd245};
ram[49682] = {9'd47,10'd248};
ram[49683] = {9'd51,10'd251};
ram[49684] = {9'd54,10'd254};
ram[49685] = {9'd57,10'd257};
ram[49686] = {9'd60,10'd260};
ram[49687] = {9'd63,10'd263};
ram[49688] = {9'd66,10'd267};
ram[49689] = {9'd69,10'd270};
ram[49690] = {9'd73,10'd273};
ram[49691] = {9'd76,10'd276};
ram[49692] = {9'd79,10'd279};
ram[49693] = {9'd82,10'd282};
ram[49694] = {9'd85,10'd285};
ram[49695] = {9'd88,10'd289};
ram[49696] = {9'd91,10'd292};
ram[49697] = {9'd95,10'd295};
ram[49698] = {9'd98,10'd298};
ram[49699] = {-9'd99,10'd301};
ram[49700] = {-9'd96,10'd304};
ram[49701] = {-9'd93,10'd307};
ram[49702] = {-9'd90,10'd311};
ram[49703] = {-9'd87,10'd314};
ram[49704] = {-9'd84,10'd317};
ram[49705] = {-9'd81,10'd320};
ram[49706] = {-9'd77,10'd323};
ram[49707] = {-9'd74,10'd326};
ram[49708] = {-9'd71,10'd329};
ram[49709] = {-9'd68,10'd333};
ram[49710] = {-9'd65,10'd336};
ram[49711] = {-9'd62,10'd339};
ram[49712] = {-9'd59,10'd342};
ram[49713] = {-9'd55,10'd345};
ram[49714] = {-9'd52,10'd348};
ram[49715] = {-9'd49,10'd351};
ram[49716] = {-9'd46,10'd354};
ram[49717] = {-9'd43,10'd358};
ram[49718] = {-9'd40,10'd361};
ram[49719] = {-9'd37,10'd364};
ram[49720] = {-9'd33,10'd367};
ram[49721] = {-9'd30,10'd370};
ram[49722] = {-9'd27,10'd373};
ram[49723] = {-9'd24,10'd376};
ram[49724] = {-9'd21,10'd380};
ram[49725] = {-9'd18,10'd383};
ram[49726] = {-9'd15,10'd386};
ram[49727] = {-9'd11,10'd389};
ram[49728] = {-9'd8,10'd392};
ram[49729] = {-9'd5,10'd395};
ram[49730] = {-9'd2,10'd398};
ram[49731] = {9'd1,-10'd399};
ram[49732] = {9'd4,-10'd396};
ram[49733] = {9'd7,-10'd393};
ram[49734] = {9'd10,-10'd390};
ram[49735] = {9'd14,-10'd387};
ram[49736] = {9'd17,-10'd384};
ram[49737] = {9'd20,-10'd381};
ram[49738] = {9'd23,-10'd377};
ram[49739] = {9'd26,-10'd374};
ram[49740] = {9'd29,-10'd371};
ram[49741] = {9'd32,-10'd368};
ram[49742] = {9'd36,-10'd365};
ram[49743] = {9'd39,-10'd362};
ram[49744] = {9'd42,-10'd359};
ram[49745] = {9'd45,-10'd355};
ram[49746] = {9'd48,-10'd352};
ram[49747] = {9'd51,-10'd349};
ram[49748] = {9'd54,-10'd346};
ram[49749] = {9'd58,-10'd343};
ram[49750] = {9'd61,-10'd340};
ram[49751] = {9'd64,-10'd337};
ram[49752] = {9'd67,-10'd334};
ram[49753] = {9'd70,-10'd330};
ram[49754] = {9'd73,-10'd327};
ram[49755] = {9'd76,-10'd324};
ram[49756] = {9'd80,-10'd321};
ram[49757] = {9'd83,-10'd318};
ram[49758] = {9'd86,-10'd315};
ram[49759] = {9'd89,-10'd312};
ram[49760] = {9'd92,-10'd308};
ram[49761] = {9'd95,-10'd305};
ram[49762] = {9'd98,-10'd302};
ram[49763] = {-9'd99,-10'd299};
ram[49764] = {-9'd96,-10'd296};
ram[49765] = {-9'd92,-10'd293};
ram[49766] = {-9'd89,-10'd290};
ram[49767] = {-9'd86,-10'd286};
ram[49768] = {-9'd83,-10'd283};
ram[49769] = {-9'd80,-10'd280};
ram[49770] = {-9'd77,-10'd277};
ram[49771] = {-9'd74,-10'd274};
ram[49772] = {-9'd70,-10'd271};
ram[49773] = {-9'd67,-10'd268};
ram[49774] = {-9'd64,-10'd264};
ram[49775] = {-9'd61,-10'd261};
ram[49776] = {-9'd58,-10'd258};
ram[49777] = {-9'd55,-10'd255};
ram[49778] = {-9'd52,-10'd252};
ram[49779] = {-9'd48,-10'd249};
ram[49780] = {-9'd45,-10'd246};
ram[49781] = {-9'd42,-10'd242};
ram[49782] = {-9'd39,-10'd239};
ram[49783] = {-9'd36,-10'd236};
ram[49784] = {-9'd33,-10'd233};
ram[49785] = {-9'd30,-10'd230};
ram[49786] = {-9'd26,-10'd227};
ram[49787] = {-9'd23,-10'd224};
ram[49788] = {-9'd20,-10'd220};
ram[49789] = {-9'd17,-10'd217};
ram[49790] = {-9'd14,-10'd214};
ram[49791] = {-9'd11,-10'd211};
ram[49792] = {-9'd11,-10'd211};
ram[49793] = {-9'd8,-10'd208};
ram[49794] = {-9'd4,-10'd205};
ram[49795] = {-9'd1,-10'd202};
ram[49796] = {9'd2,-10'd198};
ram[49797] = {9'd5,-10'd195};
ram[49798] = {9'd8,-10'd192};
ram[49799] = {9'd11,-10'd189};
ram[49800] = {9'd14,-10'd186};
ram[49801] = {9'd18,-10'd183};
ram[49802] = {9'd21,-10'd180};
ram[49803] = {9'd24,-10'd176};
ram[49804] = {9'd27,-10'd173};
ram[49805] = {9'd30,-10'd170};
ram[49806] = {9'd33,-10'd167};
ram[49807] = {9'd36,-10'd164};
ram[49808] = {9'd40,-10'd161};
ram[49809] = {9'd43,-10'd158};
ram[49810] = {9'd46,-10'd154};
ram[49811] = {9'd49,-10'd151};
ram[49812] = {9'd52,-10'd148};
ram[49813] = {9'd55,-10'd145};
ram[49814] = {9'd58,-10'd142};
ram[49815] = {9'd62,-10'd139};
ram[49816] = {9'd65,-10'd136};
ram[49817] = {9'd68,-10'd132};
ram[49818] = {9'd71,-10'd129};
ram[49819] = {9'd74,-10'd126};
ram[49820] = {9'd77,-10'd123};
ram[49821] = {9'd80,-10'd120};
ram[49822] = {9'd84,-10'd117};
ram[49823] = {9'd87,-10'd114};
ram[49824] = {9'd90,-10'd110};
ram[49825] = {9'd93,-10'd107};
ram[49826] = {9'd96,-10'd104};
ram[49827] = {9'd99,-10'd101};
ram[49828] = {-9'd98,-10'd98};
ram[49829] = {-9'd95,-10'd95};
ram[49830] = {-9'd92,-10'd92};
ram[49831] = {-9'd88,-10'd88};
ram[49832] = {-9'd85,-10'd85};
ram[49833] = {-9'd82,-10'd82};
ram[49834] = {-9'd79,-10'd79};
ram[49835] = {-9'd76,-10'd76};
ram[49836] = {-9'd73,-10'd73};
ram[49837] = {-9'd70,-10'd70};
ram[49838] = {-9'd66,-10'd66};
ram[49839] = {-9'd63,-10'd63};
ram[49840] = {-9'd60,-10'd60};
ram[49841] = {-9'd57,-10'd57};
ram[49842] = {-9'd54,-10'd54};
ram[49843] = {-9'd51,-10'd51};
ram[49844] = {-9'd48,-10'd48};
ram[49845] = {-9'd44,-10'd44};
ram[49846] = {-9'd41,-10'd41};
ram[49847] = {-9'd38,-10'd38};
ram[49848] = {-9'd35,-10'd35};
ram[49849] = {-9'd32,-10'd32};
ram[49850] = {-9'd29,-10'd29};
ram[49851] = {-9'd26,-10'd26};
ram[49852] = {-9'd22,-10'd22};
ram[49853] = {-9'd19,-10'd19};
ram[49854] = {-9'd16,-10'd16};
ram[49855] = {-9'd13,-10'd13};
ram[49856] = {-9'd10,-10'd10};
ram[49857] = {-9'd7,-10'd7};
ram[49858] = {-9'd4,-10'd4};
ram[49859] = {9'd0,10'd0};
ram[49860] = {9'd3,10'd3};
ram[49861] = {9'd6,10'd6};
ram[49862] = {9'd9,10'd9};
ram[49863] = {9'd12,10'd12};
ram[49864] = {9'd15,10'd15};
ram[49865] = {9'd18,10'd18};
ram[49866] = {9'd21,10'd21};
ram[49867] = {9'd25,10'd25};
ram[49868] = {9'd28,10'd28};
ram[49869] = {9'd31,10'd31};
ram[49870] = {9'd34,10'd34};
ram[49871] = {9'd37,10'd37};
ram[49872] = {9'd40,10'd40};
ram[49873] = {9'd43,10'd43};
ram[49874] = {9'd47,10'd47};
ram[49875] = {9'd50,10'd50};
ram[49876] = {9'd53,10'd53};
ram[49877] = {9'd56,10'd56};
ram[49878] = {9'd59,10'd59};
ram[49879] = {9'd62,10'd62};
ram[49880] = {9'd65,10'd65};
ram[49881] = {9'd69,10'd69};
ram[49882] = {9'd72,10'd72};
ram[49883] = {9'd75,10'd75};
ram[49884] = {9'd78,10'd78};
ram[49885] = {9'd81,10'd81};
ram[49886] = {9'd84,10'd84};
ram[49887] = {9'd87,10'd87};
ram[49888] = {9'd91,10'd91};
ram[49889] = {9'd94,10'd94};
ram[49890] = {9'd97,10'd97};
ram[49891] = {-9'd100,10'd100};
ram[49892] = {-9'd97,10'd103};
ram[49893] = {-9'd94,10'd106};
ram[49894] = {-9'd91,10'd109};
ram[49895] = {-9'd88,10'd113};
ram[49896] = {-9'd85,10'd116};
ram[49897] = {-9'd81,10'd119};
ram[49898] = {-9'd78,10'd122};
ram[49899] = {-9'd75,10'd125};
ram[49900] = {-9'd72,10'd128};
ram[49901] = {-9'd69,10'd131};
ram[49902] = {-9'd66,10'd135};
ram[49903] = {-9'd63,10'd138};
ram[49904] = {-9'd59,10'd141};
ram[49905] = {-9'd56,10'd144};
ram[49906] = {-9'd53,10'd147};
ram[49907] = {-9'd50,10'd150};
ram[49908] = {-9'd47,10'd153};
ram[49909] = {-9'd44,10'd157};
ram[49910] = {-9'd41,10'd160};
ram[49911] = {-9'd37,10'd163};
ram[49912] = {-9'd34,10'd166};
ram[49913] = {-9'd31,10'd169};
ram[49914] = {-9'd28,10'd172};
ram[49915] = {-9'd25,10'd175};
ram[49916] = {-9'd22,10'd179};
ram[49917] = {-9'd19,10'd182};
ram[49918] = {-9'd15,10'd185};
ram[49919] = {-9'd12,10'd188};
ram[49920] = {-9'd12,10'd188};
ram[49921] = {-9'd9,10'd191};
ram[49922] = {-9'd6,10'd194};
ram[49923] = {-9'd3,10'd197};
ram[49924] = {9'd0,10'd201};
ram[49925] = {9'd3,10'd204};
ram[49926] = {9'd7,10'd207};
ram[49927] = {9'd10,10'd210};
ram[49928] = {9'd13,10'd213};
ram[49929] = {9'd16,10'd216};
ram[49930] = {9'd19,10'd219};
ram[49931] = {9'd22,10'd223};
ram[49932] = {9'd25,10'd226};
ram[49933] = {9'd29,10'd229};
ram[49934] = {9'd32,10'd232};
ram[49935] = {9'd35,10'd235};
ram[49936] = {9'd38,10'd238};
ram[49937] = {9'd41,10'd241};
ram[49938] = {9'd44,10'd245};
ram[49939] = {9'd47,10'd248};
ram[49940] = {9'd51,10'd251};
ram[49941] = {9'd54,10'd254};
ram[49942] = {9'd57,10'd257};
ram[49943] = {9'd60,10'd260};
ram[49944] = {9'd63,10'd263};
ram[49945] = {9'd66,10'd267};
ram[49946] = {9'd69,10'd270};
ram[49947] = {9'd73,10'd273};
ram[49948] = {9'd76,10'd276};
ram[49949] = {9'd79,10'd279};
ram[49950] = {9'd82,10'd282};
ram[49951] = {9'd85,10'd285};
ram[49952] = {9'd88,10'd289};
ram[49953] = {9'd91,10'd292};
ram[49954] = {9'd95,10'd295};
ram[49955] = {9'd98,10'd298};
ram[49956] = {-9'd99,10'd301};
ram[49957] = {-9'd96,10'd304};
ram[49958] = {-9'd93,10'd307};
ram[49959] = {-9'd90,10'd311};
ram[49960] = {-9'd87,10'd314};
ram[49961] = {-9'd84,10'd317};
ram[49962] = {-9'd81,10'd320};
ram[49963] = {-9'd77,10'd323};
ram[49964] = {-9'd74,10'd326};
ram[49965] = {-9'd71,10'd329};
ram[49966] = {-9'd68,10'd333};
ram[49967] = {-9'd65,10'd336};
ram[49968] = {-9'd62,10'd339};
ram[49969] = {-9'd59,10'd342};
ram[49970] = {-9'd55,10'd345};
ram[49971] = {-9'd52,10'd348};
ram[49972] = {-9'd49,10'd351};
ram[49973] = {-9'd46,10'd354};
ram[49974] = {-9'd43,10'd358};
ram[49975] = {-9'd40,10'd361};
ram[49976] = {-9'd37,10'd364};
ram[49977] = {-9'd33,10'd367};
ram[49978] = {-9'd30,10'd370};
ram[49979] = {-9'd27,10'd373};
ram[49980] = {-9'd24,10'd376};
ram[49981] = {-9'd21,10'd380};
ram[49982] = {-9'd18,10'd383};
ram[49983] = {-9'd15,10'd386};
ram[49984] = {-9'd11,10'd389};
ram[49985] = {-9'd8,10'd392};
ram[49986] = {-9'd5,10'd395};
ram[49987] = {-9'd2,10'd398};
ram[49988] = {9'd1,-10'd399};
ram[49989] = {9'd4,-10'd396};
ram[49990] = {9'd7,-10'd393};
ram[49991] = {9'd10,-10'd390};
ram[49992] = {9'd14,-10'd387};
ram[49993] = {9'd17,-10'd384};
ram[49994] = {9'd20,-10'd381};
ram[49995] = {9'd23,-10'd377};
ram[49996] = {9'd26,-10'd374};
ram[49997] = {9'd29,-10'd371};
ram[49998] = {9'd32,-10'd368};
ram[49999] = {9'd36,-10'd365};
ram[50000] = {9'd39,-10'd362};
ram[50001] = {9'd42,-10'd359};
ram[50002] = {9'd45,-10'd355};
ram[50003] = {9'd48,-10'd352};
ram[50004] = {9'd51,-10'd349};
ram[50005] = {9'd54,-10'd346};
ram[50006] = {9'd58,-10'd343};
ram[50007] = {9'd61,-10'd340};
ram[50008] = {9'd64,-10'd337};
ram[50009] = {9'd67,-10'd334};
ram[50010] = {9'd70,-10'd330};
ram[50011] = {9'd73,-10'd327};
ram[50012] = {9'd76,-10'd324};
ram[50013] = {9'd80,-10'd321};
ram[50014] = {9'd83,-10'd318};
ram[50015] = {9'd86,-10'd315};
ram[50016] = {9'd89,-10'd312};
ram[50017] = {9'd92,-10'd308};
ram[50018] = {9'd95,-10'd305};
ram[50019] = {9'd98,-10'd302};
ram[50020] = {-9'd99,-10'd299};
ram[50021] = {-9'd96,-10'd296};
ram[50022] = {-9'd92,-10'd293};
ram[50023] = {-9'd89,-10'd290};
ram[50024] = {-9'd86,-10'd286};
ram[50025] = {-9'd83,-10'd283};
ram[50026] = {-9'd80,-10'd280};
ram[50027] = {-9'd77,-10'd277};
ram[50028] = {-9'd74,-10'd274};
ram[50029] = {-9'd70,-10'd271};
ram[50030] = {-9'd67,-10'd268};
ram[50031] = {-9'd64,-10'd264};
ram[50032] = {-9'd61,-10'd261};
ram[50033] = {-9'd58,-10'd258};
ram[50034] = {-9'd55,-10'd255};
ram[50035] = {-9'd52,-10'd252};
ram[50036] = {-9'd48,-10'd249};
ram[50037] = {-9'd45,-10'd246};
ram[50038] = {-9'd42,-10'd242};
ram[50039] = {-9'd39,-10'd239};
ram[50040] = {-9'd36,-10'd236};
ram[50041] = {-9'd33,-10'd233};
ram[50042] = {-9'd30,-10'd230};
ram[50043] = {-9'd26,-10'd227};
ram[50044] = {-9'd23,-10'd224};
ram[50045] = {-9'd20,-10'd220};
ram[50046] = {-9'd17,-10'd217};
ram[50047] = {-9'd14,-10'd214};
ram[50048] = {-9'd14,-10'd214};
ram[50049] = {-9'd11,-10'd211};
ram[50050] = {-9'd8,-10'd208};
ram[50051] = {-9'd4,-10'd205};
ram[50052] = {-9'd1,-10'd202};
ram[50053] = {9'd2,-10'd198};
ram[50054] = {9'd5,-10'd195};
ram[50055] = {9'd8,-10'd192};
ram[50056] = {9'd11,-10'd189};
ram[50057] = {9'd14,-10'd186};
ram[50058] = {9'd18,-10'd183};
ram[50059] = {9'd21,-10'd180};
ram[50060] = {9'd24,-10'd176};
ram[50061] = {9'd27,-10'd173};
ram[50062] = {9'd30,-10'd170};
ram[50063] = {9'd33,-10'd167};
ram[50064] = {9'd36,-10'd164};
ram[50065] = {9'd40,-10'd161};
ram[50066] = {9'd43,-10'd158};
ram[50067] = {9'd46,-10'd154};
ram[50068] = {9'd49,-10'd151};
ram[50069] = {9'd52,-10'd148};
ram[50070] = {9'd55,-10'd145};
ram[50071] = {9'd58,-10'd142};
ram[50072] = {9'd62,-10'd139};
ram[50073] = {9'd65,-10'd136};
ram[50074] = {9'd68,-10'd132};
ram[50075] = {9'd71,-10'd129};
ram[50076] = {9'd74,-10'd126};
ram[50077] = {9'd77,-10'd123};
ram[50078] = {9'd80,-10'd120};
ram[50079] = {9'd84,-10'd117};
ram[50080] = {9'd87,-10'd114};
ram[50081] = {9'd90,-10'd110};
ram[50082] = {9'd93,-10'd107};
ram[50083] = {9'd96,-10'd104};
ram[50084] = {9'd99,-10'd101};
ram[50085] = {-9'd98,-10'd98};
ram[50086] = {-9'd95,-10'd95};
ram[50087] = {-9'd92,-10'd92};
ram[50088] = {-9'd88,-10'd88};
ram[50089] = {-9'd85,-10'd85};
ram[50090] = {-9'd82,-10'd82};
ram[50091] = {-9'd79,-10'd79};
ram[50092] = {-9'd76,-10'd76};
ram[50093] = {-9'd73,-10'd73};
ram[50094] = {-9'd70,-10'd70};
ram[50095] = {-9'd66,-10'd66};
ram[50096] = {-9'd63,-10'd63};
ram[50097] = {-9'd60,-10'd60};
ram[50098] = {-9'd57,-10'd57};
ram[50099] = {-9'd54,-10'd54};
ram[50100] = {-9'd51,-10'd51};
ram[50101] = {-9'd48,-10'd48};
ram[50102] = {-9'd44,-10'd44};
ram[50103] = {-9'd41,-10'd41};
ram[50104] = {-9'd38,-10'd38};
ram[50105] = {-9'd35,-10'd35};
ram[50106] = {-9'd32,-10'd32};
ram[50107] = {-9'd29,-10'd29};
ram[50108] = {-9'd26,-10'd26};
ram[50109] = {-9'd22,-10'd22};
ram[50110] = {-9'd19,-10'd19};
ram[50111] = {-9'd16,-10'd16};
ram[50112] = {-9'd13,-10'd13};
ram[50113] = {-9'd10,-10'd10};
ram[50114] = {-9'd7,-10'd7};
ram[50115] = {-9'd4,-10'd4};
ram[50116] = {9'd0,10'd0};
ram[50117] = {9'd3,10'd3};
ram[50118] = {9'd6,10'd6};
ram[50119] = {9'd9,10'd9};
ram[50120] = {9'd12,10'd12};
ram[50121] = {9'd15,10'd15};
ram[50122] = {9'd18,10'd18};
ram[50123] = {9'd21,10'd21};
ram[50124] = {9'd25,10'd25};
ram[50125] = {9'd28,10'd28};
ram[50126] = {9'd31,10'd31};
ram[50127] = {9'd34,10'd34};
ram[50128] = {9'd37,10'd37};
ram[50129] = {9'd40,10'd40};
ram[50130] = {9'd43,10'd43};
ram[50131] = {9'd47,10'd47};
ram[50132] = {9'd50,10'd50};
ram[50133] = {9'd53,10'd53};
ram[50134] = {9'd56,10'd56};
ram[50135] = {9'd59,10'd59};
ram[50136] = {9'd62,10'd62};
ram[50137] = {9'd65,10'd65};
ram[50138] = {9'd69,10'd69};
ram[50139] = {9'd72,10'd72};
ram[50140] = {9'd75,10'd75};
ram[50141] = {9'd78,10'd78};
ram[50142] = {9'd81,10'd81};
ram[50143] = {9'd84,10'd84};
ram[50144] = {9'd87,10'd87};
ram[50145] = {9'd91,10'd91};
ram[50146] = {9'd94,10'd94};
ram[50147] = {9'd97,10'd97};
ram[50148] = {-9'd100,10'd100};
ram[50149] = {-9'd97,10'd103};
ram[50150] = {-9'd94,10'd106};
ram[50151] = {-9'd91,10'd109};
ram[50152] = {-9'd88,10'd113};
ram[50153] = {-9'd85,10'd116};
ram[50154] = {-9'd81,10'd119};
ram[50155] = {-9'd78,10'd122};
ram[50156] = {-9'd75,10'd125};
ram[50157] = {-9'd72,10'd128};
ram[50158] = {-9'd69,10'd131};
ram[50159] = {-9'd66,10'd135};
ram[50160] = {-9'd63,10'd138};
ram[50161] = {-9'd59,10'd141};
ram[50162] = {-9'd56,10'd144};
ram[50163] = {-9'd53,10'd147};
ram[50164] = {-9'd50,10'd150};
ram[50165] = {-9'd47,10'd153};
ram[50166] = {-9'd44,10'd157};
ram[50167] = {-9'd41,10'd160};
ram[50168] = {-9'd37,10'd163};
ram[50169] = {-9'd34,10'd166};
ram[50170] = {-9'd31,10'd169};
ram[50171] = {-9'd28,10'd172};
ram[50172] = {-9'd25,10'd175};
ram[50173] = {-9'd22,10'd179};
ram[50174] = {-9'd19,10'd182};
ram[50175] = {-9'd15,10'd185};
ram[50176] = {-9'd15,10'd185};
ram[50177] = {-9'd12,10'd188};
ram[50178] = {-9'd9,10'd191};
ram[50179] = {-9'd6,10'd194};
ram[50180] = {-9'd3,10'd197};
ram[50181] = {9'd0,10'd201};
ram[50182] = {9'd3,10'd204};
ram[50183] = {9'd7,10'd207};
ram[50184] = {9'd10,10'd210};
ram[50185] = {9'd13,10'd213};
ram[50186] = {9'd16,10'd216};
ram[50187] = {9'd19,10'd219};
ram[50188] = {9'd22,10'd223};
ram[50189] = {9'd25,10'd226};
ram[50190] = {9'd29,10'd229};
ram[50191] = {9'd32,10'd232};
ram[50192] = {9'd35,10'd235};
ram[50193] = {9'd38,10'd238};
ram[50194] = {9'd41,10'd241};
ram[50195] = {9'd44,10'd245};
ram[50196] = {9'd47,10'd248};
ram[50197] = {9'd51,10'd251};
ram[50198] = {9'd54,10'd254};
ram[50199] = {9'd57,10'd257};
ram[50200] = {9'd60,10'd260};
ram[50201] = {9'd63,10'd263};
ram[50202] = {9'd66,10'd267};
ram[50203] = {9'd69,10'd270};
ram[50204] = {9'd73,10'd273};
ram[50205] = {9'd76,10'd276};
ram[50206] = {9'd79,10'd279};
ram[50207] = {9'd82,10'd282};
ram[50208] = {9'd85,10'd285};
ram[50209] = {9'd88,10'd289};
ram[50210] = {9'd91,10'd292};
ram[50211] = {9'd95,10'd295};
ram[50212] = {9'd98,10'd298};
ram[50213] = {-9'd99,10'd301};
ram[50214] = {-9'd96,10'd304};
ram[50215] = {-9'd93,10'd307};
ram[50216] = {-9'd90,10'd311};
ram[50217] = {-9'd87,10'd314};
ram[50218] = {-9'd84,10'd317};
ram[50219] = {-9'd81,10'd320};
ram[50220] = {-9'd77,10'd323};
ram[50221] = {-9'd74,10'd326};
ram[50222] = {-9'd71,10'd329};
ram[50223] = {-9'd68,10'd333};
ram[50224] = {-9'd65,10'd336};
ram[50225] = {-9'd62,10'd339};
ram[50226] = {-9'd59,10'd342};
ram[50227] = {-9'd55,10'd345};
ram[50228] = {-9'd52,10'd348};
ram[50229] = {-9'd49,10'd351};
ram[50230] = {-9'd46,10'd354};
ram[50231] = {-9'd43,10'd358};
ram[50232] = {-9'd40,10'd361};
ram[50233] = {-9'd37,10'd364};
ram[50234] = {-9'd33,10'd367};
ram[50235] = {-9'd30,10'd370};
ram[50236] = {-9'd27,10'd373};
ram[50237] = {-9'd24,10'd376};
ram[50238] = {-9'd21,10'd380};
ram[50239] = {-9'd18,10'd383};
ram[50240] = {-9'd15,10'd386};
ram[50241] = {-9'd11,10'd389};
ram[50242] = {-9'd8,10'd392};
ram[50243] = {-9'd5,10'd395};
ram[50244] = {-9'd2,10'd398};
ram[50245] = {9'd1,-10'd399};
ram[50246] = {9'd4,-10'd396};
ram[50247] = {9'd7,-10'd393};
ram[50248] = {9'd10,-10'd390};
ram[50249] = {9'd14,-10'd387};
ram[50250] = {9'd17,-10'd384};
ram[50251] = {9'd20,-10'd381};
ram[50252] = {9'd23,-10'd377};
ram[50253] = {9'd26,-10'd374};
ram[50254] = {9'd29,-10'd371};
ram[50255] = {9'd32,-10'd368};
ram[50256] = {9'd36,-10'd365};
ram[50257] = {9'd39,-10'd362};
ram[50258] = {9'd42,-10'd359};
ram[50259] = {9'd45,-10'd355};
ram[50260] = {9'd48,-10'd352};
ram[50261] = {9'd51,-10'd349};
ram[50262] = {9'd54,-10'd346};
ram[50263] = {9'd58,-10'd343};
ram[50264] = {9'd61,-10'd340};
ram[50265] = {9'd64,-10'd337};
ram[50266] = {9'd67,-10'd334};
ram[50267] = {9'd70,-10'd330};
ram[50268] = {9'd73,-10'd327};
ram[50269] = {9'd76,-10'd324};
ram[50270] = {9'd80,-10'd321};
ram[50271] = {9'd83,-10'd318};
ram[50272] = {9'd86,-10'd315};
ram[50273] = {9'd89,-10'd312};
ram[50274] = {9'd92,-10'd308};
ram[50275] = {9'd95,-10'd305};
ram[50276] = {9'd98,-10'd302};
ram[50277] = {-9'd99,-10'd299};
ram[50278] = {-9'd96,-10'd296};
ram[50279] = {-9'd92,-10'd293};
ram[50280] = {-9'd89,-10'd290};
ram[50281] = {-9'd86,-10'd286};
ram[50282] = {-9'd83,-10'd283};
ram[50283] = {-9'd80,-10'd280};
ram[50284] = {-9'd77,-10'd277};
ram[50285] = {-9'd74,-10'd274};
ram[50286] = {-9'd70,-10'd271};
ram[50287] = {-9'd67,-10'd268};
ram[50288] = {-9'd64,-10'd264};
ram[50289] = {-9'd61,-10'd261};
ram[50290] = {-9'd58,-10'd258};
ram[50291] = {-9'd55,-10'd255};
ram[50292] = {-9'd52,-10'd252};
ram[50293] = {-9'd48,-10'd249};
ram[50294] = {-9'd45,-10'd246};
ram[50295] = {-9'd42,-10'd242};
ram[50296] = {-9'd39,-10'd239};
ram[50297] = {-9'd36,-10'd236};
ram[50298] = {-9'd33,-10'd233};
ram[50299] = {-9'd30,-10'd230};
ram[50300] = {-9'd26,-10'd227};
ram[50301] = {-9'd23,-10'd224};
ram[50302] = {-9'd20,-10'd220};
ram[50303] = {-9'd17,-10'd217};
ram[50304] = {-9'd17,-10'd217};
ram[50305] = {-9'd14,-10'd214};
ram[50306] = {-9'd11,-10'd211};
ram[50307] = {-9'd8,-10'd208};
ram[50308] = {-9'd4,-10'd205};
ram[50309] = {-9'd1,-10'd202};
ram[50310] = {9'd2,-10'd198};
ram[50311] = {9'd5,-10'd195};
ram[50312] = {9'd8,-10'd192};
ram[50313] = {9'd11,-10'd189};
ram[50314] = {9'd14,-10'd186};
ram[50315] = {9'd18,-10'd183};
ram[50316] = {9'd21,-10'd180};
ram[50317] = {9'd24,-10'd176};
ram[50318] = {9'd27,-10'd173};
ram[50319] = {9'd30,-10'd170};
ram[50320] = {9'd33,-10'd167};
ram[50321] = {9'd36,-10'd164};
ram[50322] = {9'd40,-10'd161};
ram[50323] = {9'd43,-10'd158};
ram[50324] = {9'd46,-10'd154};
ram[50325] = {9'd49,-10'd151};
ram[50326] = {9'd52,-10'd148};
ram[50327] = {9'd55,-10'd145};
ram[50328] = {9'd58,-10'd142};
ram[50329] = {9'd62,-10'd139};
ram[50330] = {9'd65,-10'd136};
ram[50331] = {9'd68,-10'd132};
ram[50332] = {9'd71,-10'd129};
ram[50333] = {9'd74,-10'd126};
ram[50334] = {9'd77,-10'd123};
ram[50335] = {9'd80,-10'd120};
ram[50336] = {9'd84,-10'd117};
ram[50337] = {9'd87,-10'd114};
ram[50338] = {9'd90,-10'd110};
ram[50339] = {9'd93,-10'd107};
ram[50340] = {9'd96,-10'd104};
ram[50341] = {9'd99,-10'd101};
ram[50342] = {-9'd98,-10'd98};
ram[50343] = {-9'd95,-10'd95};
ram[50344] = {-9'd92,-10'd92};
ram[50345] = {-9'd88,-10'd88};
ram[50346] = {-9'd85,-10'd85};
ram[50347] = {-9'd82,-10'd82};
ram[50348] = {-9'd79,-10'd79};
ram[50349] = {-9'd76,-10'd76};
ram[50350] = {-9'd73,-10'd73};
ram[50351] = {-9'd70,-10'd70};
ram[50352] = {-9'd66,-10'd66};
ram[50353] = {-9'd63,-10'd63};
ram[50354] = {-9'd60,-10'd60};
ram[50355] = {-9'd57,-10'd57};
ram[50356] = {-9'd54,-10'd54};
ram[50357] = {-9'd51,-10'd51};
ram[50358] = {-9'd48,-10'd48};
ram[50359] = {-9'd44,-10'd44};
ram[50360] = {-9'd41,-10'd41};
ram[50361] = {-9'd38,-10'd38};
ram[50362] = {-9'd35,-10'd35};
ram[50363] = {-9'd32,-10'd32};
ram[50364] = {-9'd29,-10'd29};
ram[50365] = {-9'd26,-10'd26};
ram[50366] = {-9'd22,-10'd22};
ram[50367] = {-9'd19,-10'd19};
ram[50368] = {-9'd16,-10'd16};
ram[50369] = {-9'd13,-10'd13};
ram[50370] = {-9'd10,-10'd10};
ram[50371] = {-9'd7,-10'd7};
ram[50372] = {-9'd4,-10'd4};
ram[50373] = {9'd0,10'd0};
ram[50374] = {9'd3,10'd3};
ram[50375] = {9'd6,10'd6};
ram[50376] = {9'd9,10'd9};
ram[50377] = {9'd12,10'd12};
ram[50378] = {9'd15,10'd15};
ram[50379] = {9'd18,10'd18};
ram[50380] = {9'd21,10'd21};
ram[50381] = {9'd25,10'd25};
ram[50382] = {9'd28,10'd28};
ram[50383] = {9'd31,10'd31};
ram[50384] = {9'd34,10'd34};
ram[50385] = {9'd37,10'd37};
ram[50386] = {9'd40,10'd40};
ram[50387] = {9'd43,10'd43};
ram[50388] = {9'd47,10'd47};
ram[50389] = {9'd50,10'd50};
ram[50390] = {9'd53,10'd53};
ram[50391] = {9'd56,10'd56};
ram[50392] = {9'd59,10'd59};
ram[50393] = {9'd62,10'd62};
ram[50394] = {9'd65,10'd65};
ram[50395] = {9'd69,10'd69};
ram[50396] = {9'd72,10'd72};
ram[50397] = {9'd75,10'd75};
ram[50398] = {9'd78,10'd78};
ram[50399] = {9'd81,10'd81};
ram[50400] = {9'd84,10'd84};
ram[50401] = {9'd87,10'd87};
ram[50402] = {9'd91,10'd91};
ram[50403] = {9'd94,10'd94};
ram[50404] = {9'd97,10'd97};
ram[50405] = {-9'd100,10'd100};
ram[50406] = {-9'd97,10'd103};
ram[50407] = {-9'd94,10'd106};
ram[50408] = {-9'd91,10'd109};
ram[50409] = {-9'd88,10'd113};
ram[50410] = {-9'd85,10'd116};
ram[50411] = {-9'd81,10'd119};
ram[50412] = {-9'd78,10'd122};
ram[50413] = {-9'd75,10'd125};
ram[50414] = {-9'd72,10'd128};
ram[50415] = {-9'd69,10'd131};
ram[50416] = {-9'd66,10'd135};
ram[50417] = {-9'd63,10'd138};
ram[50418] = {-9'd59,10'd141};
ram[50419] = {-9'd56,10'd144};
ram[50420] = {-9'd53,10'd147};
ram[50421] = {-9'd50,10'd150};
ram[50422] = {-9'd47,10'd153};
ram[50423] = {-9'd44,10'd157};
ram[50424] = {-9'd41,10'd160};
ram[50425] = {-9'd37,10'd163};
ram[50426] = {-9'd34,10'd166};
ram[50427] = {-9'd31,10'd169};
ram[50428] = {-9'd28,10'd172};
ram[50429] = {-9'd25,10'd175};
ram[50430] = {-9'd22,10'd179};
ram[50431] = {-9'd19,10'd182};
ram[50432] = {-9'd19,10'd182};
ram[50433] = {-9'd15,10'd185};
ram[50434] = {-9'd12,10'd188};
ram[50435] = {-9'd9,10'd191};
ram[50436] = {-9'd6,10'd194};
ram[50437] = {-9'd3,10'd197};
ram[50438] = {9'd0,10'd201};
ram[50439] = {9'd3,10'd204};
ram[50440] = {9'd7,10'd207};
ram[50441] = {9'd10,10'd210};
ram[50442] = {9'd13,10'd213};
ram[50443] = {9'd16,10'd216};
ram[50444] = {9'd19,10'd219};
ram[50445] = {9'd22,10'd223};
ram[50446] = {9'd25,10'd226};
ram[50447] = {9'd29,10'd229};
ram[50448] = {9'd32,10'd232};
ram[50449] = {9'd35,10'd235};
ram[50450] = {9'd38,10'd238};
ram[50451] = {9'd41,10'd241};
ram[50452] = {9'd44,10'd245};
ram[50453] = {9'd47,10'd248};
ram[50454] = {9'd51,10'd251};
ram[50455] = {9'd54,10'd254};
ram[50456] = {9'd57,10'd257};
ram[50457] = {9'd60,10'd260};
ram[50458] = {9'd63,10'd263};
ram[50459] = {9'd66,10'd267};
ram[50460] = {9'd69,10'd270};
ram[50461] = {9'd73,10'd273};
ram[50462] = {9'd76,10'd276};
ram[50463] = {9'd79,10'd279};
ram[50464] = {9'd82,10'd282};
ram[50465] = {9'd85,10'd285};
ram[50466] = {9'd88,10'd289};
ram[50467] = {9'd91,10'd292};
ram[50468] = {9'd95,10'd295};
ram[50469] = {9'd98,10'd298};
ram[50470] = {-9'd99,10'd301};
ram[50471] = {-9'd96,10'd304};
ram[50472] = {-9'd93,10'd307};
ram[50473] = {-9'd90,10'd311};
ram[50474] = {-9'd87,10'd314};
ram[50475] = {-9'd84,10'd317};
ram[50476] = {-9'd81,10'd320};
ram[50477] = {-9'd77,10'd323};
ram[50478] = {-9'd74,10'd326};
ram[50479] = {-9'd71,10'd329};
ram[50480] = {-9'd68,10'd333};
ram[50481] = {-9'd65,10'd336};
ram[50482] = {-9'd62,10'd339};
ram[50483] = {-9'd59,10'd342};
ram[50484] = {-9'd55,10'd345};
ram[50485] = {-9'd52,10'd348};
ram[50486] = {-9'd49,10'd351};
ram[50487] = {-9'd46,10'd354};
ram[50488] = {-9'd43,10'd358};
ram[50489] = {-9'd40,10'd361};
ram[50490] = {-9'd37,10'd364};
ram[50491] = {-9'd33,10'd367};
ram[50492] = {-9'd30,10'd370};
ram[50493] = {-9'd27,10'd373};
ram[50494] = {-9'd24,10'd376};
ram[50495] = {-9'd21,10'd380};
ram[50496] = {-9'd18,10'd383};
ram[50497] = {-9'd15,10'd386};
ram[50498] = {-9'd11,10'd389};
ram[50499] = {-9'd8,10'd392};
ram[50500] = {-9'd5,10'd395};
ram[50501] = {-9'd2,10'd398};
ram[50502] = {9'd1,-10'd399};
ram[50503] = {9'd4,-10'd396};
ram[50504] = {9'd7,-10'd393};
ram[50505] = {9'd10,-10'd390};
ram[50506] = {9'd14,-10'd387};
ram[50507] = {9'd17,-10'd384};
ram[50508] = {9'd20,-10'd381};
ram[50509] = {9'd23,-10'd377};
ram[50510] = {9'd26,-10'd374};
ram[50511] = {9'd29,-10'd371};
ram[50512] = {9'd32,-10'd368};
ram[50513] = {9'd36,-10'd365};
ram[50514] = {9'd39,-10'd362};
ram[50515] = {9'd42,-10'd359};
ram[50516] = {9'd45,-10'd355};
ram[50517] = {9'd48,-10'd352};
ram[50518] = {9'd51,-10'd349};
ram[50519] = {9'd54,-10'd346};
ram[50520] = {9'd58,-10'd343};
ram[50521] = {9'd61,-10'd340};
ram[50522] = {9'd64,-10'd337};
ram[50523] = {9'd67,-10'd334};
ram[50524] = {9'd70,-10'd330};
ram[50525] = {9'd73,-10'd327};
ram[50526] = {9'd76,-10'd324};
ram[50527] = {9'd80,-10'd321};
ram[50528] = {9'd83,-10'd318};
ram[50529] = {9'd86,-10'd315};
ram[50530] = {9'd89,-10'd312};
ram[50531] = {9'd92,-10'd308};
ram[50532] = {9'd95,-10'd305};
ram[50533] = {9'd98,-10'd302};
ram[50534] = {-9'd99,-10'd299};
ram[50535] = {-9'd96,-10'd296};
ram[50536] = {-9'd92,-10'd293};
ram[50537] = {-9'd89,-10'd290};
ram[50538] = {-9'd86,-10'd286};
ram[50539] = {-9'd83,-10'd283};
ram[50540] = {-9'd80,-10'd280};
ram[50541] = {-9'd77,-10'd277};
ram[50542] = {-9'd74,-10'd274};
ram[50543] = {-9'd70,-10'd271};
ram[50544] = {-9'd67,-10'd268};
ram[50545] = {-9'd64,-10'd264};
ram[50546] = {-9'd61,-10'd261};
ram[50547] = {-9'd58,-10'd258};
ram[50548] = {-9'd55,-10'd255};
ram[50549] = {-9'd52,-10'd252};
ram[50550] = {-9'd48,-10'd249};
ram[50551] = {-9'd45,-10'd246};
ram[50552] = {-9'd42,-10'd242};
ram[50553] = {-9'd39,-10'd239};
ram[50554] = {-9'd36,-10'd236};
ram[50555] = {-9'd33,-10'd233};
ram[50556] = {-9'd30,-10'd230};
ram[50557] = {-9'd26,-10'd227};
ram[50558] = {-9'd23,-10'd224};
ram[50559] = {-9'd20,-10'd220};
ram[50560] = {-9'd20,-10'd220};
ram[50561] = {-9'd17,-10'd217};
ram[50562] = {-9'd14,-10'd214};
ram[50563] = {-9'd11,-10'd211};
ram[50564] = {-9'd8,-10'd208};
ram[50565] = {-9'd4,-10'd205};
ram[50566] = {-9'd1,-10'd202};
ram[50567] = {9'd2,-10'd198};
ram[50568] = {9'd5,-10'd195};
ram[50569] = {9'd8,-10'd192};
ram[50570] = {9'd11,-10'd189};
ram[50571] = {9'd14,-10'd186};
ram[50572] = {9'd18,-10'd183};
ram[50573] = {9'd21,-10'd180};
ram[50574] = {9'd24,-10'd176};
ram[50575] = {9'd27,-10'd173};
ram[50576] = {9'd30,-10'd170};
ram[50577] = {9'd33,-10'd167};
ram[50578] = {9'd36,-10'd164};
ram[50579] = {9'd40,-10'd161};
ram[50580] = {9'd43,-10'd158};
ram[50581] = {9'd46,-10'd154};
ram[50582] = {9'd49,-10'd151};
ram[50583] = {9'd52,-10'd148};
ram[50584] = {9'd55,-10'd145};
ram[50585] = {9'd58,-10'd142};
ram[50586] = {9'd62,-10'd139};
ram[50587] = {9'd65,-10'd136};
ram[50588] = {9'd68,-10'd132};
ram[50589] = {9'd71,-10'd129};
ram[50590] = {9'd74,-10'd126};
ram[50591] = {9'd77,-10'd123};
ram[50592] = {9'd80,-10'd120};
ram[50593] = {9'd84,-10'd117};
ram[50594] = {9'd87,-10'd114};
ram[50595] = {9'd90,-10'd110};
ram[50596] = {9'd93,-10'd107};
ram[50597] = {9'd96,-10'd104};
ram[50598] = {9'd99,-10'd101};
ram[50599] = {-9'd98,-10'd98};
ram[50600] = {-9'd95,-10'd95};
ram[50601] = {-9'd92,-10'd92};
ram[50602] = {-9'd88,-10'd88};
ram[50603] = {-9'd85,-10'd85};
ram[50604] = {-9'd82,-10'd82};
ram[50605] = {-9'd79,-10'd79};
ram[50606] = {-9'd76,-10'd76};
ram[50607] = {-9'd73,-10'd73};
ram[50608] = {-9'd70,-10'd70};
ram[50609] = {-9'd66,-10'd66};
ram[50610] = {-9'd63,-10'd63};
ram[50611] = {-9'd60,-10'd60};
ram[50612] = {-9'd57,-10'd57};
ram[50613] = {-9'd54,-10'd54};
ram[50614] = {-9'd51,-10'd51};
ram[50615] = {-9'd48,-10'd48};
ram[50616] = {-9'd44,-10'd44};
ram[50617] = {-9'd41,-10'd41};
ram[50618] = {-9'd38,-10'd38};
ram[50619] = {-9'd35,-10'd35};
ram[50620] = {-9'd32,-10'd32};
ram[50621] = {-9'd29,-10'd29};
ram[50622] = {-9'd26,-10'd26};
ram[50623] = {-9'd22,-10'd22};
ram[50624] = {-9'd19,-10'd19};
ram[50625] = {-9'd16,-10'd16};
ram[50626] = {-9'd13,-10'd13};
ram[50627] = {-9'd10,-10'd10};
ram[50628] = {-9'd7,-10'd7};
ram[50629] = {-9'd4,-10'd4};
ram[50630] = {9'd0,10'd0};
ram[50631] = {9'd3,10'd3};
ram[50632] = {9'd6,10'd6};
ram[50633] = {9'd9,10'd9};
ram[50634] = {9'd12,10'd12};
ram[50635] = {9'd15,10'd15};
ram[50636] = {9'd18,10'd18};
ram[50637] = {9'd21,10'd21};
ram[50638] = {9'd25,10'd25};
ram[50639] = {9'd28,10'd28};
ram[50640] = {9'd31,10'd31};
ram[50641] = {9'd34,10'd34};
ram[50642] = {9'd37,10'd37};
ram[50643] = {9'd40,10'd40};
ram[50644] = {9'd43,10'd43};
ram[50645] = {9'd47,10'd47};
ram[50646] = {9'd50,10'd50};
ram[50647] = {9'd53,10'd53};
ram[50648] = {9'd56,10'd56};
ram[50649] = {9'd59,10'd59};
ram[50650] = {9'd62,10'd62};
ram[50651] = {9'd65,10'd65};
ram[50652] = {9'd69,10'd69};
ram[50653] = {9'd72,10'd72};
ram[50654] = {9'd75,10'd75};
ram[50655] = {9'd78,10'd78};
ram[50656] = {9'd81,10'd81};
ram[50657] = {9'd84,10'd84};
ram[50658] = {9'd87,10'd87};
ram[50659] = {9'd91,10'd91};
ram[50660] = {9'd94,10'd94};
ram[50661] = {9'd97,10'd97};
ram[50662] = {-9'd100,10'd100};
ram[50663] = {-9'd97,10'd103};
ram[50664] = {-9'd94,10'd106};
ram[50665] = {-9'd91,10'd109};
ram[50666] = {-9'd88,10'd113};
ram[50667] = {-9'd85,10'd116};
ram[50668] = {-9'd81,10'd119};
ram[50669] = {-9'd78,10'd122};
ram[50670] = {-9'd75,10'd125};
ram[50671] = {-9'd72,10'd128};
ram[50672] = {-9'd69,10'd131};
ram[50673] = {-9'd66,10'd135};
ram[50674] = {-9'd63,10'd138};
ram[50675] = {-9'd59,10'd141};
ram[50676] = {-9'd56,10'd144};
ram[50677] = {-9'd53,10'd147};
ram[50678] = {-9'd50,10'd150};
ram[50679] = {-9'd47,10'd153};
ram[50680] = {-9'd44,10'd157};
ram[50681] = {-9'd41,10'd160};
ram[50682] = {-9'd37,10'd163};
ram[50683] = {-9'd34,10'd166};
ram[50684] = {-9'd31,10'd169};
ram[50685] = {-9'd28,10'd172};
ram[50686] = {-9'd25,10'd175};
ram[50687] = {-9'd22,10'd179};
ram[50688] = {-9'd22,10'd179};
ram[50689] = {-9'd19,10'd182};
ram[50690] = {-9'd15,10'd185};
ram[50691] = {-9'd12,10'd188};
ram[50692] = {-9'd9,10'd191};
ram[50693] = {-9'd6,10'd194};
ram[50694] = {-9'd3,10'd197};
ram[50695] = {9'd0,10'd201};
ram[50696] = {9'd3,10'd204};
ram[50697] = {9'd7,10'd207};
ram[50698] = {9'd10,10'd210};
ram[50699] = {9'd13,10'd213};
ram[50700] = {9'd16,10'd216};
ram[50701] = {9'd19,10'd219};
ram[50702] = {9'd22,10'd223};
ram[50703] = {9'd25,10'd226};
ram[50704] = {9'd29,10'd229};
ram[50705] = {9'd32,10'd232};
ram[50706] = {9'd35,10'd235};
ram[50707] = {9'd38,10'd238};
ram[50708] = {9'd41,10'd241};
ram[50709] = {9'd44,10'd245};
ram[50710] = {9'd47,10'd248};
ram[50711] = {9'd51,10'd251};
ram[50712] = {9'd54,10'd254};
ram[50713] = {9'd57,10'd257};
ram[50714] = {9'd60,10'd260};
ram[50715] = {9'd63,10'd263};
ram[50716] = {9'd66,10'd267};
ram[50717] = {9'd69,10'd270};
ram[50718] = {9'd73,10'd273};
ram[50719] = {9'd76,10'd276};
ram[50720] = {9'd79,10'd279};
ram[50721] = {9'd82,10'd282};
ram[50722] = {9'd85,10'd285};
ram[50723] = {9'd88,10'd289};
ram[50724] = {9'd91,10'd292};
ram[50725] = {9'd95,10'd295};
ram[50726] = {9'd98,10'd298};
ram[50727] = {-9'd99,10'd301};
ram[50728] = {-9'd96,10'd304};
ram[50729] = {-9'd93,10'd307};
ram[50730] = {-9'd90,10'd311};
ram[50731] = {-9'd87,10'd314};
ram[50732] = {-9'd84,10'd317};
ram[50733] = {-9'd81,10'd320};
ram[50734] = {-9'd77,10'd323};
ram[50735] = {-9'd74,10'd326};
ram[50736] = {-9'd71,10'd329};
ram[50737] = {-9'd68,10'd333};
ram[50738] = {-9'd65,10'd336};
ram[50739] = {-9'd62,10'd339};
ram[50740] = {-9'd59,10'd342};
ram[50741] = {-9'd55,10'd345};
ram[50742] = {-9'd52,10'd348};
ram[50743] = {-9'd49,10'd351};
ram[50744] = {-9'd46,10'd354};
ram[50745] = {-9'd43,10'd358};
ram[50746] = {-9'd40,10'd361};
ram[50747] = {-9'd37,10'd364};
ram[50748] = {-9'd33,10'd367};
ram[50749] = {-9'd30,10'd370};
ram[50750] = {-9'd27,10'd373};
ram[50751] = {-9'd24,10'd376};
ram[50752] = {-9'd21,10'd380};
ram[50753] = {-9'd18,10'd383};
ram[50754] = {-9'd15,10'd386};
ram[50755] = {-9'd11,10'd389};
ram[50756] = {-9'd8,10'd392};
ram[50757] = {-9'd5,10'd395};
ram[50758] = {-9'd2,10'd398};
ram[50759] = {9'd1,-10'd399};
ram[50760] = {9'd4,-10'd396};
ram[50761] = {9'd7,-10'd393};
ram[50762] = {9'd10,-10'd390};
ram[50763] = {9'd14,-10'd387};
ram[50764] = {9'd17,-10'd384};
ram[50765] = {9'd20,-10'd381};
ram[50766] = {9'd23,-10'd377};
ram[50767] = {9'd26,-10'd374};
ram[50768] = {9'd29,-10'd371};
ram[50769] = {9'd32,-10'd368};
ram[50770] = {9'd36,-10'd365};
ram[50771] = {9'd39,-10'd362};
ram[50772] = {9'd42,-10'd359};
ram[50773] = {9'd45,-10'd355};
ram[50774] = {9'd48,-10'd352};
ram[50775] = {9'd51,-10'd349};
ram[50776] = {9'd54,-10'd346};
ram[50777] = {9'd58,-10'd343};
ram[50778] = {9'd61,-10'd340};
ram[50779] = {9'd64,-10'd337};
ram[50780] = {9'd67,-10'd334};
ram[50781] = {9'd70,-10'd330};
ram[50782] = {9'd73,-10'd327};
ram[50783] = {9'd76,-10'd324};
ram[50784] = {9'd80,-10'd321};
ram[50785] = {9'd83,-10'd318};
ram[50786] = {9'd86,-10'd315};
ram[50787] = {9'd89,-10'd312};
ram[50788] = {9'd92,-10'd308};
ram[50789] = {9'd95,-10'd305};
ram[50790] = {9'd98,-10'd302};
ram[50791] = {-9'd99,-10'd299};
ram[50792] = {-9'd96,-10'd296};
ram[50793] = {-9'd92,-10'd293};
ram[50794] = {-9'd89,-10'd290};
ram[50795] = {-9'd86,-10'd286};
ram[50796] = {-9'd83,-10'd283};
ram[50797] = {-9'd80,-10'd280};
ram[50798] = {-9'd77,-10'd277};
ram[50799] = {-9'd74,-10'd274};
ram[50800] = {-9'd70,-10'd271};
ram[50801] = {-9'd67,-10'd268};
ram[50802] = {-9'd64,-10'd264};
ram[50803] = {-9'd61,-10'd261};
ram[50804] = {-9'd58,-10'd258};
ram[50805] = {-9'd55,-10'd255};
ram[50806] = {-9'd52,-10'd252};
ram[50807] = {-9'd48,-10'd249};
ram[50808] = {-9'd45,-10'd246};
ram[50809] = {-9'd42,-10'd242};
ram[50810] = {-9'd39,-10'd239};
ram[50811] = {-9'd36,-10'd236};
ram[50812] = {-9'd33,-10'd233};
ram[50813] = {-9'd30,-10'd230};
ram[50814] = {-9'd26,-10'd227};
ram[50815] = {-9'd23,-10'd224};
ram[50816] = {-9'd23,-10'd224};
ram[50817] = {-9'd20,-10'd220};
ram[50818] = {-9'd17,-10'd217};
ram[50819] = {-9'd14,-10'd214};
ram[50820] = {-9'd11,-10'd211};
ram[50821] = {-9'd8,-10'd208};
ram[50822] = {-9'd4,-10'd205};
ram[50823] = {-9'd1,-10'd202};
ram[50824] = {9'd2,-10'd198};
ram[50825] = {9'd5,-10'd195};
ram[50826] = {9'd8,-10'd192};
ram[50827] = {9'd11,-10'd189};
ram[50828] = {9'd14,-10'd186};
ram[50829] = {9'd18,-10'd183};
ram[50830] = {9'd21,-10'd180};
ram[50831] = {9'd24,-10'd176};
ram[50832] = {9'd27,-10'd173};
ram[50833] = {9'd30,-10'd170};
ram[50834] = {9'd33,-10'd167};
ram[50835] = {9'd36,-10'd164};
ram[50836] = {9'd40,-10'd161};
ram[50837] = {9'd43,-10'd158};
ram[50838] = {9'd46,-10'd154};
ram[50839] = {9'd49,-10'd151};
ram[50840] = {9'd52,-10'd148};
ram[50841] = {9'd55,-10'd145};
ram[50842] = {9'd58,-10'd142};
ram[50843] = {9'd62,-10'd139};
ram[50844] = {9'd65,-10'd136};
ram[50845] = {9'd68,-10'd132};
ram[50846] = {9'd71,-10'd129};
ram[50847] = {9'd74,-10'd126};
ram[50848] = {9'd77,-10'd123};
ram[50849] = {9'd80,-10'd120};
ram[50850] = {9'd84,-10'd117};
ram[50851] = {9'd87,-10'd114};
ram[50852] = {9'd90,-10'd110};
ram[50853] = {9'd93,-10'd107};
ram[50854] = {9'd96,-10'd104};
ram[50855] = {9'd99,-10'd101};
ram[50856] = {-9'd98,-10'd98};
ram[50857] = {-9'd95,-10'd95};
ram[50858] = {-9'd92,-10'd92};
ram[50859] = {-9'd88,-10'd88};
ram[50860] = {-9'd85,-10'd85};
ram[50861] = {-9'd82,-10'd82};
ram[50862] = {-9'd79,-10'd79};
ram[50863] = {-9'd76,-10'd76};
ram[50864] = {-9'd73,-10'd73};
ram[50865] = {-9'd70,-10'd70};
ram[50866] = {-9'd66,-10'd66};
ram[50867] = {-9'd63,-10'd63};
ram[50868] = {-9'd60,-10'd60};
ram[50869] = {-9'd57,-10'd57};
ram[50870] = {-9'd54,-10'd54};
ram[50871] = {-9'd51,-10'd51};
ram[50872] = {-9'd48,-10'd48};
ram[50873] = {-9'd44,-10'd44};
ram[50874] = {-9'd41,-10'd41};
ram[50875] = {-9'd38,-10'd38};
ram[50876] = {-9'd35,-10'd35};
ram[50877] = {-9'd32,-10'd32};
ram[50878] = {-9'd29,-10'd29};
ram[50879] = {-9'd26,-10'd26};
ram[50880] = {-9'd22,-10'd22};
ram[50881] = {-9'd19,-10'd19};
ram[50882] = {-9'd16,-10'd16};
ram[50883] = {-9'd13,-10'd13};
ram[50884] = {-9'd10,-10'd10};
ram[50885] = {-9'd7,-10'd7};
ram[50886] = {-9'd4,-10'd4};
ram[50887] = {9'd0,10'd0};
ram[50888] = {9'd3,10'd3};
ram[50889] = {9'd6,10'd6};
ram[50890] = {9'd9,10'd9};
ram[50891] = {9'd12,10'd12};
ram[50892] = {9'd15,10'd15};
ram[50893] = {9'd18,10'd18};
ram[50894] = {9'd21,10'd21};
ram[50895] = {9'd25,10'd25};
ram[50896] = {9'd28,10'd28};
ram[50897] = {9'd31,10'd31};
ram[50898] = {9'd34,10'd34};
ram[50899] = {9'd37,10'd37};
ram[50900] = {9'd40,10'd40};
ram[50901] = {9'd43,10'd43};
ram[50902] = {9'd47,10'd47};
ram[50903] = {9'd50,10'd50};
ram[50904] = {9'd53,10'd53};
ram[50905] = {9'd56,10'd56};
ram[50906] = {9'd59,10'd59};
ram[50907] = {9'd62,10'd62};
ram[50908] = {9'd65,10'd65};
ram[50909] = {9'd69,10'd69};
ram[50910] = {9'd72,10'd72};
ram[50911] = {9'd75,10'd75};
ram[50912] = {9'd78,10'd78};
ram[50913] = {9'd81,10'd81};
ram[50914] = {9'd84,10'd84};
ram[50915] = {9'd87,10'd87};
ram[50916] = {9'd91,10'd91};
ram[50917] = {9'd94,10'd94};
ram[50918] = {9'd97,10'd97};
ram[50919] = {-9'd100,10'd100};
ram[50920] = {-9'd97,10'd103};
ram[50921] = {-9'd94,10'd106};
ram[50922] = {-9'd91,10'd109};
ram[50923] = {-9'd88,10'd113};
ram[50924] = {-9'd85,10'd116};
ram[50925] = {-9'd81,10'd119};
ram[50926] = {-9'd78,10'd122};
ram[50927] = {-9'd75,10'd125};
ram[50928] = {-9'd72,10'd128};
ram[50929] = {-9'd69,10'd131};
ram[50930] = {-9'd66,10'd135};
ram[50931] = {-9'd63,10'd138};
ram[50932] = {-9'd59,10'd141};
ram[50933] = {-9'd56,10'd144};
ram[50934] = {-9'd53,10'd147};
ram[50935] = {-9'd50,10'd150};
ram[50936] = {-9'd47,10'd153};
ram[50937] = {-9'd44,10'd157};
ram[50938] = {-9'd41,10'd160};
ram[50939] = {-9'd37,10'd163};
ram[50940] = {-9'd34,10'd166};
ram[50941] = {-9'd31,10'd169};
ram[50942] = {-9'd28,10'd172};
ram[50943] = {-9'd25,10'd175};
ram[50944] = {-9'd25,10'd175};
ram[50945] = {-9'd22,10'd179};
ram[50946] = {-9'd19,10'd182};
ram[50947] = {-9'd15,10'd185};
ram[50948] = {-9'd12,10'd188};
ram[50949] = {-9'd9,10'd191};
ram[50950] = {-9'd6,10'd194};
ram[50951] = {-9'd3,10'd197};
ram[50952] = {9'd0,10'd201};
ram[50953] = {9'd3,10'd204};
ram[50954] = {9'd7,10'd207};
ram[50955] = {9'd10,10'd210};
ram[50956] = {9'd13,10'd213};
ram[50957] = {9'd16,10'd216};
ram[50958] = {9'd19,10'd219};
ram[50959] = {9'd22,10'd223};
ram[50960] = {9'd25,10'd226};
ram[50961] = {9'd29,10'd229};
ram[50962] = {9'd32,10'd232};
ram[50963] = {9'd35,10'd235};
ram[50964] = {9'd38,10'd238};
ram[50965] = {9'd41,10'd241};
ram[50966] = {9'd44,10'd245};
ram[50967] = {9'd47,10'd248};
ram[50968] = {9'd51,10'd251};
ram[50969] = {9'd54,10'd254};
ram[50970] = {9'd57,10'd257};
ram[50971] = {9'd60,10'd260};
ram[50972] = {9'd63,10'd263};
ram[50973] = {9'd66,10'd267};
ram[50974] = {9'd69,10'd270};
ram[50975] = {9'd73,10'd273};
ram[50976] = {9'd76,10'd276};
ram[50977] = {9'd79,10'd279};
ram[50978] = {9'd82,10'd282};
ram[50979] = {9'd85,10'd285};
ram[50980] = {9'd88,10'd289};
ram[50981] = {9'd91,10'd292};
ram[50982] = {9'd95,10'd295};
ram[50983] = {9'd98,10'd298};
ram[50984] = {-9'd99,10'd301};
ram[50985] = {-9'd96,10'd304};
ram[50986] = {-9'd93,10'd307};
ram[50987] = {-9'd90,10'd311};
ram[50988] = {-9'd87,10'd314};
ram[50989] = {-9'd84,10'd317};
ram[50990] = {-9'd81,10'd320};
ram[50991] = {-9'd77,10'd323};
ram[50992] = {-9'd74,10'd326};
ram[50993] = {-9'd71,10'd329};
ram[50994] = {-9'd68,10'd333};
ram[50995] = {-9'd65,10'd336};
ram[50996] = {-9'd62,10'd339};
ram[50997] = {-9'd59,10'd342};
ram[50998] = {-9'd55,10'd345};
ram[50999] = {-9'd52,10'd348};
ram[51000] = {-9'd49,10'd351};
ram[51001] = {-9'd46,10'd354};
ram[51002] = {-9'd43,10'd358};
ram[51003] = {-9'd40,10'd361};
ram[51004] = {-9'd37,10'd364};
ram[51005] = {-9'd33,10'd367};
ram[51006] = {-9'd30,10'd370};
ram[51007] = {-9'd27,10'd373};
ram[51008] = {-9'd24,10'd376};
ram[51009] = {-9'd21,10'd380};
ram[51010] = {-9'd18,10'd383};
ram[51011] = {-9'd15,10'd386};
ram[51012] = {-9'd11,10'd389};
ram[51013] = {-9'd8,10'd392};
ram[51014] = {-9'd5,10'd395};
ram[51015] = {-9'd2,10'd398};
ram[51016] = {9'd1,-10'd399};
ram[51017] = {9'd4,-10'd396};
ram[51018] = {9'd7,-10'd393};
ram[51019] = {9'd10,-10'd390};
ram[51020] = {9'd14,-10'd387};
ram[51021] = {9'd17,-10'd384};
ram[51022] = {9'd20,-10'd381};
ram[51023] = {9'd23,-10'd377};
ram[51024] = {9'd26,-10'd374};
ram[51025] = {9'd29,-10'd371};
ram[51026] = {9'd32,-10'd368};
ram[51027] = {9'd36,-10'd365};
ram[51028] = {9'd39,-10'd362};
ram[51029] = {9'd42,-10'd359};
ram[51030] = {9'd45,-10'd355};
ram[51031] = {9'd48,-10'd352};
ram[51032] = {9'd51,-10'd349};
ram[51033] = {9'd54,-10'd346};
ram[51034] = {9'd58,-10'd343};
ram[51035] = {9'd61,-10'd340};
ram[51036] = {9'd64,-10'd337};
ram[51037] = {9'd67,-10'd334};
ram[51038] = {9'd70,-10'd330};
ram[51039] = {9'd73,-10'd327};
ram[51040] = {9'd76,-10'd324};
ram[51041] = {9'd80,-10'd321};
ram[51042] = {9'd83,-10'd318};
ram[51043] = {9'd86,-10'd315};
ram[51044] = {9'd89,-10'd312};
ram[51045] = {9'd92,-10'd308};
ram[51046] = {9'd95,-10'd305};
ram[51047] = {9'd98,-10'd302};
ram[51048] = {-9'd99,-10'd299};
ram[51049] = {-9'd96,-10'd296};
ram[51050] = {-9'd92,-10'd293};
ram[51051] = {-9'd89,-10'd290};
ram[51052] = {-9'd86,-10'd286};
ram[51053] = {-9'd83,-10'd283};
ram[51054] = {-9'd80,-10'd280};
ram[51055] = {-9'd77,-10'd277};
ram[51056] = {-9'd74,-10'd274};
ram[51057] = {-9'd70,-10'd271};
ram[51058] = {-9'd67,-10'd268};
ram[51059] = {-9'd64,-10'd264};
ram[51060] = {-9'd61,-10'd261};
ram[51061] = {-9'd58,-10'd258};
ram[51062] = {-9'd55,-10'd255};
ram[51063] = {-9'd52,-10'd252};
ram[51064] = {-9'd48,-10'd249};
ram[51065] = {-9'd45,-10'd246};
ram[51066] = {-9'd42,-10'd242};
ram[51067] = {-9'd39,-10'd239};
ram[51068] = {-9'd36,-10'd236};
ram[51069] = {-9'd33,-10'd233};
ram[51070] = {-9'd30,-10'd230};
ram[51071] = {-9'd26,-10'd227};
ram[51072] = {-9'd26,-10'd227};
ram[51073] = {-9'd23,-10'd224};
ram[51074] = {-9'd20,-10'd220};
ram[51075] = {-9'd17,-10'd217};
ram[51076] = {-9'd14,-10'd214};
ram[51077] = {-9'd11,-10'd211};
ram[51078] = {-9'd8,-10'd208};
ram[51079] = {-9'd4,-10'd205};
ram[51080] = {-9'd1,-10'd202};
ram[51081] = {9'd2,-10'd198};
ram[51082] = {9'd5,-10'd195};
ram[51083] = {9'd8,-10'd192};
ram[51084] = {9'd11,-10'd189};
ram[51085] = {9'd14,-10'd186};
ram[51086] = {9'd18,-10'd183};
ram[51087] = {9'd21,-10'd180};
ram[51088] = {9'd24,-10'd176};
ram[51089] = {9'd27,-10'd173};
ram[51090] = {9'd30,-10'd170};
ram[51091] = {9'd33,-10'd167};
ram[51092] = {9'd36,-10'd164};
ram[51093] = {9'd40,-10'd161};
ram[51094] = {9'd43,-10'd158};
ram[51095] = {9'd46,-10'd154};
ram[51096] = {9'd49,-10'd151};
ram[51097] = {9'd52,-10'd148};
ram[51098] = {9'd55,-10'd145};
ram[51099] = {9'd58,-10'd142};
ram[51100] = {9'd62,-10'd139};
ram[51101] = {9'd65,-10'd136};
ram[51102] = {9'd68,-10'd132};
ram[51103] = {9'd71,-10'd129};
ram[51104] = {9'd74,-10'd126};
ram[51105] = {9'd77,-10'd123};
ram[51106] = {9'd80,-10'd120};
ram[51107] = {9'd84,-10'd117};
ram[51108] = {9'd87,-10'd114};
ram[51109] = {9'd90,-10'd110};
ram[51110] = {9'd93,-10'd107};
ram[51111] = {9'd96,-10'd104};
ram[51112] = {9'd99,-10'd101};
ram[51113] = {-9'd98,-10'd98};
ram[51114] = {-9'd95,-10'd95};
ram[51115] = {-9'd92,-10'd92};
ram[51116] = {-9'd88,-10'd88};
ram[51117] = {-9'd85,-10'd85};
ram[51118] = {-9'd82,-10'd82};
ram[51119] = {-9'd79,-10'd79};
ram[51120] = {-9'd76,-10'd76};
ram[51121] = {-9'd73,-10'd73};
ram[51122] = {-9'd70,-10'd70};
ram[51123] = {-9'd66,-10'd66};
ram[51124] = {-9'd63,-10'd63};
ram[51125] = {-9'd60,-10'd60};
ram[51126] = {-9'd57,-10'd57};
ram[51127] = {-9'd54,-10'd54};
ram[51128] = {-9'd51,-10'd51};
ram[51129] = {-9'd48,-10'd48};
ram[51130] = {-9'd44,-10'd44};
ram[51131] = {-9'd41,-10'd41};
ram[51132] = {-9'd38,-10'd38};
ram[51133] = {-9'd35,-10'd35};
ram[51134] = {-9'd32,-10'd32};
ram[51135] = {-9'd29,-10'd29};
ram[51136] = {-9'd26,-10'd26};
ram[51137] = {-9'd22,-10'd22};
ram[51138] = {-9'd19,-10'd19};
ram[51139] = {-9'd16,-10'd16};
ram[51140] = {-9'd13,-10'd13};
ram[51141] = {-9'd10,-10'd10};
ram[51142] = {-9'd7,-10'd7};
ram[51143] = {-9'd4,-10'd4};
ram[51144] = {9'd0,10'd0};
ram[51145] = {9'd3,10'd3};
ram[51146] = {9'd6,10'd6};
ram[51147] = {9'd9,10'd9};
ram[51148] = {9'd12,10'd12};
ram[51149] = {9'd15,10'd15};
ram[51150] = {9'd18,10'd18};
ram[51151] = {9'd21,10'd21};
ram[51152] = {9'd25,10'd25};
ram[51153] = {9'd28,10'd28};
ram[51154] = {9'd31,10'd31};
ram[51155] = {9'd34,10'd34};
ram[51156] = {9'd37,10'd37};
ram[51157] = {9'd40,10'd40};
ram[51158] = {9'd43,10'd43};
ram[51159] = {9'd47,10'd47};
ram[51160] = {9'd50,10'd50};
ram[51161] = {9'd53,10'd53};
ram[51162] = {9'd56,10'd56};
ram[51163] = {9'd59,10'd59};
ram[51164] = {9'd62,10'd62};
ram[51165] = {9'd65,10'd65};
ram[51166] = {9'd69,10'd69};
ram[51167] = {9'd72,10'd72};
ram[51168] = {9'd75,10'd75};
ram[51169] = {9'd78,10'd78};
ram[51170] = {9'd81,10'd81};
ram[51171] = {9'd84,10'd84};
ram[51172] = {9'd87,10'd87};
ram[51173] = {9'd91,10'd91};
ram[51174] = {9'd94,10'd94};
ram[51175] = {9'd97,10'd97};
ram[51176] = {-9'd100,10'd100};
ram[51177] = {-9'd97,10'd103};
ram[51178] = {-9'd94,10'd106};
ram[51179] = {-9'd91,10'd109};
ram[51180] = {-9'd88,10'd113};
ram[51181] = {-9'd85,10'd116};
ram[51182] = {-9'd81,10'd119};
ram[51183] = {-9'd78,10'd122};
ram[51184] = {-9'd75,10'd125};
ram[51185] = {-9'd72,10'd128};
ram[51186] = {-9'd69,10'd131};
ram[51187] = {-9'd66,10'd135};
ram[51188] = {-9'd63,10'd138};
ram[51189] = {-9'd59,10'd141};
ram[51190] = {-9'd56,10'd144};
ram[51191] = {-9'd53,10'd147};
ram[51192] = {-9'd50,10'd150};
ram[51193] = {-9'd47,10'd153};
ram[51194] = {-9'd44,10'd157};
ram[51195] = {-9'd41,10'd160};
ram[51196] = {-9'd37,10'd163};
ram[51197] = {-9'd34,10'd166};
ram[51198] = {-9'd31,10'd169};
ram[51199] = {-9'd28,10'd172};
ram[51200] = {-9'd28,10'd172};
ram[51201] = {-9'd25,10'd175};
ram[51202] = {-9'd22,10'd179};
ram[51203] = {-9'd19,10'd182};
ram[51204] = {-9'd15,10'd185};
ram[51205] = {-9'd12,10'd188};
ram[51206] = {-9'd9,10'd191};
ram[51207] = {-9'd6,10'd194};
ram[51208] = {-9'd3,10'd197};
ram[51209] = {9'd0,10'd201};
ram[51210] = {9'd3,10'd204};
ram[51211] = {9'd7,10'd207};
ram[51212] = {9'd10,10'd210};
ram[51213] = {9'd13,10'd213};
ram[51214] = {9'd16,10'd216};
ram[51215] = {9'd19,10'd219};
ram[51216] = {9'd22,10'd223};
ram[51217] = {9'd25,10'd226};
ram[51218] = {9'd29,10'd229};
ram[51219] = {9'd32,10'd232};
ram[51220] = {9'd35,10'd235};
ram[51221] = {9'd38,10'd238};
ram[51222] = {9'd41,10'd241};
ram[51223] = {9'd44,10'd245};
ram[51224] = {9'd47,10'd248};
ram[51225] = {9'd51,10'd251};
ram[51226] = {9'd54,10'd254};
ram[51227] = {9'd57,10'd257};
ram[51228] = {9'd60,10'd260};
ram[51229] = {9'd63,10'd263};
ram[51230] = {9'd66,10'd267};
ram[51231] = {9'd69,10'd270};
ram[51232] = {9'd73,10'd273};
ram[51233] = {9'd76,10'd276};
ram[51234] = {9'd79,10'd279};
ram[51235] = {9'd82,10'd282};
ram[51236] = {9'd85,10'd285};
ram[51237] = {9'd88,10'd289};
ram[51238] = {9'd91,10'd292};
ram[51239] = {9'd95,10'd295};
ram[51240] = {9'd98,10'd298};
ram[51241] = {-9'd99,10'd301};
ram[51242] = {-9'd96,10'd304};
ram[51243] = {-9'd93,10'd307};
ram[51244] = {-9'd90,10'd311};
ram[51245] = {-9'd87,10'd314};
ram[51246] = {-9'd84,10'd317};
ram[51247] = {-9'd81,10'd320};
ram[51248] = {-9'd77,10'd323};
ram[51249] = {-9'd74,10'd326};
ram[51250] = {-9'd71,10'd329};
ram[51251] = {-9'd68,10'd333};
ram[51252] = {-9'd65,10'd336};
ram[51253] = {-9'd62,10'd339};
ram[51254] = {-9'd59,10'd342};
ram[51255] = {-9'd55,10'd345};
ram[51256] = {-9'd52,10'd348};
ram[51257] = {-9'd49,10'd351};
ram[51258] = {-9'd46,10'd354};
ram[51259] = {-9'd43,10'd358};
ram[51260] = {-9'd40,10'd361};
ram[51261] = {-9'd37,10'd364};
ram[51262] = {-9'd33,10'd367};
ram[51263] = {-9'd30,10'd370};
ram[51264] = {-9'd27,10'd373};
ram[51265] = {-9'd24,10'd376};
ram[51266] = {-9'd21,10'd380};
ram[51267] = {-9'd18,10'd383};
ram[51268] = {-9'd15,10'd386};
ram[51269] = {-9'd11,10'd389};
ram[51270] = {-9'd8,10'd392};
ram[51271] = {-9'd5,10'd395};
ram[51272] = {-9'd2,10'd398};
ram[51273] = {9'd1,-10'd399};
ram[51274] = {9'd4,-10'd396};
ram[51275] = {9'd7,-10'd393};
ram[51276] = {9'd10,-10'd390};
ram[51277] = {9'd14,-10'd387};
ram[51278] = {9'd17,-10'd384};
ram[51279] = {9'd20,-10'd381};
ram[51280] = {9'd23,-10'd377};
ram[51281] = {9'd26,-10'd374};
ram[51282] = {9'd29,-10'd371};
ram[51283] = {9'd32,-10'd368};
ram[51284] = {9'd36,-10'd365};
ram[51285] = {9'd39,-10'd362};
ram[51286] = {9'd42,-10'd359};
ram[51287] = {9'd45,-10'd355};
ram[51288] = {9'd48,-10'd352};
ram[51289] = {9'd51,-10'd349};
ram[51290] = {9'd54,-10'd346};
ram[51291] = {9'd58,-10'd343};
ram[51292] = {9'd61,-10'd340};
ram[51293] = {9'd64,-10'd337};
ram[51294] = {9'd67,-10'd334};
ram[51295] = {9'd70,-10'd330};
ram[51296] = {9'd73,-10'd327};
ram[51297] = {9'd76,-10'd324};
ram[51298] = {9'd80,-10'd321};
ram[51299] = {9'd83,-10'd318};
ram[51300] = {9'd86,-10'd315};
ram[51301] = {9'd89,-10'd312};
ram[51302] = {9'd92,-10'd308};
ram[51303] = {9'd95,-10'd305};
ram[51304] = {9'd98,-10'd302};
ram[51305] = {-9'd99,-10'd299};
ram[51306] = {-9'd96,-10'd296};
ram[51307] = {-9'd92,-10'd293};
ram[51308] = {-9'd89,-10'd290};
ram[51309] = {-9'd86,-10'd286};
ram[51310] = {-9'd83,-10'd283};
ram[51311] = {-9'd80,-10'd280};
ram[51312] = {-9'd77,-10'd277};
ram[51313] = {-9'd74,-10'd274};
ram[51314] = {-9'd70,-10'd271};
ram[51315] = {-9'd67,-10'd268};
ram[51316] = {-9'd64,-10'd264};
ram[51317] = {-9'd61,-10'd261};
ram[51318] = {-9'd58,-10'd258};
ram[51319] = {-9'd55,-10'd255};
ram[51320] = {-9'd52,-10'd252};
ram[51321] = {-9'd48,-10'd249};
ram[51322] = {-9'd45,-10'd246};
ram[51323] = {-9'd42,-10'd242};
ram[51324] = {-9'd39,-10'd239};
ram[51325] = {-9'd36,-10'd236};
ram[51326] = {-9'd33,-10'd233};
ram[51327] = {-9'd30,-10'd230};
ram[51328] = {-9'd30,-10'd230};
ram[51329] = {-9'd26,-10'd227};
ram[51330] = {-9'd23,-10'd224};
ram[51331] = {-9'd20,-10'd220};
ram[51332] = {-9'd17,-10'd217};
ram[51333] = {-9'd14,-10'd214};
ram[51334] = {-9'd11,-10'd211};
ram[51335] = {-9'd8,-10'd208};
ram[51336] = {-9'd4,-10'd205};
ram[51337] = {-9'd1,-10'd202};
ram[51338] = {9'd2,-10'd198};
ram[51339] = {9'd5,-10'd195};
ram[51340] = {9'd8,-10'd192};
ram[51341] = {9'd11,-10'd189};
ram[51342] = {9'd14,-10'd186};
ram[51343] = {9'd18,-10'd183};
ram[51344] = {9'd21,-10'd180};
ram[51345] = {9'd24,-10'd176};
ram[51346] = {9'd27,-10'd173};
ram[51347] = {9'd30,-10'd170};
ram[51348] = {9'd33,-10'd167};
ram[51349] = {9'd36,-10'd164};
ram[51350] = {9'd40,-10'd161};
ram[51351] = {9'd43,-10'd158};
ram[51352] = {9'd46,-10'd154};
ram[51353] = {9'd49,-10'd151};
ram[51354] = {9'd52,-10'd148};
ram[51355] = {9'd55,-10'd145};
ram[51356] = {9'd58,-10'd142};
ram[51357] = {9'd62,-10'd139};
ram[51358] = {9'd65,-10'd136};
ram[51359] = {9'd68,-10'd132};
ram[51360] = {9'd71,-10'd129};
ram[51361] = {9'd74,-10'd126};
ram[51362] = {9'd77,-10'd123};
ram[51363] = {9'd80,-10'd120};
ram[51364] = {9'd84,-10'd117};
ram[51365] = {9'd87,-10'd114};
ram[51366] = {9'd90,-10'd110};
ram[51367] = {9'd93,-10'd107};
ram[51368] = {9'd96,-10'd104};
ram[51369] = {9'd99,-10'd101};
ram[51370] = {-9'd98,-10'd98};
ram[51371] = {-9'd95,-10'd95};
ram[51372] = {-9'd92,-10'd92};
ram[51373] = {-9'd88,-10'd88};
ram[51374] = {-9'd85,-10'd85};
ram[51375] = {-9'd82,-10'd82};
ram[51376] = {-9'd79,-10'd79};
ram[51377] = {-9'd76,-10'd76};
ram[51378] = {-9'd73,-10'd73};
ram[51379] = {-9'd70,-10'd70};
ram[51380] = {-9'd66,-10'd66};
ram[51381] = {-9'd63,-10'd63};
ram[51382] = {-9'd60,-10'd60};
ram[51383] = {-9'd57,-10'd57};
ram[51384] = {-9'd54,-10'd54};
ram[51385] = {-9'd51,-10'd51};
ram[51386] = {-9'd48,-10'd48};
ram[51387] = {-9'd44,-10'd44};
ram[51388] = {-9'd41,-10'd41};
ram[51389] = {-9'd38,-10'd38};
ram[51390] = {-9'd35,-10'd35};
ram[51391] = {-9'd32,-10'd32};
ram[51392] = {-9'd29,-10'd29};
ram[51393] = {-9'd26,-10'd26};
ram[51394] = {-9'd22,-10'd22};
ram[51395] = {-9'd19,-10'd19};
ram[51396] = {-9'd16,-10'd16};
ram[51397] = {-9'd13,-10'd13};
ram[51398] = {-9'd10,-10'd10};
ram[51399] = {-9'd7,-10'd7};
ram[51400] = {-9'd4,-10'd4};
ram[51401] = {9'd0,10'd0};
ram[51402] = {9'd3,10'd3};
ram[51403] = {9'd6,10'd6};
ram[51404] = {9'd9,10'd9};
ram[51405] = {9'd12,10'd12};
ram[51406] = {9'd15,10'd15};
ram[51407] = {9'd18,10'd18};
ram[51408] = {9'd21,10'd21};
ram[51409] = {9'd25,10'd25};
ram[51410] = {9'd28,10'd28};
ram[51411] = {9'd31,10'd31};
ram[51412] = {9'd34,10'd34};
ram[51413] = {9'd37,10'd37};
ram[51414] = {9'd40,10'd40};
ram[51415] = {9'd43,10'd43};
ram[51416] = {9'd47,10'd47};
ram[51417] = {9'd50,10'd50};
ram[51418] = {9'd53,10'd53};
ram[51419] = {9'd56,10'd56};
ram[51420] = {9'd59,10'd59};
ram[51421] = {9'd62,10'd62};
ram[51422] = {9'd65,10'd65};
ram[51423] = {9'd69,10'd69};
ram[51424] = {9'd72,10'd72};
ram[51425] = {9'd75,10'd75};
ram[51426] = {9'd78,10'd78};
ram[51427] = {9'd81,10'd81};
ram[51428] = {9'd84,10'd84};
ram[51429] = {9'd87,10'd87};
ram[51430] = {9'd91,10'd91};
ram[51431] = {9'd94,10'd94};
ram[51432] = {9'd97,10'd97};
ram[51433] = {-9'd100,10'd100};
ram[51434] = {-9'd97,10'd103};
ram[51435] = {-9'd94,10'd106};
ram[51436] = {-9'd91,10'd109};
ram[51437] = {-9'd88,10'd113};
ram[51438] = {-9'd85,10'd116};
ram[51439] = {-9'd81,10'd119};
ram[51440] = {-9'd78,10'd122};
ram[51441] = {-9'd75,10'd125};
ram[51442] = {-9'd72,10'd128};
ram[51443] = {-9'd69,10'd131};
ram[51444] = {-9'd66,10'd135};
ram[51445] = {-9'd63,10'd138};
ram[51446] = {-9'd59,10'd141};
ram[51447] = {-9'd56,10'd144};
ram[51448] = {-9'd53,10'd147};
ram[51449] = {-9'd50,10'd150};
ram[51450] = {-9'd47,10'd153};
ram[51451] = {-9'd44,10'd157};
ram[51452] = {-9'd41,10'd160};
ram[51453] = {-9'd37,10'd163};
ram[51454] = {-9'd34,10'd166};
ram[51455] = {-9'd31,10'd169};
ram[51456] = {-9'd31,10'd169};
ram[51457] = {-9'd28,10'd172};
ram[51458] = {-9'd25,10'd175};
ram[51459] = {-9'd22,10'd179};
ram[51460] = {-9'd19,10'd182};
ram[51461] = {-9'd15,10'd185};
ram[51462] = {-9'd12,10'd188};
ram[51463] = {-9'd9,10'd191};
ram[51464] = {-9'd6,10'd194};
ram[51465] = {-9'd3,10'd197};
ram[51466] = {9'd0,10'd201};
ram[51467] = {9'd3,10'd204};
ram[51468] = {9'd7,10'd207};
ram[51469] = {9'd10,10'd210};
ram[51470] = {9'd13,10'd213};
ram[51471] = {9'd16,10'd216};
ram[51472] = {9'd19,10'd219};
ram[51473] = {9'd22,10'd223};
ram[51474] = {9'd25,10'd226};
ram[51475] = {9'd29,10'd229};
ram[51476] = {9'd32,10'd232};
ram[51477] = {9'd35,10'd235};
ram[51478] = {9'd38,10'd238};
ram[51479] = {9'd41,10'd241};
ram[51480] = {9'd44,10'd245};
ram[51481] = {9'd47,10'd248};
ram[51482] = {9'd51,10'd251};
ram[51483] = {9'd54,10'd254};
ram[51484] = {9'd57,10'd257};
ram[51485] = {9'd60,10'd260};
ram[51486] = {9'd63,10'd263};
ram[51487] = {9'd66,10'd267};
ram[51488] = {9'd69,10'd270};
ram[51489] = {9'd73,10'd273};
ram[51490] = {9'd76,10'd276};
ram[51491] = {9'd79,10'd279};
ram[51492] = {9'd82,10'd282};
ram[51493] = {9'd85,10'd285};
ram[51494] = {9'd88,10'd289};
ram[51495] = {9'd91,10'd292};
ram[51496] = {9'd95,10'd295};
ram[51497] = {9'd98,10'd298};
ram[51498] = {-9'd99,10'd301};
ram[51499] = {-9'd96,10'd304};
ram[51500] = {-9'd93,10'd307};
ram[51501] = {-9'd90,10'd311};
ram[51502] = {-9'd87,10'd314};
ram[51503] = {-9'd84,10'd317};
ram[51504] = {-9'd81,10'd320};
ram[51505] = {-9'd77,10'd323};
ram[51506] = {-9'd74,10'd326};
ram[51507] = {-9'd71,10'd329};
ram[51508] = {-9'd68,10'd333};
ram[51509] = {-9'd65,10'd336};
ram[51510] = {-9'd62,10'd339};
ram[51511] = {-9'd59,10'd342};
ram[51512] = {-9'd55,10'd345};
ram[51513] = {-9'd52,10'd348};
ram[51514] = {-9'd49,10'd351};
ram[51515] = {-9'd46,10'd354};
ram[51516] = {-9'd43,10'd358};
ram[51517] = {-9'd40,10'd361};
ram[51518] = {-9'd37,10'd364};
ram[51519] = {-9'd33,10'd367};
ram[51520] = {-9'd30,10'd370};
ram[51521] = {-9'd27,10'd373};
ram[51522] = {-9'd24,10'd376};
ram[51523] = {-9'd21,10'd380};
ram[51524] = {-9'd18,10'd383};
ram[51525] = {-9'd15,10'd386};
ram[51526] = {-9'd11,10'd389};
ram[51527] = {-9'd8,10'd392};
ram[51528] = {-9'd5,10'd395};
ram[51529] = {-9'd2,10'd398};
ram[51530] = {9'd1,-10'd399};
ram[51531] = {9'd4,-10'd396};
ram[51532] = {9'd7,-10'd393};
ram[51533] = {9'd10,-10'd390};
ram[51534] = {9'd14,-10'd387};
ram[51535] = {9'd17,-10'd384};
ram[51536] = {9'd20,-10'd381};
ram[51537] = {9'd23,-10'd377};
ram[51538] = {9'd26,-10'd374};
ram[51539] = {9'd29,-10'd371};
ram[51540] = {9'd32,-10'd368};
ram[51541] = {9'd36,-10'd365};
ram[51542] = {9'd39,-10'd362};
ram[51543] = {9'd42,-10'd359};
ram[51544] = {9'd45,-10'd355};
ram[51545] = {9'd48,-10'd352};
ram[51546] = {9'd51,-10'd349};
ram[51547] = {9'd54,-10'd346};
ram[51548] = {9'd58,-10'd343};
ram[51549] = {9'd61,-10'd340};
ram[51550] = {9'd64,-10'd337};
ram[51551] = {9'd67,-10'd334};
ram[51552] = {9'd70,-10'd330};
ram[51553] = {9'd73,-10'd327};
ram[51554] = {9'd76,-10'd324};
ram[51555] = {9'd80,-10'd321};
ram[51556] = {9'd83,-10'd318};
ram[51557] = {9'd86,-10'd315};
ram[51558] = {9'd89,-10'd312};
ram[51559] = {9'd92,-10'd308};
ram[51560] = {9'd95,-10'd305};
ram[51561] = {9'd98,-10'd302};
ram[51562] = {-9'd99,-10'd299};
ram[51563] = {-9'd96,-10'd296};
ram[51564] = {-9'd92,-10'd293};
ram[51565] = {-9'd89,-10'd290};
ram[51566] = {-9'd86,-10'd286};
ram[51567] = {-9'd83,-10'd283};
ram[51568] = {-9'd80,-10'd280};
ram[51569] = {-9'd77,-10'd277};
ram[51570] = {-9'd74,-10'd274};
ram[51571] = {-9'd70,-10'd271};
ram[51572] = {-9'd67,-10'd268};
ram[51573] = {-9'd64,-10'd264};
ram[51574] = {-9'd61,-10'd261};
ram[51575] = {-9'd58,-10'd258};
ram[51576] = {-9'd55,-10'd255};
ram[51577] = {-9'd52,-10'd252};
ram[51578] = {-9'd48,-10'd249};
ram[51579] = {-9'd45,-10'd246};
ram[51580] = {-9'd42,-10'd242};
ram[51581] = {-9'd39,-10'd239};
ram[51582] = {-9'd36,-10'd236};
ram[51583] = {-9'd33,-10'd233};
ram[51584] = {-9'd33,-10'd233};
ram[51585] = {-9'd30,-10'd230};
ram[51586] = {-9'd26,-10'd227};
ram[51587] = {-9'd23,-10'd224};
ram[51588] = {-9'd20,-10'd220};
ram[51589] = {-9'd17,-10'd217};
ram[51590] = {-9'd14,-10'd214};
ram[51591] = {-9'd11,-10'd211};
ram[51592] = {-9'd8,-10'd208};
ram[51593] = {-9'd4,-10'd205};
ram[51594] = {-9'd1,-10'd202};
ram[51595] = {9'd2,-10'd198};
ram[51596] = {9'd5,-10'd195};
ram[51597] = {9'd8,-10'd192};
ram[51598] = {9'd11,-10'd189};
ram[51599] = {9'd14,-10'd186};
ram[51600] = {9'd18,-10'd183};
ram[51601] = {9'd21,-10'd180};
ram[51602] = {9'd24,-10'd176};
ram[51603] = {9'd27,-10'd173};
ram[51604] = {9'd30,-10'd170};
ram[51605] = {9'd33,-10'd167};
ram[51606] = {9'd36,-10'd164};
ram[51607] = {9'd40,-10'd161};
ram[51608] = {9'd43,-10'd158};
ram[51609] = {9'd46,-10'd154};
ram[51610] = {9'd49,-10'd151};
ram[51611] = {9'd52,-10'd148};
ram[51612] = {9'd55,-10'd145};
ram[51613] = {9'd58,-10'd142};
ram[51614] = {9'd62,-10'd139};
ram[51615] = {9'd65,-10'd136};
ram[51616] = {9'd68,-10'd132};
ram[51617] = {9'd71,-10'd129};
ram[51618] = {9'd74,-10'd126};
ram[51619] = {9'd77,-10'd123};
ram[51620] = {9'd80,-10'd120};
ram[51621] = {9'd84,-10'd117};
ram[51622] = {9'd87,-10'd114};
ram[51623] = {9'd90,-10'd110};
ram[51624] = {9'd93,-10'd107};
ram[51625] = {9'd96,-10'd104};
ram[51626] = {9'd99,-10'd101};
ram[51627] = {-9'd98,-10'd98};
ram[51628] = {-9'd95,-10'd95};
ram[51629] = {-9'd92,-10'd92};
ram[51630] = {-9'd88,-10'd88};
ram[51631] = {-9'd85,-10'd85};
ram[51632] = {-9'd82,-10'd82};
ram[51633] = {-9'd79,-10'd79};
ram[51634] = {-9'd76,-10'd76};
ram[51635] = {-9'd73,-10'd73};
ram[51636] = {-9'd70,-10'd70};
ram[51637] = {-9'd66,-10'd66};
ram[51638] = {-9'd63,-10'd63};
ram[51639] = {-9'd60,-10'd60};
ram[51640] = {-9'd57,-10'd57};
ram[51641] = {-9'd54,-10'd54};
ram[51642] = {-9'd51,-10'd51};
ram[51643] = {-9'd48,-10'd48};
ram[51644] = {-9'd44,-10'd44};
ram[51645] = {-9'd41,-10'd41};
ram[51646] = {-9'd38,-10'd38};
ram[51647] = {-9'd35,-10'd35};
ram[51648] = {-9'd32,-10'd32};
ram[51649] = {-9'd29,-10'd29};
ram[51650] = {-9'd26,-10'd26};
ram[51651] = {-9'd22,-10'd22};
ram[51652] = {-9'd19,-10'd19};
ram[51653] = {-9'd16,-10'd16};
ram[51654] = {-9'd13,-10'd13};
ram[51655] = {-9'd10,-10'd10};
ram[51656] = {-9'd7,-10'd7};
ram[51657] = {-9'd4,-10'd4};
ram[51658] = {9'd0,10'd0};
ram[51659] = {9'd3,10'd3};
ram[51660] = {9'd6,10'd6};
ram[51661] = {9'd9,10'd9};
ram[51662] = {9'd12,10'd12};
ram[51663] = {9'd15,10'd15};
ram[51664] = {9'd18,10'd18};
ram[51665] = {9'd21,10'd21};
ram[51666] = {9'd25,10'd25};
ram[51667] = {9'd28,10'd28};
ram[51668] = {9'd31,10'd31};
ram[51669] = {9'd34,10'd34};
ram[51670] = {9'd37,10'd37};
ram[51671] = {9'd40,10'd40};
ram[51672] = {9'd43,10'd43};
ram[51673] = {9'd47,10'd47};
ram[51674] = {9'd50,10'd50};
ram[51675] = {9'd53,10'd53};
ram[51676] = {9'd56,10'd56};
ram[51677] = {9'd59,10'd59};
ram[51678] = {9'd62,10'd62};
ram[51679] = {9'd65,10'd65};
ram[51680] = {9'd69,10'd69};
ram[51681] = {9'd72,10'd72};
ram[51682] = {9'd75,10'd75};
ram[51683] = {9'd78,10'd78};
ram[51684] = {9'd81,10'd81};
ram[51685] = {9'd84,10'd84};
ram[51686] = {9'd87,10'd87};
ram[51687] = {9'd91,10'd91};
ram[51688] = {9'd94,10'd94};
ram[51689] = {9'd97,10'd97};
ram[51690] = {-9'd100,10'd100};
ram[51691] = {-9'd97,10'd103};
ram[51692] = {-9'd94,10'd106};
ram[51693] = {-9'd91,10'd109};
ram[51694] = {-9'd88,10'd113};
ram[51695] = {-9'd85,10'd116};
ram[51696] = {-9'd81,10'd119};
ram[51697] = {-9'd78,10'd122};
ram[51698] = {-9'd75,10'd125};
ram[51699] = {-9'd72,10'd128};
ram[51700] = {-9'd69,10'd131};
ram[51701] = {-9'd66,10'd135};
ram[51702] = {-9'd63,10'd138};
ram[51703] = {-9'd59,10'd141};
ram[51704] = {-9'd56,10'd144};
ram[51705] = {-9'd53,10'd147};
ram[51706] = {-9'd50,10'd150};
ram[51707] = {-9'd47,10'd153};
ram[51708] = {-9'd44,10'd157};
ram[51709] = {-9'd41,10'd160};
ram[51710] = {-9'd37,10'd163};
ram[51711] = {-9'd34,10'd166};
ram[51712] = {-9'd34,10'd166};
ram[51713] = {-9'd31,10'd169};
ram[51714] = {-9'd28,10'd172};
ram[51715] = {-9'd25,10'd175};
ram[51716] = {-9'd22,10'd179};
ram[51717] = {-9'd19,10'd182};
ram[51718] = {-9'd15,10'd185};
ram[51719] = {-9'd12,10'd188};
ram[51720] = {-9'd9,10'd191};
ram[51721] = {-9'd6,10'd194};
ram[51722] = {-9'd3,10'd197};
ram[51723] = {9'd0,10'd201};
ram[51724] = {9'd3,10'd204};
ram[51725] = {9'd7,10'd207};
ram[51726] = {9'd10,10'd210};
ram[51727] = {9'd13,10'd213};
ram[51728] = {9'd16,10'd216};
ram[51729] = {9'd19,10'd219};
ram[51730] = {9'd22,10'd223};
ram[51731] = {9'd25,10'd226};
ram[51732] = {9'd29,10'd229};
ram[51733] = {9'd32,10'd232};
ram[51734] = {9'd35,10'd235};
ram[51735] = {9'd38,10'd238};
ram[51736] = {9'd41,10'd241};
ram[51737] = {9'd44,10'd245};
ram[51738] = {9'd47,10'd248};
ram[51739] = {9'd51,10'd251};
ram[51740] = {9'd54,10'd254};
ram[51741] = {9'd57,10'd257};
ram[51742] = {9'd60,10'd260};
ram[51743] = {9'd63,10'd263};
ram[51744] = {9'd66,10'd267};
ram[51745] = {9'd69,10'd270};
ram[51746] = {9'd73,10'd273};
ram[51747] = {9'd76,10'd276};
ram[51748] = {9'd79,10'd279};
ram[51749] = {9'd82,10'd282};
ram[51750] = {9'd85,10'd285};
ram[51751] = {9'd88,10'd289};
ram[51752] = {9'd91,10'd292};
ram[51753] = {9'd95,10'd295};
ram[51754] = {9'd98,10'd298};
ram[51755] = {-9'd99,10'd301};
ram[51756] = {-9'd96,10'd304};
ram[51757] = {-9'd93,10'd307};
ram[51758] = {-9'd90,10'd311};
ram[51759] = {-9'd87,10'd314};
ram[51760] = {-9'd84,10'd317};
ram[51761] = {-9'd81,10'd320};
ram[51762] = {-9'd77,10'd323};
ram[51763] = {-9'd74,10'd326};
ram[51764] = {-9'd71,10'd329};
ram[51765] = {-9'd68,10'd333};
ram[51766] = {-9'd65,10'd336};
ram[51767] = {-9'd62,10'd339};
ram[51768] = {-9'd59,10'd342};
ram[51769] = {-9'd55,10'd345};
ram[51770] = {-9'd52,10'd348};
ram[51771] = {-9'd49,10'd351};
ram[51772] = {-9'd46,10'd354};
ram[51773] = {-9'd43,10'd358};
ram[51774] = {-9'd40,10'd361};
ram[51775] = {-9'd37,10'd364};
ram[51776] = {-9'd33,10'd367};
ram[51777] = {-9'd30,10'd370};
ram[51778] = {-9'd27,10'd373};
ram[51779] = {-9'd24,10'd376};
ram[51780] = {-9'd21,10'd380};
ram[51781] = {-9'd18,10'd383};
ram[51782] = {-9'd15,10'd386};
ram[51783] = {-9'd11,10'd389};
ram[51784] = {-9'd8,10'd392};
ram[51785] = {-9'd5,10'd395};
ram[51786] = {-9'd2,10'd398};
ram[51787] = {9'd1,-10'd399};
ram[51788] = {9'd4,-10'd396};
ram[51789] = {9'd7,-10'd393};
ram[51790] = {9'd10,-10'd390};
ram[51791] = {9'd14,-10'd387};
ram[51792] = {9'd17,-10'd384};
ram[51793] = {9'd20,-10'd381};
ram[51794] = {9'd23,-10'd377};
ram[51795] = {9'd26,-10'd374};
ram[51796] = {9'd29,-10'd371};
ram[51797] = {9'd32,-10'd368};
ram[51798] = {9'd36,-10'd365};
ram[51799] = {9'd39,-10'd362};
ram[51800] = {9'd42,-10'd359};
ram[51801] = {9'd45,-10'd355};
ram[51802] = {9'd48,-10'd352};
ram[51803] = {9'd51,-10'd349};
ram[51804] = {9'd54,-10'd346};
ram[51805] = {9'd58,-10'd343};
ram[51806] = {9'd61,-10'd340};
ram[51807] = {9'd64,-10'd337};
ram[51808] = {9'd67,-10'd334};
ram[51809] = {9'd70,-10'd330};
ram[51810] = {9'd73,-10'd327};
ram[51811] = {9'd76,-10'd324};
ram[51812] = {9'd80,-10'd321};
ram[51813] = {9'd83,-10'd318};
ram[51814] = {9'd86,-10'd315};
ram[51815] = {9'd89,-10'd312};
ram[51816] = {9'd92,-10'd308};
ram[51817] = {9'd95,-10'd305};
ram[51818] = {9'd98,-10'd302};
ram[51819] = {-9'd99,-10'd299};
ram[51820] = {-9'd96,-10'd296};
ram[51821] = {-9'd92,-10'd293};
ram[51822] = {-9'd89,-10'd290};
ram[51823] = {-9'd86,-10'd286};
ram[51824] = {-9'd83,-10'd283};
ram[51825] = {-9'd80,-10'd280};
ram[51826] = {-9'd77,-10'd277};
ram[51827] = {-9'd74,-10'd274};
ram[51828] = {-9'd70,-10'd271};
ram[51829] = {-9'd67,-10'd268};
ram[51830] = {-9'd64,-10'd264};
ram[51831] = {-9'd61,-10'd261};
ram[51832] = {-9'd58,-10'd258};
ram[51833] = {-9'd55,-10'd255};
ram[51834] = {-9'd52,-10'd252};
ram[51835] = {-9'd48,-10'd249};
ram[51836] = {-9'd45,-10'd246};
ram[51837] = {-9'd42,-10'd242};
ram[51838] = {-9'd39,-10'd239};
ram[51839] = {-9'd36,-10'd236};
ram[51840] = {-9'd36,-10'd236};
ram[51841] = {-9'd33,-10'd233};
ram[51842] = {-9'd30,-10'd230};
ram[51843] = {-9'd26,-10'd227};
ram[51844] = {-9'd23,-10'd224};
ram[51845] = {-9'd20,-10'd220};
ram[51846] = {-9'd17,-10'd217};
ram[51847] = {-9'd14,-10'd214};
ram[51848] = {-9'd11,-10'd211};
ram[51849] = {-9'd8,-10'd208};
ram[51850] = {-9'd4,-10'd205};
ram[51851] = {-9'd1,-10'd202};
ram[51852] = {9'd2,-10'd198};
ram[51853] = {9'd5,-10'd195};
ram[51854] = {9'd8,-10'd192};
ram[51855] = {9'd11,-10'd189};
ram[51856] = {9'd14,-10'd186};
ram[51857] = {9'd18,-10'd183};
ram[51858] = {9'd21,-10'd180};
ram[51859] = {9'd24,-10'd176};
ram[51860] = {9'd27,-10'd173};
ram[51861] = {9'd30,-10'd170};
ram[51862] = {9'd33,-10'd167};
ram[51863] = {9'd36,-10'd164};
ram[51864] = {9'd40,-10'd161};
ram[51865] = {9'd43,-10'd158};
ram[51866] = {9'd46,-10'd154};
ram[51867] = {9'd49,-10'd151};
ram[51868] = {9'd52,-10'd148};
ram[51869] = {9'd55,-10'd145};
ram[51870] = {9'd58,-10'd142};
ram[51871] = {9'd62,-10'd139};
ram[51872] = {9'd65,-10'd136};
ram[51873] = {9'd68,-10'd132};
ram[51874] = {9'd71,-10'd129};
ram[51875] = {9'd74,-10'd126};
ram[51876] = {9'd77,-10'd123};
ram[51877] = {9'd80,-10'd120};
ram[51878] = {9'd84,-10'd117};
ram[51879] = {9'd87,-10'd114};
ram[51880] = {9'd90,-10'd110};
ram[51881] = {9'd93,-10'd107};
ram[51882] = {9'd96,-10'd104};
ram[51883] = {9'd99,-10'd101};
ram[51884] = {-9'd98,-10'd98};
ram[51885] = {-9'd95,-10'd95};
ram[51886] = {-9'd92,-10'd92};
ram[51887] = {-9'd88,-10'd88};
ram[51888] = {-9'd85,-10'd85};
ram[51889] = {-9'd82,-10'd82};
ram[51890] = {-9'd79,-10'd79};
ram[51891] = {-9'd76,-10'd76};
ram[51892] = {-9'd73,-10'd73};
ram[51893] = {-9'd70,-10'd70};
ram[51894] = {-9'd66,-10'd66};
ram[51895] = {-9'd63,-10'd63};
ram[51896] = {-9'd60,-10'd60};
ram[51897] = {-9'd57,-10'd57};
ram[51898] = {-9'd54,-10'd54};
ram[51899] = {-9'd51,-10'd51};
ram[51900] = {-9'd48,-10'd48};
ram[51901] = {-9'd44,-10'd44};
ram[51902] = {-9'd41,-10'd41};
ram[51903] = {-9'd38,-10'd38};
ram[51904] = {-9'd35,-10'd35};
ram[51905] = {-9'd32,-10'd32};
ram[51906] = {-9'd29,-10'd29};
ram[51907] = {-9'd26,-10'd26};
ram[51908] = {-9'd22,-10'd22};
ram[51909] = {-9'd19,-10'd19};
ram[51910] = {-9'd16,-10'd16};
ram[51911] = {-9'd13,-10'd13};
ram[51912] = {-9'd10,-10'd10};
ram[51913] = {-9'd7,-10'd7};
ram[51914] = {-9'd4,-10'd4};
ram[51915] = {9'd0,10'd0};
ram[51916] = {9'd3,10'd3};
ram[51917] = {9'd6,10'd6};
ram[51918] = {9'd9,10'd9};
ram[51919] = {9'd12,10'd12};
ram[51920] = {9'd15,10'd15};
ram[51921] = {9'd18,10'd18};
ram[51922] = {9'd21,10'd21};
ram[51923] = {9'd25,10'd25};
ram[51924] = {9'd28,10'd28};
ram[51925] = {9'd31,10'd31};
ram[51926] = {9'd34,10'd34};
ram[51927] = {9'd37,10'd37};
ram[51928] = {9'd40,10'd40};
ram[51929] = {9'd43,10'd43};
ram[51930] = {9'd47,10'd47};
ram[51931] = {9'd50,10'd50};
ram[51932] = {9'd53,10'd53};
ram[51933] = {9'd56,10'd56};
ram[51934] = {9'd59,10'd59};
ram[51935] = {9'd62,10'd62};
ram[51936] = {9'd65,10'd65};
ram[51937] = {9'd69,10'd69};
ram[51938] = {9'd72,10'd72};
ram[51939] = {9'd75,10'd75};
ram[51940] = {9'd78,10'd78};
ram[51941] = {9'd81,10'd81};
ram[51942] = {9'd84,10'd84};
ram[51943] = {9'd87,10'd87};
ram[51944] = {9'd91,10'd91};
ram[51945] = {9'd94,10'd94};
ram[51946] = {9'd97,10'd97};
ram[51947] = {-9'd100,10'd100};
ram[51948] = {-9'd97,10'd103};
ram[51949] = {-9'd94,10'd106};
ram[51950] = {-9'd91,10'd109};
ram[51951] = {-9'd88,10'd113};
ram[51952] = {-9'd85,10'd116};
ram[51953] = {-9'd81,10'd119};
ram[51954] = {-9'd78,10'd122};
ram[51955] = {-9'd75,10'd125};
ram[51956] = {-9'd72,10'd128};
ram[51957] = {-9'd69,10'd131};
ram[51958] = {-9'd66,10'd135};
ram[51959] = {-9'd63,10'd138};
ram[51960] = {-9'd59,10'd141};
ram[51961] = {-9'd56,10'd144};
ram[51962] = {-9'd53,10'd147};
ram[51963] = {-9'd50,10'd150};
ram[51964] = {-9'd47,10'd153};
ram[51965] = {-9'd44,10'd157};
ram[51966] = {-9'd41,10'd160};
ram[51967] = {-9'd37,10'd163};
ram[51968] = {-9'd37,10'd163};
ram[51969] = {-9'd34,10'd166};
ram[51970] = {-9'd31,10'd169};
ram[51971] = {-9'd28,10'd172};
ram[51972] = {-9'd25,10'd175};
ram[51973] = {-9'd22,10'd179};
ram[51974] = {-9'd19,10'd182};
ram[51975] = {-9'd15,10'd185};
ram[51976] = {-9'd12,10'd188};
ram[51977] = {-9'd9,10'd191};
ram[51978] = {-9'd6,10'd194};
ram[51979] = {-9'd3,10'd197};
ram[51980] = {9'd0,10'd201};
ram[51981] = {9'd3,10'd204};
ram[51982] = {9'd7,10'd207};
ram[51983] = {9'd10,10'd210};
ram[51984] = {9'd13,10'd213};
ram[51985] = {9'd16,10'd216};
ram[51986] = {9'd19,10'd219};
ram[51987] = {9'd22,10'd223};
ram[51988] = {9'd25,10'd226};
ram[51989] = {9'd29,10'd229};
ram[51990] = {9'd32,10'd232};
ram[51991] = {9'd35,10'd235};
ram[51992] = {9'd38,10'd238};
ram[51993] = {9'd41,10'd241};
ram[51994] = {9'd44,10'd245};
ram[51995] = {9'd47,10'd248};
ram[51996] = {9'd51,10'd251};
ram[51997] = {9'd54,10'd254};
ram[51998] = {9'd57,10'd257};
ram[51999] = {9'd60,10'd260};
ram[52000] = {9'd63,10'd263};
ram[52001] = {9'd66,10'd267};
ram[52002] = {9'd69,10'd270};
ram[52003] = {9'd73,10'd273};
ram[52004] = {9'd76,10'd276};
ram[52005] = {9'd79,10'd279};
ram[52006] = {9'd82,10'd282};
ram[52007] = {9'd85,10'd285};
ram[52008] = {9'd88,10'd289};
ram[52009] = {9'd91,10'd292};
ram[52010] = {9'd95,10'd295};
ram[52011] = {9'd98,10'd298};
ram[52012] = {-9'd99,10'd301};
ram[52013] = {-9'd96,10'd304};
ram[52014] = {-9'd93,10'd307};
ram[52015] = {-9'd90,10'd311};
ram[52016] = {-9'd87,10'd314};
ram[52017] = {-9'd84,10'd317};
ram[52018] = {-9'd81,10'd320};
ram[52019] = {-9'd77,10'd323};
ram[52020] = {-9'd74,10'd326};
ram[52021] = {-9'd71,10'd329};
ram[52022] = {-9'd68,10'd333};
ram[52023] = {-9'd65,10'd336};
ram[52024] = {-9'd62,10'd339};
ram[52025] = {-9'd59,10'd342};
ram[52026] = {-9'd55,10'd345};
ram[52027] = {-9'd52,10'd348};
ram[52028] = {-9'd49,10'd351};
ram[52029] = {-9'd46,10'd354};
ram[52030] = {-9'd43,10'd358};
ram[52031] = {-9'd40,10'd361};
ram[52032] = {-9'd37,10'd364};
ram[52033] = {-9'd33,10'd367};
ram[52034] = {-9'd30,10'd370};
ram[52035] = {-9'd27,10'd373};
ram[52036] = {-9'd24,10'd376};
ram[52037] = {-9'd21,10'd380};
ram[52038] = {-9'd18,10'd383};
ram[52039] = {-9'd15,10'd386};
ram[52040] = {-9'd11,10'd389};
ram[52041] = {-9'd8,10'd392};
ram[52042] = {-9'd5,10'd395};
ram[52043] = {-9'd2,10'd398};
ram[52044] = {9'd1,-10'd399};
ram[52045] = {9'd4,-10'd396};
ram[52046] = {9'd7,-10'd393};
ram[52047] = {9'd10,-10'd390};
ram[52048] = {9'd14,-10'd387};
ram[52049] = {9'd17,-10'd384};
ram[52050] = {9'd20,-10'd381};
ram[52051] = {9'd23,-10'd377};
ram[52052] = {9'd26,-10'd374};
ram[52053] = {9'd29,-10'd371};
ram[52054] = {9'd32,-10'd368};
ram[52055] = {9'd36,-10'd365};
ram[52056] = {9'd39,-10'd362};
ram[52057] = {9'd42,-10'd359};
ram[52058] = {9'd45,-10'd355};
ram[52059] = {9'd48,-10'd352};
ram[52060] = {9'd51,-10'd349};
ram[52061] = {9'd54,-10'd346};
ram[52062] = {9'd58,-10'd343};
ram[52063] = {9'd61,-10'd340};
ram[52064] = {9'd64,-10'd337};
ram[52065] = {9'd67,-10'd334};
ram[52066] = {9'd70,-10'd330};
ram[52067] = {9'd73,-10'd327};
ram[52068] = {9'd76,-10'd324};
ram[52069] = {9'd80,-10'd321};
ram[52070] = {9'd83,-10'd318};
ram[52071] = {9'd86,-10'd315};
ram[52072] = {9'd89,-10'd312};
ram[52073] = {9'd92,-10'd308};
ram[52074] = {9'd95,-10'd305};
ram[52075] = {9'd98,-10'd302};
ram[52076] = {-9'd99,-10'd299};
ram[52077] = {-9'd96,-10'd296};
ram[52078] = {-9'd92,-10'd293};
ram[52079] = {-9'd89,-10'd290};
ram[52080] = {-9'd86,-10'd286};
ram[52081] = {-9'd83,-10'd283};
ram[52082] = {-9'd80,-10'd280};
ram[52083] = {-9'd77,-10'd277};
ram[52084] = {-9'd74,-10'd274};
ram[52085] = {-9'd70,-10'd271};
ram[52086] = {-9'd67,-10'd268};
ram[52087] = {-9'd64,-10'd264};
ram[52088] = {-9'd61,-10'd261};
ram[52089] = {-9'd58,-10'd258};
ram[52090] = {-9'd55,-10'd255};
ram[52091] = {-9'd52,-10'd252};
ram[52092] = {-9'd48,-10'd249};
ram[52093] = {-9'd45,-10'd246};
ram[52094] = {-9'd42,-10'd242};
ram[52095] = {-9'd39,-10'd239};
ram[52096] = {-9'd39,-10'd239};
ram[52097] = {-9'd36,-10'd236};
ram[52098] = {-9'd33,-10'd233};
ram[52099] = {-9'd30,-10'd230};
ram[52100] = {-9'd26,-10'd227};
ram[52101] = {-9'd23,-10'd224};
ram[52102] = {-9'd20,-10'd220};
ram[52103] = {-9'd17,-10'd217};
ram[52104] = {-9'd14,-10'd214};
ram[52105] = {-9'd11,-10'd211};
ram[52106] = {-9'd8,-10'd208};
ram[52107] = {-9'd4,-10'd205};
ram[52108] = {-9'd1,-10'd202};
ram[52109] = {9'd2,-10'd198};
ram[52110] = {9'd5,-10'd195};
ram[52111] = {9'd8,-10'd192};
ram[52112] = {9'd11,-10'd189};
ram[52113] = {9'd14,-10'd186};
ram[52114] = {9'd18,-10'd183};
ram[52115] = {9'd21,-10'd180};
ram[52116] = {9'd24,-10'd176};
ram[52117] = {9'd27,-10'd173};
ram[52118] = {9'd30,-10'd170};
ram[52119] = {9'd33,-10'd167};
ram[52120] = {9'd36,-10'd164};
ram[52121] = {9'd40,-10'd161};
ram[52122] = {9'd43,-10'd158};
ram[52123] = {9'd46,-10'd154};
ram[52124] = {9'd49,-10'd151};
ram[52125] = {9'd52,-10'd148};
ram[52126] = {9'd55,-10'd145};
ram[52127] = {9'd58,-10'd142};
ram[52128] = {9'd62,-10'd139};
ram[52129] = {9'd65,-10'd136};
ram[52130] = {9'd68,-10'd132};
ram[52131] = {9'd71,-10'd129};
ram[52132] = {9'd74,-10'd126};
ram[52133] = {9'd77,-10'd123};
ram[52134] = {9'd80,-10'd120};
ram[52135] = {9'd84,-10'd117};
ram[52136] = {9'd87,-10'd114};
ram[52137] = {9'd90,-10'd110};
ram[52138] = {9'd93,-10'd107};
ram[52139] = {9'd96,-10'd104};
ram[52140] = {9'd99,-10'd101};
ram[52141] = {-9'd98,-10'd98};
ram[52142] = {-9'd95,-10'd95};
ram[52143] = {-9'd92,-10'd92};
ram[52144] = {-9'd88,-10'd88};
ram[52145] = {-9'd85,-10'd85};
ram[52146] = {-9'd82,-10'd82};
ram[52147] = {-9'd79,-10'd79};
ram[52148] = {-9'd76,-10'd76};
ram[52149] = {-9'd73,-10'd73};
ram[52150] = {-9'd70,-10'd70};
ram[52151] = {-9'd66,-10'd66};
ram[52152] = {-9'd63,-10'd63};
ram[52153] = {-9'd60,-10'd60};
ram[52154] = {-9'd57,-10'd57};
ram[52155] = {-9'd54,-10'd54};
ram[52156] = {-9'd51,-10'd51};
ram[52157] = {-9'd48,-10'd48};
ram[52158] = {-9'd44,-10'd44};
ram[52159] = {-9'd41,-10'd41};
ram[52160] = {-9'd38,-10'd38};
ram[52161] = {-9'd35,-10'd35};
ram[52162] = {-9'd32,-10'd32};
ram[52163] = {-9'd29,-10'd29};
ram[52164] = {-9'd26,-10'd26};
ram[52165] = {-9'd22,-10'd22};
ram[52166] = {-9'd19,-10'd19};
ram[52167] = {-9'd16,-10'd16};
ram[52168] = {-9'd13,-10'd13};
ram[52169] = {-9'd10,-10'd10};
ram[52170] = {-9'd7,-10'd7};
ram[52171] = {-9'd4,-10'd4};
ram[52172] = {9'd0,10'd0};
ram[52173] = {9'd3,10'd3};
ram[52174] = {9'd6,10'd6};
ram[52175] = {9'd9,10'd9};
ram[52176] = {9'd12,10'd12};
ram[52177] = {9'd15,10'd15};
ram[52178] = {9'd18,10'd18};
ram[52179] = {9'd21,10'd21};
ram[52180] = {9'd25,10'd25};
ram[52181] = {9'd28,10'd28};
ram[52182] = {9'd31,10'd31};
ram[52183] = {9'd34,10'd34};
ram[52184] = {9'd37,10'd37};
ram[52185] = {9'd40,10'd40};
ram[52186] = {9'd43,10'd43};
ram[52187] = {9'd47,10'd47};
ram[52188] = {9'd50,10'd50};
ram[52189] = {9'd53,10'd53};
ram[52190] = {9'd56,10'd56};
ram[52191] = {9'd59,10'd59};
ram[52192] = {9'd62,10'd62};
ram[52193] = {9'd65,10'd65};
ram[52194] = {9'd69,10'd69};
ram[52195] = {9'd72,10'd72};
ram[52196] = {9'd75,10'd75};
ram[52197] = {9'd78,10'd78};
ram[52198] = {9'd81,10'd81};
ram[52199] = {9'd84,10'd84};
ram[52200] = {9'd87,10'd87};
ram[52201] = {9'd91,10'd91};
ram[52202] = {9'd94,10'd94};
ram[52203] = {9'd97,10'd97};
ram[52204] = {-9'd100,10'd100};
ram[52205] = {-9'd97,10'd103};
ram[52206] = {-9'd94,10'd106};
ram[52207] = {-9'd91,10'd109};
ram[52208] = {-9'd88,10'd113};
ram[52209] = {-9'd85,10'd116};
ram[52210] = {-9'd81,10'd119};
ram[52211] = {-9'd78,10'd122};
ram[52212] = {-9'd75,10'd125};
ram[52213] = {-9'd72,10'd128};
ram[52214] = {-9'd69,10'd131};
ram[52215] = {-9'd66,10'd135};
ram[52216] = {-9'd63,10'd138};
ram[52217] = {-9'd59,10'd141};
ram[52218] = {-9'd56,10'd144};
ram[52219] = {-9'd53,10'd147};
ram[52220] = {-9'd50,10'd150};
ram[52221] = {-9'd47,10'd153};
ram[52222] = {-9'd44,10'd157};
ram[52223] = {-9'd41,10'd160};
ram[52224] = {-9'd41,10'd160};
ram[52225] = {-9'd37,10'd163};
ram[52226] = {-9'd34,10'd166};
ram[52227] = {-9'd31,10'd169};
ram[52228] = {-9'd28,10'd172};
ram[52229] = {-9'd25,10'd175};
ram[52230] = {-9'd22,10'd179};
ram[52231] = {-9'd19,10'd182};
ram[52232] = {-9'd15,10'd185};
ram[52233] = {-9'd12,10'd188};
ram[52234] = {-9'd9,10'd191};
ram[52235] = {-9'd6,10'd194};
ram[52236] = {-9'd3,10'd197};
ram[52237] = {9'd0,10'd201};
ram[52238] = {9'd3,10'd204};
ram[52239] = {9'd7,10'd207};
ram[52240] = {9'd10,10'd210};
ram[52241] = {9'd13,10'd213};
ram[52242] = {9'd16,10'd216};
ram[52243] = {9'd19,10'd219};
ram[52244] = {9'd22,10'd223};
ram[52245] = {9'd25,10'd226};
ram[52246] = {9'd29,10'd229};
ram[52247] = {9'd32,10'd232};
ram[52248] = {9'd35,10'd235};
ram[52249] = {9'd38,10'd238};
ram[52250] = {9'd41,10'd241};
ram[52251] = {9'd44,10'd245};
ram[52252] = {9'd47,10'd248};
ram[52253] = {9'd51,10'd251};
ram[52254] = {9'd54,10'd254};
ram[52255] = {9'd57,10'd257};
ram[52256] = {9'd60,10'd260};
ram[52257] = {9'd63,10'd263};
ram[52258] = {9'd66,10'd267};
ram[52259] = {9'd69,10'd270};
ram[52260] = {9'd73,10'd273};
ram[52261] = {9'd76,10'd276};
ram[52262] = {9'd79,10'd279};
ram[52263] = {9'd82,10'd282};
ram[52264] = {9'd85,10'd285};
ram[52265] = {9'd88,10'd289};
ram[52266] = {9'd91,10'd292};
ram[52267] = {9'd95,10'd295};
ram[52268] = {9'd98,10'd298};
ram[52269] = {-9'd99,10'd301};
ram[52270] = {-9'd96,10'd304};
ram[52271] = {-9'd93,10'd307};
ram[52272] = {-9'd90,10'd311};
ram[52273] = {-9'd87,10'd314};
ram[52274] = {-9'd84,10'd317};
ram[52275] = {-9'd81,10'd320};
ram[52276] = {-9'd77,10'd323};
ram[52277] = {-9'd74,10'd326};
ram[52278] = {-9'd71,10'd329};
ram[52279] = {-9'd68,10'd333};
ram[52280] = {-9'd65,10'd336};
ram[52281] = {-9'd62,10'd339};
ram[52282] = {-9'd59,10'd342};
ram[52283] = {-9'd55,10'd345};
ram[52284] = {-9'd52,10'd348};
ram[52285] = {-9'd49,10'd351};
ram[52286] = {-9'd46,10'd354};
ram[52287] = {-9'd43,10'd358};
ram[52288] = {-9'd40,10'd361};
ram[52289] = {-9'd37,10'd364};
ram[52290] = {-9'd33,10'd367};
ram[52291] = {-9'd30,10'd370};
ram[52292] = {-9'd27,10'd373};
ram[52293] = {-9'd24,10'd376};
ram[52294] = {-9'd21,10'd380};
ram[52295] = {-9'd18,10'd383};
ram[52296] = {-9'd15,10'd386};
ram[52297] = {-9'd11,10'd389};
ram[52298] = {-9'd8,10'd392};
ram[52299] = {-9'd5,10'd395};
ram[52300] = {-9'd2,10'd398};
ram[52301] = {9'd1,-10'd399};
ram[52302] = {9'd4,-10'd396};
ram[52303] = {9'd7,-10'd393};
ram[52304] = {9'd10,-10'd390};
ram[52305] = {9'd14,-10'd387};
ram[52306] = {9'd17,-10'd384};
ram[52307] = {9'd20,-10'd381};
ram[52308] = {9'd23,-10'd377};
ram[52309] = {9'd26,-10'd374};
ram[52310] = {9'd29,-10'd371};
ram[52311] = {9'd32,-10'd368};
ram[52312] = {9'd36,-10'd365};
ram[52313] = {9'd39,-10'd362};
ram[52314] = {9'd42,-10'd359};
ram[52315] = {9'd45,-10'd355};
ram[52316] = {9'd48,-10'd352};
ram[52317] = {9'd51,-10'd349};
ram[52318] = {9'd54,-10'd346};
ram[52319] = {9'd58,-10'd343};
ram[52320] = {9'd61,-10'd340};
ram[52321] = {9'd64,-10'd337};
ram[52322] = {9'd67,-10'd334};
ram[52323] = {9'd70,-10'd330};
ram[52324] = {9'd73,-10'd327};
ram[52325] = {9'd76,-10'd324};
ram[52326] = {9'd80,-10'd321};
ram[52327] = {9'd83,-10'd318};
ram[52328] = {9'd86,-10'd315};
ram[52329] = {9'd89,-10'd312};
ram[52330] = {9'd92,-10'd308};
ram[52331] = {9'd95,-10'd305};
ram[52332] = {9'd98,-10'd302};
ram[52333] = {-9'd99,-10'd299};
ram[52334] = {-9'd96,-10'd296};
ram[52335] = {-9'd92,-10'd293};
ram[52336] = {-9'd89,-10'd290};
ram[52337] = {-9'd86,-10'd286};
ram[52338] = {-9'd83,-10'd283};
ram[52339] = {-9'd80,-10'd280};
ram[52340] = {-9'd77,-10'd277};
ram[52341] = {-9'd74,-10'd274};
ram[52342] = {-9'd70,-10'd271};
ram[52343] = {-9'd67,-10'd268};
ram[52344] = {-9'd64,-10'd264};
ram[52345] = {-9'd61,-10'd261};
ram[52346] = {-9'd58,-10'd258};
ram[52347] = {-9'd55,-10'd255};
ram[52348] = {-9'd52,-10'd252};
ram[52349] = {-9'd48,-10'd249};
ram[52350] = {-9'd45,-10'd246};
ram[52351] = {-9'd42,-10'd242};
ram[52352] = {-9'd42,-10'd242};
ram[52353] = {-9'd39,-10'd239};
ram[52354] = {-9'd36,-10'd236};
ram[52355] = {-9'd33,-10'd233};
ram[52356] = {-9'd30,-10'd230};
ram[52357] = {-9'd26,-10'd227};
ram[52358] = {-9'd23,-10'd224};
ram[52359] = {-9'd20,-10'd220};
ram[52360] = {-9'd17,-10'd217};
ram[52361] = {-9'd14,-10'd214};
ram[52362] = {-9'd11,-10'd211};
ram[52363] = {-9'd8,-10'd208};
ram[52364] = {-9'd4,-10'd205};
ram[52365] = {-9'd1,-10'd202};
ram[52366] = {9'd2,-10'd198};
ram[52367] = {9'd5,-10'd195};
ram[52368] = {9'd8,-10'd192};
ram[52369] = {9'd11,-10'd189};
ram[52370] = {9'd14,-10'd186};
ram[52371] = {9'd18,-10'd183};
ram[52372] = {9'd21,-10'd180};
ram[52373] = {9'd24,-10'd176};
ram[52374] = {9'd27,-10'd173};
ram[52375] = {9'd30,-10'd170};
ram[52376] = {9'd33,-10'd167};
ram[52377] = {9'd36,-10'd164};
ram[52378] = {9'd40,-10'd161};
ram[52379] = {9'd43,-10'd158};
ram[52380] = {9'd46,-10'd154};
ram[52381] = {9'd49,-10'd151};
ram[52382] = {9'd52,-10'd148};
ram[52383] = {9'd55,-10'd145};
ram[52384] = {9'd58,-10'd142};
ram[52385] = {9'd62,-10'd139};
ram[52386] = {9'd65,-10'd136};
ram[52387] = {9'd68,-10'd132};
ram[52388] = {9'd71,-10'd129};
ram[52389] = {9'd74,-10'd126};
ram[52390] = {9'd77,-10'd123};
ram[52391] = {9'd80,-10'd120};
ram[52392] = {9'd84,-10'd117};
ram[52393] = {9'd87,-10'd114};
ram[52394] = {9'd90,-10'd110};
ram[52395] = {9'd93,-10'd107};
ram[52396] = {9'd96,-10'd104};
ram[52397] = {9'd99,-10'd101};
ram[52398] = {-9'd98,-10'd98};
ram[52399] = {-9'd95,-10'd95};
ram[52400] = {-9'd92,-10'd92};
ram[52401] = {-9'd88,-10'd88};
ram[52402] = {-9'd85,-10'd85};
ram[52403] = {-9'd82,-10'd82};
ram[52404] = {-9'd79,-10'd79};
ram[52405] = {-9'd76,-10'd76};
ram[52406] = {-9'd73,-10'd73};
ram[52407] = {-9'd70,-10'd70};
ram[52408] = {-9'd66,-10'd66};
ram[52409] = {-9'd63,-10'd63};
ram[52410] = {-9'd60,-10'd60};
ram[52411] = {-9'd57,-10'd57};
ram[52412] = {-9'd54,-10'd54};
ram[52413] = {-9'd51,-10'd51};
ram[52414] = {-9'd48,-10'd48};
ram[52415] = {-9'd44,-10'd44};
ram[52416] = {-9'd41,-10'd41};
ram[52417] = {-9'd38,-10'd38};
ram[52418] = {-9'd35,-10'd35};
ram[52419] = {-9'd32,-10'd32};
ram[52420] = {-9'd29,-10'd29};
ram[52421] = {-9'd26,-10'd26};
ram[52422] = {-9'd22,-10'd22};
ram[52423] = {-9'd19,-10'd19};
ram[52424] = {-9'd16,-10'd16};
ram[52425] = {-9'd13,-10'd13};
ram[52426] = {-9'd10,-10'd10};
ram[52427] = {-9'd7,-10'd7};
ram[52428] = {-9'd4,-10'd4};
ram[52429] = {9'd0,10'd0};
ram[52430] = {9'd3,10'd3};
ram[52431] = {9'd6,10'd6};
ram[52432] = {9'd9,10'd9};
ram[52433] = {9'd12,10'd12};
ram[52434] = {9'd15,10'd15};
ram[52435] = {9'd18,10'd18};
ram[52436] = {9'd21,10'd21};
ram[52437] = {9'd25,10'd25};
ram[52438] = {9'd28,10'd28};
ram[52439] = {9'd31,10'd31};
ram[52440] = {9'd34,10'd34};
ram[52441] = {9'd37,10'd37};
ram[52442] = {9'd40,10'd40};
ram[52443] = {9'd43,10'd43};
ram[52444] = {9'd47,10'd47};
ram[52445] = {9'd50,10'd50};
ram[52446] = {9'd53,10'd53};
ram[52447] = {9'd56,10'd56};
ram[52448] = {9'd59,10'd59};
ram[52449] = {9'd62,10'd62};
ram[52450] = {9'd65,10'd65};
ram[52451] = {9'd69,10'd69};
ram[52452] = {9'd72,10'd72};
ram[52453] = {9'd75,10'd75};
ram[52454] = {9'd78,10'd78};
ram[52455] = {9'd81,10'd81};
ram[52456] = {9'd84,10'd84};
ram[52457] = {9'd87,10'd87};
ram[52458] = {9'd91,10'd91};
ram[52459] = {9'd94,10'd94};
ram[52460] = {9'd97,10'd97};
ram[52461] = {-9'd100,10'd100};
ram[52462] = {-9'd97,10'd103};
ram[52463] = {-9'd94,10'd106};
ram[52464] = {-9'd91,10'd109};
ram[52465] = {-9'd88,10'd113};
ram[52466] = {-9'd85,10'd116};
ram[52467] = {-9'd81,10'd119};
ram[52468] = {-9'd78,10'd122};
ram[52469] = {-9'd75,10'd125};
ram[52470] = {-9'd72,10'd128};
ram[52471] = {-9'd69,10'd131};
ram[52472] = {-9'd66,10'd135};
ram[52473] = {-9'd63,10'd138};
ram[52474] = {-9'd59,10'd141};
ram[52475] = {-9'd56,10'd144};
ram[52476] = {-9'd53,10'd147};
ram[52477] = {-9'd50,10'd150};
ram[52478] = {-9'd47,10'd153};
ram[52479] = {-9'd44,10'd157};
ram[52480] = {-9'd44,10'd157};
ram[52481] = {-9'd41,10'd160};
ram[52482] = {-9'd37,10'd163};
ram[52483] = {-9'd34,10'd166};
ram[52484] = {-9'd31,10'd169};
ram[52485] = {-9'd28,10'd172};
ram[52486] = {-9'd25,10'd175};
ram[52487] = {-9'd22,10'd179};
ram[52488] = {-9'd19,10'd182};
ram[52489] = {-9'd15,10'd185};
ram[52490] = {-9'd12,10'd188};
ram[52491] = {-9'd9,10'd191};
ram[52492] = {-9'd6,10'd194};
ram[52493] = {-9'd3,10'd197};
ram[52494] = {9'd0,10'd201};
ram[52495] = {9'd3,10'd204};
ram[52496] = {9'd7,10'd207};
ram[52497] = {9'd10,10'd210};
ram[52498] = {9'd13,10'd213};
ram[52499] = {9'd16,10'd216};
ram[52500] = {9'd19,10'd219};
ram[52501] = {9'd22,10'd223};
ram[52502] = {9'd25,10'd226};
ram[52503] = {9'd29,10'd229};
ram[52504] = {9'd32,10'd232};
ram[52505] = {9'd35,10'd235};
ram[52506] = {9'd38,10'd238};
ram[52507] = {9'd41,10'd241};
ram[52508] = {9'd44,10'd245};
ram[52509] = {9'd47,10'd248};
ram[52510] = {9'd51,10'd251};
ram[52511] = {9'd54,10'd254};
ram[52512] = {9'd57,10'd257};
ram[52513] = {9'd60,10'd260};
ram[52514] = {9'd63,10'd263};
ram[52515] = {9'd66,10'd267};
ram[52516] = {9'd69,10'd270};
ram[52517] = {9'd73,10'd273};
ram[52518] = {9'd76,10'd276};
ram[52519] = {9'd79,10'd279};
ram[52520] = {9'd82,10'd282};
ram[52521] = {9'd85,10'd285};
ram[52522] = {9'd88,10'd289};
ram[52523] = {9'd91,10'd292};
ram[52524] = {9'd95,10'd295};
ram[52525] = {9'd98,10'd298};
ram[52526] = {-9'd99,10'd301};
ram[52527] = {-9'd96,10'd304};
ram[52528] = {-9'd93,10'd307};
ram[52529] = {-9'd90,10'd311};
ram[52530] = {-9'd87,10'd314};
ram[52531] = {-9'd84,10'd317};
ram[52532] = {-9'd81,10'd320};
ram[52533] = {-9'd77,10'd323};
ram[52534] = {-9'd74,10'd326};
ram[52535] = {-9'd71,10'd329};
ram[52536] = {-9'd68,10'd333};
ram[52537] = {-9'd65,10'd336};
ram[52538] = {-9'd62,10'd339};
ram[52539] = {-9'd59,10'd342};
ram[52540] = {-9'd55,10'd345};
ram[52541] = {-9'd52,10'd348};
ram[52542] = {-9'd49,10'd351};
ram[52543] = {-9'd46,10'd354};
ram[52544] = {-9'd43,10'd358};
ram[52545] = {-9'd40,10'd361};
ram[52546] = {-9'd37,10'd364};
ram[52547] = {-9'd33,10'd367};
ram[52548] = {-9'd30,10'd370};
ram[52549] = {-9'd27,10'd373};
ram[52550] = {-9'd24,10'd376};
ram[52551] = {-9'd21,10'd380};
ram[52552] = {-9'd18,10'd383};
ram[52553] = {-9'd15,10'd386};
ram[52554] = {-9'd11,10'd389};
ram[52555] = {-9'd8,10'd392};
ram[52556] = {-9'd5,10'd395};
ram[52557] = {-9'd2,10'd398};
ram[52558] = {9'd1,-10'd399};
ram[52559] = {9'd4,-10'd396};
ram[52560] = {9'd7,-10'd393};
ram[52561] = {9'd10,-10'd390};
ram[52562] = {9'd14,-10'd387};
ram[52563] = {9'd17,-10'd384};
ram[52564] = {9'd20,-10'd381};
ram[52565] = {9'd23,-10'd377};
ram[52566] = {9'd26,-10'd374};
ram[52567] = {9'd29,-10'd371};
ram[52568] = {9'd32,-10'd368};
ram[52569] = {9'd36,-10'd365};
ram[52570] = {9'd39,-10'd362};
ram[52571] = {9'd42,-10'd359};
ram[52572] = {9'd45,-10'd355};
ram[52573] = {9'd48,-10'd352};
ram[52574] = {9'd51,-10'd349};
ram[52575] = {9'd54,-10'd346};
ram[52576] = {9'd58,-10'd343};
ram[52577] = {9'd61,-10'd340};
ram[52578] = {9'd64,-10'd337};
ram[52579] = {9'd67,-10'd334};
ram[52580] = {9'd70,-10'd330};
ram[52581] = {9'd73,-10'd327};
ram[52582] = {9'd76,-10'd324};
ram[52583] = {9'd80,-10'd321};
ram[52584] = {9'd83,-10'd318};
ram[52585] = {9'd86,-10'd315};
ram[52586] = {9'd89,-10'd312};
ram[52587] = {9'd92,-10'd308};
ram[52588] = {9'd95,-10'd305};
ram[52589] = {9'd98,-10'd302};
ram[52590] = {-9'd99,-10'd299};
ram[52591] = {-9'd96,-10'd296};
ram[52592] = {-9'd92,-10'd293};
ram[52593] = {-9'd89,-10'd290};
ram[52594] = {-9'd86,-10'd286};
ram[52595] = {-9'd83,-10'd283};
ram[52596] = {-9'd80,-10'd280};
ram[52597] = {-9'd77,-10'd277};
ram[52598] = {-9'd74,-10'd274};
ram[52599] = {-9'd70,-10'd271};
ram[52600] = {-9'd67,-10'd268};
ram[52601] = {-9'd64,-10'd264};
ram[52602] = {-9'd61,-10'd261};
ram[52603] = {-9'd58,-10'd258};
ram[52604] = {-9'd55,-10'd255};
ram[52605] = {-9'd52,-10'd252};
ram[52606] = {-9'd48,-10'd249};
ram[52607] = {-9'd45,-10'd246};
ram[52608] = {-9'd45,-10'd246};
ram[52609] = {-9'd42,-10'd242};
ram[52610] = {-9'd39,-10'd239};
ram[52611] = {-9'd36,-10'd236};
ram[52612] = {-9'd33,-10'd233};
ram[52613] = {-9'd30,-10'd230};
ram[52614] = {-9'd26,-10'd227};
ram[52615] = {-9'd23,-10'd224};
ram[52616] = {-9'd20,-10'd220};
ram[52617] = {-9'd17,-10'd217};
ram[52618] = {-9'd14,-10'd214};
ram[52619] = {-9'd11,-10'd211};
ram[52620] = {-9'd8,-10'd208};
ram[52621] = {-9'd4,-10'd205};
ram[52622] = {-9'd1,-10'd202};
ram[52623] = {9'd2,-10'd198};
ram[52624] = {9'd5,-10'd195};
ram[52625] = {9'd8,-10'd192};
ram[52626] = {9'd11,-10'd189};
ram[52627] = {9'd14,-10'd186};
ram[52628] = {9'd18,-10'd183};
ram[52629] = {9'd21,-10'd180};
ram[52630] = {9'd24,-10'd176};
ram[52631] = {9'd27,-10'd173};
ram[52632] = {9'd30,-10'd170};
ram[52633] = {9'd33,-10'd167};
ram[52634] = {9'd36,-10'd164};
ram[52635] = {9'd40,-10'd161};
ram[52636] = {9'd43,-10'd158};
ram[52637] = {9'd46,-10'd154};
ram[52638] = {9'd49,-10'd151};
ram[52639] = {9'd52,-10'd148};
ram[52640] = {9'd55,-10'd145};
ram[52641] = {9'd58,-10'd142};
ram[52642] = {9'd62,-10'd139};
ram[52643] = {9'd65,-10'd136};
ram[52644] = {9'd68,-10'd132};
ram[52645] = {9'd71,-10'd129};
ram[52646] = {9'd74,-10'd126};
ram[52647] = {9'd77,-10'd123};
ram[52648] = {9'd80,-10'd120};
ram[52649] = {9'd84,-10'd117};
ram[52650] = {9'd87,-10'd114};
ram[52651] = {9'd90,-10'd110};
ram[52652] = {9'd93,-10'd107};
ram[52653] = {9'd96,-10'd104};
ram[52654] = {9'd99,-10'd101};
ram[52655] = {-9'd98,-10'd98};
ram[52656] = {-9'd95,-10'd95};
ram[52657] = {-9'd92,-10'd92};
ram[52658] = {-9'd88,-10'd88};
ram[52659] = {-9'd85,-10'd85};
ram[52660] = {-9'd82,-10'd82};
ram[52661] = {-9'd79,-10'd79};
ram[52662] = {-9'd76,-10'd76};
ram[52663] = {-9'd73,-10'd73};
ram[52664] = {-9'd70,-10'd70};
ram[52665] = {-9'd66,-10'd66};
ram[52666] = {-9'd63,-10'd63};
ram[52667] = {-9'd60,-10'd60};
ram[52668] = {-9'd57,-10'd57};
ram[52669] = {-9'd54,-10'd54};
ram[52670] = {-9'd51,-10'd51};
ram[52671] = {-9'd48,-10'd48};
ram[52672] = {-9'd44,-10'd44};
ram[52673] = {-9'd41,-10'd41};
ram[52674] = {-9'd38,-10'd38};
ram[52675] = {-9'd35,-10'd35};
ram[52676] = {-9'd32,-10'd32};
ram[52677] = {-9'd29,-10'd29};
ram[52678] = {-9'd26,-10'd26};
ram[52679] = {-9'd22,-10'd22};
ram[52680] = {-9'd19,-10'd19};
ram[52681] = {-9'd16,-10'd16};
ram[52682] = {-9'd13,-10'd13};
ram[52683] = {-9'd10,-10'd10};
ram[52684] = {-9'd7,-10'd7};
ram[52685] = {-9'd4,-10'd4};
ram[52686] = {9'd0,10'd0};
ram[52687] = {9'd3,10'd3};
ram[52688] = {9'd6,10'd6};
ram[52689] = {9'd9,10'd9};
ram[52690] = {9'd12,10'd12};
ram[52691] = {9'd15,10'd15};
ram[52692] = {9'd18,10'd18};
ram[52693] = {9'd21,10'd21};
ram[52694] = {9'd25,10'd25};
ram[52695] = {9'd28,10'd28};
ram[52696] = {9'd31,10'd31};
ram[52697] = {9'd34,10'd34};
ram[52698] = {9'd37,10'd37};
ram[52699] = {9'd40,10'd40};
ram[52700] = {9'd43,10'd43};
ram[52701] = {9'd47,10'd47};
ram[52702] = {9'd50,10'd50};
ram[52703] = {9'd53,10'd53};
ram[52704] = {9'd56,10'd56};
ram[52705] = {9'd59,10'd59};
ram[52706] = {9'd62,10'd62};
ram[52707] = {9'd65,10'd65};
ram[52708] = {9'd69,10'd69};
ram[52709] = {9'd72,10'd72};
ram[52710] = {9'd75,10'd75};
ram[52711] = {9'd78,10'd78};
ram[52712] = {9'd81,10'd81};
ram[52713] = {9'd84,10'd84};
ram[52714] = {9'd87,10'd87};
ram[52715] = {9'd91,10'd91};
ram[52716] = {9'd94,10'd94};
ram[52717] = {9'd97,10'd97};
ram[52718] = {-9'd100,10'd100};
ram[52719] = {-9'd97,10'd103};
ram[52720] = {-9'd94,10'd106};
ram[52721] = {-9'd91,10'd109};
ram[52722] = {-9'd88,10'd113};
ram[52723] = {-9'd85,10'd116};
ram[52724] = {-9'd81,10'd119};
ram[52725] = {-9'd78,10'd122};
ram[52726] = {-9'd75,10'd125};
ram[52727] = {-9'd72,10'd128};
ram[52728] = {-9'd69,10'd131};
ram[52729] = {-9'd66,10'd135};
ram[52730] = {-9'd63,10'd138};
ram[52731] = {-9'd59,10'd141};
ram[52732] = {-9'd56,10'd144};
ram[52733] = {-9'd53,10'd147};
ram[52734] = {-9'd50,10'd150};
ram[52735] = {-9'd47,10'd153};
ram[52736] = {-9'd47,10'd153};
ram[52737] = {-9'd44,10'd157};
ram[52738] = {-9'd41,10'd160};
ram[52739] = {-9'd37,10'd163};
ram[52740] = {-9'd34,10'd166};
ram[52741] = {-9'd31,10'd169};
ram[52742] = {-9'd28,10'd172};
ram[52743] = {-9'd25,10'd175};
ram[52744] = {-9'd22,10'd179};
ram[52745] = {-9'd19,10'd182};
ram[52746] = {-9'd15,10'd185};
ram[52747] = {-9'd12,10'd188};
ram[52748] = {-9'd9,10'd191};
ram[52749] = {-9'd6,10'd194};
ram[52750] = {-9'd3,10'd197};
ram[52751] = {9'd0,10'd201};
ram[52752] = {9'd3,10'd204};
ram[52753] = {9'd7,10'd207};
ram[52754] = {9'd10,10'd210};
ram[52755] = {9'd13,10'd213};
ram[52756] = {9'd16,10'd216};
ram[52757] = {9'd19,10'd219};
ram[52758] = {9'd22,10'd223};
ram[52759] = {9'd25,10'd226};
ram[52760] = {9'd29,10'd229};
ram[52761] = {9'd32,10'd232};
ram[52762] = {9'd35,10'd235};
ram[52763] = {9'd38,10'd238};
ram[52764] = {9'd41,10'd241};
ram[52765] = {9'd44,10'd245};
ram[52766] = {9'd47,10'd248};
ram[52767] = {9'd51,10'd251};
ram[52768] = {9'd54,10'd254};
ram[52769] = {9'd57,10'd257};
ram[52770] = {9'd60,10'd260};
ram[52771] = {9'd63,10'd263};
ram[52772] = {9'd66,10'd267};
ram[52773] = {9'd69,10'd270};
ram[52774] = {9'd73,10'd273};
ram[52775] = {9'd76,10'd276};
ram[52776] = {9'd79,10'd279};
ram[52777] = {9'd82,10'd282};
ram[52778] = {9'd85,10'd285};
ram[52779] = {9'd88,10'd289};
ram[52780] = {9'd91,10'd292};
ram[52781] = {9'd95,10'd295};
ram[52782] = {9'd98,10'd298};
ram[52783] = {-9'd99,10'd301};
ram[52784] = {-9'd96,10'd304};
ram[52785] = {-9'd93,10'd307};
ram[52786] = {-9'd90,10'd311};
ram[52787] = {-9'd87,10'd314};
ram[52788] = {-9'd84,10'd317};
ram[52789] = {-9'd81,10'd320};
ram[52790] = {-9'd77,10'd323};
ram[52791] = {-9'd74,10'd326};
ram[52792] = {-9'd71,10'd329};
ram[52793] = {-9'd68,10'd333};
ram[52794] = {-9'd65,10'd336};
ram[52795] = {-9'd62,10'd339};
ram[52796] = {-9'd59,10'd342};
ram[52797] = {-9'd55,10'd345};
ram[52798] = {-9'd52,10'd348};
ram[52799] = {-9'd49,10'd351};
ram[52800] = {-9'd46,10'd354};
ram[52801] = {-9'd43,10'd358};
ram[52802] = {-9'd40,10'd361};
ram[52803] = {-9'd37,10'd364};
ram[52804] = {-9'd33,10'd367};
ram[52805] = {-9'd30,10'd370};
ram[52806] = {-9'd27,10'd373};
ram[52807] = {-9'd24,10'd376};
ram[52808] = {-9'd21,10'd380};
ram[52809] = {-9'd18,10'd383};
ram[52810] = {-9'd15,10'd386};
ram[52811] = {-9'd11,10'd389};
ram[52812] = {-9'd8,10'd392};
ram[52813] = {-9'd5,10'd395};
ram[52814] = {-9'd2,10'd398};
ram[52815] = {9'd1,-10'd399};
ram[52816] = {9'd4,-10'd396};
ram[52817] = {9'd7,-10'd393};
ram[52818] = {9'd10,-10'd390};
ram[52819] = {9'd14,-10'd387};
ram[52820] = {9'd17,-10'd384};
ram[52821] = {9'd20,-10'd381};
ram[52822] = {9'd23,-10'd377};
ram[52823] = {9'd26,-10'd374};
ram[52824] = {9'd29,-10'd371};
ram[52825] = {9'd32,-10'd368};
ram[52826] = {9'd36,-10'd365};
ram[52827] = {9'd39,-10'd362};
ram[52828] = {9'd42,-10'd359};
ram[52829] = {9'd45,-10'd355};
ram[52830] = {9'd48,-10'd352};
ram[52831] = {9'd51,-10'd349};
ram[52832] = {9'd54,-10'd346};
ram[52833] = {9'd58,-10'd343};
ram[52834] = {9'd61,-10'd340};
ram[52835] = {9'd64,-10'd337};
ram[52836] = {9'd67,-10'd334};
ram[52837] = {9'd70,-10'd330};
ram[52838] = {9'd73,-10'd327};
ram[52839] = {9'd76,-10'd324};
ram[52840] = {9'd80,-10'd321};
ram[52841] = {9'd83,-10'd318};
ram[52842] = {9'd86,-10'd315};
ram[52843] = {9'd89,-10'd312};
ram[52844] = {9'd92,-10'd308};
ram[52845] = {9'd95,-10'd305};
ram[52846] = {9'd98,-10'd302};
ram[52847] = {-9'd99,-10'd299};
ram[52848] = {-9'd96,-10'd296};
ram[52849] = {-9'd92,-10'd293};
ram[52850] = {-9'd89,-10'd290};
ram[52851] = {-9'd86,-10'd286};
ram[52852] = {-9'd83,-10'd283};
ram[52853] = {-9'd80,-10'd280};
ram[52854] = {-9'd77,-10'd277};
ram[52855] = {-9'd74,-10'd274};
ram[52856] = {-9'd70,-10'd271};
ram[52857] = {-9'd67,-10'd268};
ram[52858] = {-9'd64,-10'd264};
ram[52859] = {-9'd61,-10'd261};
ram[52860] = {-9'd58,-10'd258};
ram[52861] = {-9'd55,-10'd255};
ram[52862] = {-9'd52,-10'd252};
ram[52863] = {-9'd48,-10'd249};
ram[52864] = {-9'd48,-10'd249};
ram[52865] = {-9'd45,-10'd246};
ram[52866] = {-9'd42,-10'd242};
ram[52867] = {-9'd39,-10'd239};
ram[52868] = {-9'd36,-10'd236};
ram[52869] = {-9'd33,-10'd233};
ram[52870] = {-9'd30,-10'd230};
ram[52871] = {-9'd26,-10'd227};
ram[52872] = {-9'd23,-10'd224};
ram[52873] = {-9'd20,-10'd220};
ram[52874] = {-9'd17,-10'd217};
ram[52875] = {-9'd14,-10'd214};
ram[52876] = {-9'd11,-10'd211};
ram[52877] = {-9'd8,-10'd208};
ram[52878] = {-9'd4,-10'd205};
ram[52879] = {-9'd1,-10'd202};
ram[52880] = {9'd2,-10'd198};
ram[52881] = {9'd5,-10'd195};
ram[52882] = {9'd8,-10'd192};
ram[52883] = {9'd11,-10'd189};
ram[52884] = {9'd14,-10'd186};
ram[52885] = {9'd18,-10'd183};
ram[52886] = {9'd21,-10'd180};
ram[52887] = {9'd24,-10'd176};
ram[52888] = {9'd27,-10'd173};
ram[52889] = {9'd30,-10'd170};
ram[52890] = {9'd33,-10'd167};
ram[52891] = {9'd36,-10'd164};
ram[52892] = {9'd40,-10'd161};
ram[52893] = {9'd43,-10'd158};
ram[52894] = {9'd46,-10'd154};
ram[52895] = {9'd49,-10'd151};
ram[52896] = {9'd52,-10'd148};
ram[52897] = {9'd55,-10'd145};
ram[52898] = {9'd58,-10'd142};
ram[52899] = {9'd62,-10'd139};
ram[52900] = {9'd65,-10'd136};
ram[52901] = {9'd68,-10'd132};
ram[52902] = {9'd71,-10'd129};
ram[52903] = {9'd74,-10'd126};
ram[52904] = {9'd77,-10'd123};
ram[52905] = {9'd80,-10'd120};
ram[52906] = {9'd84,-10'd117};
ram[52907] = {9'd87,-10'd114};
ram[52908] = {9'd90,-10'd110};
ram[52909] = {9'd93,-10'd107};
ram[52910] = {9'd96,-10'd104};
ram[52911] = {9'd99,-10'd101};
ram[52912] = {-9'd98,-10'd98};
ram[52913] = {-9'd95,-10'd95};
ram[52914] = {-9'd92,-10'd92};
ram[52915] = {-9'd88,-10'd88};
ram[52916] = {-9'd85,-10'd85};
ram[52917] = {-9'd82,-10'd82};
ram[52918] = {-9'd79,-10'd79};
ram[52919] = {-9'd76,-10'd76};
ram[52920] = {-9'd73,-10'd73};
ram[52921] = {-9'd70,-10'd70};
ram[52922] = {-9'd66,-10'd66};
ram[52923] = {-9'd63,-10'd63};
ram[52924] = {-9'd60,-10'd60};
ram[52925] = {-9'd57,-10'd57};
ram[52926] = {-9'd54,-10'd54};
ram[52927] = {-9'd51,-10'd51};
ram[52928] = {-9'd48,-10'd48};
ram[52929] = {-9'd44,-10'd44};
ram[52930] = {-9'd41,-10'd41};
ram[52931] = {-9'd38,-10'd38};
ram[52932] = {-9'd35,-10'd35};
ram[52933] = {-9'd32,-10'd32};
ram[52934] = {-9'd29,-10'd29};
ram[52935] = {-9'd26,-10'd26};
ram[52936] = {-9'd22,-10'd22};
ram[52937] = {-9'd19,-10'd19};
ram[52938] = {-9'd16,-10'd16};
ram[52939] = {-9'd13,-10'd13};
ram[52940] = {-9'd10,-10'd10};
ram[52941] = {-9'd7,-10'd7};
ram[52942] = {-9'd4,-10'd4};
ram[52943] = {9'd0,10'd0};
ram[52944] = {9'd3,10'd3};
ram[52945] = {9'd6,10'd6};
ram[52946] = {9'd9,10'd9};
ram[52947] = {9'd12,10'd12};
ram[52948] = {9'd15,10'd15};
ram[52949] = {9'd18,10'd18};
ram[52950] = {9'd21,10'd21};
ram[52951] = {9'd25,10'd25};
ram[52952] = {9'd28,10'd28};
ram[52953] = {9'd31,10'd31};
ram[52954] = {9'd34,10'd34};
ram[52955] = {9'd37,10'd37};
ram[52956] = {9'd40,10'd40};
ram[52957] = {9'd43,10'd43};
ram[52958] = {9'd47,10'd47};
ram[52959] = {9'd50,10'd50};
ram[52960] = {9'd53,10'd53};
ram[52961] = {9'd56,10'd56};
ram[52962] = {9'd59,10'd59};
ram[52963] = {9'd62,10'd62};
ram[52964] = {9'd65,10'd65};
ram[52965] = {9'd69,10'd69};
ram[52966] = {9'd72,10'd72};
ram[52967] = {9'd75,10'd75};
ram[52968] = {9'd78,10'd78};
ram[52969] = {9'd81,10'd81};
ram[52970] = {9'd84,10'd84};
ram[52971] = {9'd87,10'd87};
ram[52972] = {9'd91,10'd91};
ram[52973] = {9'd94,10'd94};
ram[52974] = {9'd97,10'd97};
ram[52975] = {-9'd100,10'd100};
ram[52976] = {-9'd97,10'd103};
ram[52977] = {-9'd94,10'd106};
ram[52978] = {-9'd91,10'd109};
ram[52979] = {-9'd88,10'd113};
ram[52980] = {-9'd85,10'd116};
ram[52981] = {-9'd81,10'd119};
ram[52982] = {-9'd78,10'd122};
ram[52983] = {-9'd75,10'd125};
ram[52984] = {-9'd72,10'd128};
ram[52985] = {-9'd69,10'd131};
ram[52986] = {-9'd66,10'd135};
ram[52987] = {-9'd63,10'd138};
ram[52988] = {-9'd59,10'd141};
ram[52989] = {-9'd56,10'd144};
ram[52990] = {-9'd53,10'd147};
ram[52991] = {-9'd50,10'd150};
ram[52992] = {-9'd50,10'd150};
ram[52993] = {-9'd47,10'd153};
ram[52994] = {-9'd44,10'd157};
ram[52995] = {-9'd41,10'd160};
ram[52996] = {-9'd37,10'd163};
ram[52997] = {-9'd34,10'd166};
ram[52998] = {-9'd31,10'd169};
ram[52999] = {-9'd28,10'd172};
ram[53000] = {-9'd25,10'd175};
ram[53001] = {-9'd22,10'd179};
ram[53002] = {-9'd19,10'd182};
ram[53003] = {-9'd15,10'd185};
ram[53004] = {-9'd12,10'd188};
ram[53005] = {-9'd9,10'd191};
ram[53006] = {-9'd6,10'd194};
ram[53007] = {-9'd3,10'd197};
ram[53008] = {9'd0,10'd201};
ram[53009] = {9'd3,10'd204};
ram[53010] = {9'd7,10'd207};
ram[53011] = {9'd10,10'd210};
ram[53012] = {9'd13,10'd213};
ram[53013] = {9'd16,10'd216};
ram[53014] = {9'd19,10'd219};
ram[53015] = {9'd22,10'd223};
ram[53016] = {9'd25,10'd226};
ram[53017] = {9'd29,10'd229};
ram[53018] = {9'd32,10'd232};
ram[53019] = {9'd35,10'd235};
ram[53020] = {9'd38,10'd238};
ram[53021] = {9'd41,10'd241};
ram[53022] = {9'd44,10'd245};
ram[53023] = {9'd47,10'd248};
ram[53024] = {9'd51,10'd251};
ram[53025] = {9'd54,10'd254};
ram[53026] = {9'd57,10'd257};
ram[53027] = {9'd60,10'd260};
ram[53028] = {9'd63,10'd263};
ram[53029] = {9'd66,10'd267};
ram[53030] = {9'd69,10'd270};
ram[53031] = {9'd73,10'd273};
ram[53032] = {9'd76,10'd276};
ram[53033] = {9'd79,10'd279};
ram[53034] = {9'd82,10'd282};
ram[53035] = {9'd85,10'd285};
ram[53036] = {9'd88,10'd289};
ram[53037] = {9'd91,10'd292};
ram[53038] = {9'd95,10'd295};
ram[53039] = {9'd98,10'd298};
ram[53040] = {-9'd99,10'd301};
ram[53041] = {-9'd96,10'd304};
ram[53042] = {-9'd93,10'd307};
ram[53043] = {-9'd90,10'd311};
ram[53044] = {-9'd87,10'd314};
ram[53045] = {-9'd84,10'd317};
ram[53046] = {-9'd81,10'd320};
ram[53047] = {-9'd77,10'd323};
ram[53048] = {-9'd74,10'd326};
ram[53049] = {-9'd71,10'd329};
ram[53050] = {-9'd68,10'd333};
ram[53051] = {-9'd65,10'd336};
ram[53052] = {-9'd62,10'd339};
ram[53053] = {-9'd59,10'd342};
ram[53054] = {-9'd55,10'd345};
ram[53055] = {-9'd52,10'd348};
ram[53056] = {-9'd49,10'd351};
ram[53057] = {-9'd46,10'd354};
ram[53058] = {-9'd43,10'd358};
ram[53059] = {-9'd40,10'd361};
ram[53060] = {-9'd37,10'd364};
ram[53061] = {-9'd33,10'd367};
ram[53062] = {-9'd30,10'd370};
ram[53063] = {-9'd27,10'd373};
ram[53064] = {-9'd24,10'd376};
ram[53065] = {-9'd21,10'd380};
ram[53066] = {-9'd18,10'd383};
ram[53067] = {-9'd15,10'd386};
ram[53068] = {-9'd11,10'd389};
ram[53069] = {-9'd8,10'd392};
ram[53070] = {-9'd5,10'd395};
ram[53071] = {-9'd2,10'd398};
ram[53072] = {9'd1,-10'd399};
ram[53073] = {9'd4,-10'd396};
ram[53074] = {9'd7,-10'd393};
ram[53075] = {9'd10,-10'd390};
ram[53076] = {9'd14,-10'd387};
ram[53077] = {9'd17,-10'd384};
ram[53078] = {9'd20,-10'd381};
ram[53079] = {9'd23,-10'd377};
ram[53080] = {9'd26,-10'd374};
ram[53081] = {9'd29,-10'd371};
ram[53082] = {9'd32,-10'd368};
ram[53083] = {9'd36,-10'd365};
ram[53084] = {9'd39,-10'd362};
ram[53085] = {9'd42,-10'd359};
ram[53086] = {9'd45,-10'd355};
ram[53087] = {9'd48,-10'd352};
ram[53088] = {9'd51,-10'd349};
ram[53089] = {9'd54,-10'd346};
ram[53090] = {9'd58,-10'd343};
ram[53091] = {9'd61,-10'd340};
ram[53092] = {9'd64,-10'd337};
ram[53093] = {9'd67,-10'd334};
ram[53094] = {9'd70,-10'd330};
ram[53095] = {9'd73,-10'd327};
ram[53096] = {9'd76,-10'd324};
ram[53097] = {9'd80,-10'd321};
ram[53098] = {9'd83,-10'd318};
ram[53099] = {9'd86,-10'd315};
ram[53100] = {9'd89,-10'd312};
ram[53101] = {9'd92,-10'd308};
ram[53102] = {9'd95,-10'd305};
ram[53103] = {9'd98,-10'd302};
ram[53104] = {-9'd99,-10'd299};
ram[53105] = {-9'd96,-10'd296};
ram[53106] = {-9'd92,-10'd293};
ram[53107] = {-9'd89,-10'd290};
ram[53108] = {-9'd86,-10'd286};
ram[53109] = {-9'd83,-10'd283};
ram[53110] = {-9'd80,-10'd280};
ram[53111] = {-9'd77,-10'd277};
ram[53112] = {-9'd74,-10'd274};
ram[53113] = {-9'd70,-10'd271};
ram[53114] = {-9'd67,-10'd268};
ram[53115] = {-9'd64,-10'd264};
ram[53116] = {-9'd61,-10'd261};
ram[53117] = {-9'd58,-10'd258};
ram[53118] = {-9'd55,-10'd255};
ram[53119] = {-9'd52,-10'd252};
ram[53120] = {-9'd52,-10'd252};
ram[53121] = {-9'd48,-10'd249};
ram[53122] = {-9'd45,-10'd246};
ram[53123] = {-9'd42,-10'd242};
ram[53124] = {-9'd39,-10'd239};
ram[53125] = {-9'd36,-10'd236};
ram[53126] = {-9'd33,-10'd233};
ram[53127] = {-9'd30,-10'd230};
ram[53128] = {-9'd26,-10'd227};
ram[53129] = {-9'd23,-10'd224};
ram[53130] = {-9'd20,-10'd220};
ram[53131] = {-9'd17,-10'd217};
ram[53132] = {-9'd14,-10'd214};
ram[53133] = {-9'd11,-10'd211};
ram[53134] = {-9'd8,-10'd208};
ram[53135] = {-9'd4,-10'd205};
ram[53136] = {-9'd1,-10'd202};
ram[53137] = {9'd2,-10'd198};
ram[53138] = {9'd5,-10'd195};
ram[53139] = {9'd8,-10'd192};
ram[53140] = {9'd11,-10'd189};
ram[53141] = {9'd14,-10'd186};
ram[53142] = {9'd18,-10'd183};
ram[53143] = {9'd21,-10'd180};
ram[53144] = {9'd24,-10'd176};
ram[53145] = {9'd27,-10'd173};
ram[53146] = {9'd30,-10'd170};
ram[53147] = {9'd33,-10'd167};
ram[53148] = {9'd36,-10'd164};
ram[53149] = {9'd40,-10'd161};
ram[53150] = {9'd43,-10'd158};
ram[53151] = {9'd46,-10'd154};
ram[53152] = {9'd49,-10'd151};
ram[53153] = {9'd52,-10'd148};
ram[53154] = {9'd55,-10'd145};
ram[53155] = {9'd58,-10'd142};
ram[53156] = {9'd62,-10'd139};
ram[53157] = {9'd65,-10'd136};
ram[53158] = {9'd68,-10'd132};
ram[53159] = {9'd71,-10'd129};
ram[53160] = {9'd74,-10'd126};
ram[53161] = {9'd77,-10'd123};
ram[53162] = {9'd80,-10'd120};
ram[53163] = {9'd84,-10'd117};
ram[53164] = {9'd87,-10'd114};
ram[53165] = {9'd90,-10'd110};
ram[53166] = {9'd93,-10'd107};
ram[53167] = {9'd96,-10'd104};
ram[53168] = {9'd99,-10'd101};
ram[53169] = {-9'd98,-10'd98};
ram[53170] = {-9'd95,-10'd95};
ram[53171] = {-9'd92,-10'd92};
ram[53172] = {-9'd88,-10'd88};
ram[53173] = {-9'd85,-10'd85};
ram[53174] = {-9'd82,-10'd82};
ram[53175] = {-9'd79,-10'd79};
ram[53176] = {-9'd76,-10'd76};
ram[53177] = {-9'd73,-10'd73};
ram[53178] = {-9'd70,-10'd70};
ram[53179] = {-9'd66,-10'd66};
ram[53180] = {-9'd63,-10'd63};
ram[53181] = {-9'd60,-10'd60};
ram[53182] = {-9'd57,-10'd57};
ram[53183] = {-9'd54,-10'd54};
ram[53184] = {-9'd51,-10'd51};
ram[53185] = {-9'd48,-10'd48};
ram[53186] = {-9'd44,-10'd44};
ram[53187] = {-9'd41,-10'd41};
ram[53188] = {-9'd38,-10'd38};
ram[53189] = {-9'd35,-10'd35};
ram[53190] = {-9'd32,-10'd32};
ram[53191] = {-9'd29,-10'd29};
ram[53192] = {-9'd26,-10'd26};
ram[53193] = {-9'd22,-10'd22};
ram[53194] = {-9'd19,-10'd19};
ram[53195] = {-9'd16,-10'd16};
ram[53196] = {-9'd13,-10'd13};
ram[53197] = {-9'd10,-10'd10};
ram[53198] = {-9'd7,-10'd7};
ram[53199] = {-9'd4,-10'd4};
ram[53200] = {9'd0,10'd0};
ram[53201] = {9'd3,10'd3};
ram[53202] = {9'd6,10'd6};
ram[53203] = {9'd9,10'd9};
ram[53204] = {9'd12,10'd12};
ram[53205] = {9'd15,10'd15};
ram[53206] = {9'd18,10'd18};
ram[53207] = {9'd21,10'd21};
ram[53208] = {9'd25,10'd25};
ram[53209] = {9'd28,10'd28};
ram[53210] = {9'd31,10'd31};
ram[53211] = {9'd34,10'd34};
ram[53212] = {9'd37,10'd37};
ram[53213] = {9'd40,10'd40};
ram[53214] = {9'd43,10'd43};
ram[53215] = {9'd47,10'd47};
ram[53216] = {9'd50,10'd50};
ram[53217] = {9'd53,10'd53};
ram[53218] = {9'd56,10'd56};
ram[53219] = {9'd59,10'd59};
ram[53220] = {9'd62,10'd62};
ram[53221] = {9'd65,10'd65};
ram[53222] = {9'd69,10'd69};
ram[53223] = {9'd72,10'd72};
ram[53224] = {9'd75,10'd75};
ram[53225] = {9'd78,10'd78};
ram[53226] = {9'd81,10'd81};
ram[53227] = {9'd84,10'd84};
ram[53228] = {9'd87,10'd87};
ram[53229] = {9'd91,10'd91};
ram[53230] = {9'd94,10'd94};
ram[53231] = {9'd97,10'd97};
ram[53232] = {-9'd100,10'd100};
ram[53233] = {-9'd97,10'd103};
ram[53234] = {-9'd94,10'd106};
ram[53235] = {-9'd91,10'd109};
ram[53236] = {-9'd88,10'd113};
ram[53237] = {-9'd85,10'd116};
ram[53238] = {-9'd81,10'd119};
ram[53239] = {-9'd78,10'd122};
ram[53240] = {-9'd75,10'd125};
ram[53241] = {-9'd72,10'd128};
ram[53242] = {-9'd69,10'd131};
ram[53243] = {-9'd66,10'd135};
ram[53244] = {-9'd63,10'd138};
ram[53245] = {-9'd59,10'd141};
ram[53246] = {-9'd56,10'd144};
ram[53247] = {-9'd53,10'd147};
ram[53248] = {-9'd53,10'd147};
ram[53249] = {-9'd50,10'd150};
ram[53250] = {-9'd47,10'd153};
ram[53251] = {-9'd44,10'd157};
ram[53252] = {-9'd41,10'd160};
ram[53253] = {-9'd37,10'd163};
ram[53254] = {-9'd34,10'd166};
ram[53255] = {-9'd31,10'd169};
ram[53256] = {-9'd28,10'd172};
ram[53257] = {-9'd25,10'd175};
ram[53258] = {-9'd22,10'd179};
ram[53259] = {-9'd19,10'd182};
ram[53260] = {-9'd15,10'd185};
ram[53261] = {-9'd12,10'd188};
ram[53262] = {-9'd9,10'd191};
ram[53263] = {-9'd6,10'd194};
ram[53264] = {-9'd3,10'd197};
ram[53265] = {9'd0,10'd201};
ram[53266] = {9'd3,10'd204};
ram[53267] = {9'd7,10'd207};
ram[53268] = {9'd10,10'd210};
ram[53269] = {9'd13,10'd213};
ram[53270] = {9'd16,10'd216};
ram[53271] = {9'd19,10'd219};
ram[53272] = {9'd22,10'd223};
ram[53273] = {9'd25,10'd226};
ram[53274] = {9'd29,10'd229};
ram[53275] = {9'd32,10'd232};
ram[53276] = {9'd35,10'd235};
ram[53277] = {9'd38,10'd238};
ram[53278] = {9'd41,10'd241};
ram[53279] = {9'd44,10'd245};
ram[53280] = {9'd47,10'd248};
ram[53281] = {9'd51,10'd251};
ram[53282] = {9'd54,10'd254};
ram[53283] = {9'd57,10'd257};
ram[53284] = {9'd60,10'd260};
ram[53285] = {9'd63,10'd263};
ram[53286] = {9'd66,10'd267};
ram[53287] = {9'd69,10'd270};
ram[53288] = {9'd73,10'd273};
ram[53289] = {9'd76,10'd276};
ram[53290] = {9'd79,10'd279};
ram[53291] = {9'd82,10'd282};
ram[53292] = {9'd85,10'd285};
ram[53293] = {9'd88,10'd289};
ram[53294] = {9'd91,10'd292};
ram[53295] = {9'd95,10'd295};
ram[53296] = {9'd98,10'd298};
ram[53297] = {-9'd99,10'd301};
ram[53298] = {-9'd96,10'd304};
ram[53299] = {-9'd93,10'd307};
ram[53300] = {-9'd90,10'd311};
ram[53301] = {-9'd87,10'd314};
ram[53302] = {-9'd84,10'd317};
ram[53303] = {-9'd81,10'd320};
ram[53304] = {-9'd77,10'd323};
ram[53305] = {-9'd74,10'd326};
ram[53306] = {-9'd71,10'd329};
ram[53307] = {-9'd68,10'd333};
ram[53308] = {-9'd65,10'd336};
ram[53309] = {-9'd62,10'd339};
ram[53310] = {-9'd59,10'd342};
ram[53311] = {-9'd55,10'd345};
ram[53312] = {-9'd52,10'd348};
ram[53313] = {-9'd49,10'd351};
ram[53314] = {-9'd46,10'd354};
ram[53315] = {-9'd43,10'd358};
ram[53316] = {-9'd40,10'd361};
ram[53317] = {-9'd37,10'd364};
ram[53318] = {-9'd33,10'd367};
ram[53319] = {-9'd30,10'd370};
ram[53320] = {-9'd27,10'd373};
ram[53321] = {-9'd24,10'd376};
ram[53322] = {-9'd21,10'd380};
ram[53323] = {-9'd18,10'd383};
ram[53324] = {-9'd15,10'd386};
ram[53325] = {-9'd11,10'd389};
ram[53326] = {-9'd8,10'd392};
ram[53327] = {-9'd5,10'd395};
ram[53328] = {-9'd2,10'd398};
ram[53329] = {9'd1,-10'd399};
ram[53330] = {9'd4,-10'd396};
ram[53331] = {9'd7,-10'd393};
ram[53332] = {9'd10,-10'd390};
ram[53333] = {9'd14,-10'd387};
ram[53334] = {9'd17,-10'd384};
ram[53335] = {9'd20,-10'd381};
ram[53336] = {9'd23,-10'd377};
ram[53337] = {9'd26,-10'd374};
ram[53338] = {9'd29,-10'd371};
ram[53339] = {9'd32,-10'd368};
ram[53340] = {9'd36,-10'd365};
ram[53341] = {9'd39,-10'd362};
ram[53342] = {9'd42,-10'd359};
ram[53343] = {9'd45,-10'd355};
ram[53344] = {9'd48,-10'd352};
ram[53345] = {9'd51,-10'd349};
ram[53346] = {9'd54,-10'd346};
ram[53347] = {9'd58,-10'd343};
ram[53348] = {9'd61,-10'd340};
ram[53349] = {9'd64,-10'd337};
ram[53350] = {9'd67,-10'd334};
ram[53351] = {9'd70,-10'd330};
ram[53352] = {9'd73,-10'd327};
ram[53353] = {9'd76,-10'd324};
ram[53354] = {9'd80,-10'd321};
ram[53355] = {9'd83,-10'd318};
ram[53356] = {9'd86,-10'd315};
ram[53357] = {9'd89,-10'd312};
ram[53358] = {9'd92,-10'd308};
ram[53359] = {9'd95,-10'd305};
ram[53360] = {9'd98,-10'd302};
ram[53361] = {-9'd99,-10'd299};
ram[53362] = {-9'd96,-10'd296};
ram[53363] = {-9'd92,-10'd293};
ram[53364] = {-9'd89,-10'd290};
ram[53365] = {-9'd86,-10'd286};
ram[53366] = {-9'd83,-10'd283};
ram[53367] = {-9'd80,-10'd280};
ram[53368] = {-9'd77,-10'd277};
ram[53369] = {-9'd74,-10'd274};
ram[53370] = {-9'd70,-10'd271};
ram[53371] = {-9'd67,-10'd268};
ram[53372] = {-9'd64,-10'd264};
ram[53373] = {-9'd61,-10'd261};
ram[53374] = {-9'd58,-10'd258};
ram[53375] = {-9'd55,-10'd255};
ram[53376] = {-9'd55,-10'd255};
ram[53377] = {-9'd52,-10'd252};
ram[53378] = {-9'd48,-10'd249};
ram[53379] = {-9'd45,-10'd246};
ram[53380] = {-9'd42,-10'd242};
ram[53381] = {-9'd39,-10'd239};
ram[53382] = {-9'd36,-10'd236};
ram[53383] = {-9'd33,-10'd233};
ram[53384] = {-9'd30,-10'd230};
ram[53385] = {-9'd26,-10'd227};
ram[53386] = {-9'd23,-10'd224};
ram[53387] = {-9'd20,-10'd220};
ram[53388] = {-9'd17,-10'd217};
ram[53389] = {-9'd14,-10'd214};
ram[53390] = {-9'd11,-10'd211};
ram[53391] = {-9'd8,-10'd208};
ram[53392] = {-9'd4,-10'd205};
ram[53393] = {-9'd1,-10'd202};
ram[53394] = {9'd2,-10'd198};
ram[53395] = {9'd5,-10'd195};
ram[53396] = {9'd8,-10'd192};
ram[53397] = {9'd11,-10'd189};
ram[53398] = {9'd14,-10'd186};
ram[53399] = {9'd18,-10'd183};
ram[53400] = {9'd21,-10'd180};
ram[53401] = {9'd24,-10'd176};
ram[53402] = {9'd27,-10'd173};
ram[53403] = {9'd30,-10'd170};
ram[53404] = {9'd33,-10'd167};
ram[53405] = {9'd36,-10'd164};
ram[53406] = {9'd40,-10'd161};
ram[53407] = {9'd43,-10'd158};
ram[53408] = {9'd46,-10'd154};
ram[53409] = {9'd49,-10'd151};
ram[53410] = {9'd52,-10'd148};
ram[53411] = {9'd55,-10'd145};
ram[53412] = {9'd58,-10'd142};
ram[53413] = {9'd62,-10'd139};
ram[53414] = {9'd65,-10'd136};
ram[53415] = {9'd68,-10'd132};
ram[53416] = {9'd71,-10'd129};
ram[53417] = {9'd74,-10'd126};
ram[53418] = {9'd77,-10'd123};
ram[53419] = {9'd80,-10'd120};
ram[53420] = {9'd84,-10'd117};
ram[53421] = {9'd87,-10'd114};
ram[53422] = {9'd90,-10'd110};
ram[53423] = {9'd93,-10'd107};
ram[53424] = {9'd96,-10'd104};
ram[53425] = {9'd99,-10'd101};
ram[53426] = {-9'd98,-10'd98};
ram[53427] = {-9'd95,-10'd95};
ram[53428] = {-9'd92,-10'd92};
ram[53429] = {-9'd88,-10'd88};
ram[53430] = {-9'd85,-10'd85};
ram[53431] = {-9'd82,-10'd82};
ram[53432] = {-9'd79,-10'd79};
ram[53433] = {-9'd76,-10'd76};
ram[53434] = {-9'd73,-10'd73};
ram[53435] = {-9'd70,-10'd70};
ram[53436] = {-9'd66,-10'd66};
ram[53437] = {-9'd63,-10'd63};
ram[53438] = {-9'd60,-10'd60};
ram[53439] = {-9'd57,-10'd57};
ram[53440] = {-9'd54,-10'd54};
ram[53441] = {-9'd51,-10'd51};
ram[53442] = {-9'd48,-10'd48};
ram[53443] = {-9'd44,-10'd44};
ram[53444] = {-9'd41,-10'd41};
ram[53445] = {-9'd38,-10'd38};
ram[53446] = {-9'd35,-10'd35};
ram[53447] = {-9'd32,-10'd32};
ram[53448] = {-9'd29,-10'd29};
ram[53449] = {-9'd26,-10'd26};
ram[53450] = {-9'd22,-10'd22};
ram[53451] = {-9'd19,-10'd19};
ram[53452] = {-9'd16,-10'd16};
ram[53453] = {-9'd13,-10'd13};
ram[53454] = {-9'd10,-10'd10};
ram[53455] = {-9'd7,-10'd7};
ram[53456] = {-9'd4,-10'd4};
ram[53457] = {-9'd1,-10'd1};
ram[53458] = {9'd3,10'd3};
ram[53459] = {9'd6,10'd6};
ram[53460] = {9'd9,10'd9};
ram[53461] = {9'd12,10'd12};
ram[53462] = {9'd15,10'd15};
ram[53463] = {9'd18,10'd18};
ram[53464] = {9'd21,10'd21};
ram[53465] = {9'd25,10'd25};
ram[53466] = {9'd28,10'd28};
ram[53467] = {9'd31,10'd31};
ram[53468] = {9'd34,10'd34};
ram[53469] = {9'd37,10'd37};
ram[53470] = {9'd40,10'd40};
ram[53471] = {9'd43,10'd43};
ram[53472] = {9'd47,10'd47};
ram[53473] = {9'd50,10'd50};
ram[53474] = {9'd53,10'd53};
ram[53475] = {9'd56,10'd56};
ram[53476] = {9'd59,10'd59};
ram[53477] = {9'd62,10'd62};
ram[53478] = {9'd65,10'd65};
ram[53479] = {9'd69,10'd69};
ram[53480] = {9'd72,10'd72};
ram[53481] = {9'd75,10'd75};
ram[53482] = {9'd78,10'd78};
ram[53483] = {9'd81,10'd81};
ram[53484] = {9'd84,10'd84};
ram[53485] = {9'd87,10'd87};
ram[53486] = {9'd91,10'd91};
ram[53487] = {9'd94,10'd94};
ram[53488] = {9'd97,10'd97};
ram[53489] = {-9'd100,10'd100};
ram[53490] = {-9'd97,10'd103};
ram[53491] = {-9'd94,10'd106};
ram[53492] = {-9'd91,10'd109};
ram[53493] = {-9'd88,10'd113};
ram[53494] = {-9'd85,10'd116};
ram[53495] = {-9'd81,10'd119};
ram[53496] = {-9'd78,10'd122};
ram[53497] = {-9'd75,10'd125};
ram[53498] = {-9'd72,10'd128};
ram[53499] = {-9'd69,10'd131};
ram[53500] = {-9'd66,10'd135};
ram[53501] = {-9'd63,10'd138};
ram[53502] = {-9'd59,10'd141};
ram[53503] = {-9'd56,10'd144};
ram[53504] = {-9'd56,10'd144};
ram[53505] = {-9'd53,10'd147};
ram[53506] = {-9'd50,10'd150};
ram[53507] = {-9'd47,10'd153};
ram[53508] = {-9'd44,10'd157};
ram[53509] = {-9'd41,10'd160};
ram[53510] = {-9'd37,10'd163};
ram[53511] = {-9'd34,10'd166};
ram[53512] = {-9'd31,10'd169};
ram[53513] = {-9'd28,10'd172};
ram[53514] = {-9'd25,10'd175};
ram[53515] = {-9'd22,10'd179};
ram[53516] = {-9'd19,10'd182};
ram[53517] = {-9'd15,10'd185};
ram[53518] = {-9'd12,10'd188};
ram[53519] = {-9'd9,10'd191};
ram[53520] = {-9'd6,10'd194};
ram[53521] = {-9'd3,10'd197};
ram[53522] = {9'd0,10'd201};
ram[53523] = {9'd3,10'd204};
ram[53524] = {9'd7,10'd207};
ram[53525] = {9'd10,10'd210};
ram[53526] = {9'd13,10'd213};
ram[53527] = {9'd16,10'd216};
ram[53528] = {9'd19,10'd219};
ram[53529] = {9'd22,10'd223};
ram[53530] = {9'd25,10'd226};
ram[53531] = {9'd29,10'd229};
ram[53532] = {9'd32,10'd232};
ram[53533] = {9'd35,10'd235};
ram[53534] = {9'd38,10'd238};
ram[53535] = {9'd41,10'd241};
ram[53536] = {9'd44,10'd245};
ram[53537] = {9'd47,10'd248};
ram[53538] = {9'd51,10'd251};
ram[53539] = {9'd54,10'd254};
ram[53540] = {9'd57,10'd257};
ram[53541] = {9'd60,10'd260};
ram[53542] = {9'd63,10'd263};
ram[53543] = {9'd66,10'd267};
ram[53544] = {9'd69,10'd270};
ram[53545] = {9'd73,10'd273};
ram[53546] = {9'd76,10'd276};
ram[53547] = {9'd79,10'd279};
ram[53548] = {9'd82,10'd282};
ram[53549] = {9'd85,10'd285};
ram[53550] = {9'd88,10'd289};
ram[53551] = {9'd91,10'd292};
ram[53552] = {9'd95,10'd295};
ram[53553] = {9'd98,10'd298};
ram[53554] = {-9'd99,10'd301};
ram[53555] = {-9'd96,10'd304};
ram[53556] = {-9'd93,10'd307};
ram[53557] = {-9'd90,10'd311};
ram[53558] = {-9'd87,10'd314};
ram[53559] = {-9'd84,10'd317};
ram[53560] = {-9'd81,10'd320};
ram[53561] = {-9'd77,10'd323};
ram[53562] = {-9'd74,10'd326};
ram[53563] = {-9'd71,10'd329};
ram[53564] = {-9'd68,10'd333};
ram[53565] = {-9'd65,10'd336};
ram[53566] = {-9'd62,10'd339};
ram[53567] = {-9'd59,10'd342};
ram[53568] = {-9'd55,10'd345};
ram[53569] = {-9'd52,10'd348};
ram[53570] = {-9'd49,10'd351};
ram[53571] = {-9'd46,10'd354};
ram[53572] = {-9'd43,10'd358};
ram[53573] = {-9'd40,10'd361};
ram[53574] = {-9'd37,10'd364};
ram[53575] = {-9'd33,10'd367};
ram[53576] = {-9'd30,10'd370};
ram[53577] = {-9'd27,10'd373};
ram[53578] = {-9'd24,10'd376};
ram[53579] = {-9'd21,10'd380};
ram[53580] = {-9'd18,10'd383};
ram[53581] = {-9'd15,10'd386};
ram[53582] = {-9'd11,10'd389};
ram[53583] = {-9'd8,10'd392};
ram[53584] = {-9'd5,10'd395};
ram[53585] = {-9'd2,10'd398};
ram[53586] = {9'd1,-10'd399};
ram[53587] = {9'd4,-10'd396};
ram[53588] = {9'd7,-10'd393};
ram[53589] = {9'd10,-10'd390};
ram[53590] = {9'd14,-10'd387};
ram[53591] = {9'd17,-10'd384};
ram[53592] = {9'd20,-10'd381};
ram[53593] = {9'd23,-10'd377};
ram[53594] = {9'd26,-10'd374};
ram[53595] = {9'd29,-10'd371};
ram[53596] = {9'd32,-10'd368};
ram[53597] = {9'd36,-10'd365};
ram[53598] = {9'd39,-10'd362};
ram[53599] = {9'd42,-10'd359};
ram[53600] = {9'd45,-10'd355};
ram[53601] = {9'd48,-10'd352};
ram[53602] = {9'd51,-10'd349};
ram[53603] = {9'd54,-10'd346};
ram[53604] = {9'd58,-10'd343};
ram[53605] = {9'd61,-10'd340};
ram[53606] = {9'd64,-10'd337};
ram[53607] = {9'd67,-10'd334};
ram[53608] = {9'd70,-10'd330};
ram[53609] = {9'd73,-10'd327};
ram[53610] = {9'd76,-10'd324};
ram[53611] = {9'd80,-10'd321};
ram[53612] = {9'd83,-10'd318};
ram[53613] = {9'd86,-10'd315};
ram[53614] = {9'd89,-10'd312};
ram[53615] = {9'd92,-10'd308};
ram[53616] = {9'd95,-10'd305};
ram[53617] = {9'd98,-10'd302};
ram[53618] = {-9'd99,-10'd299};
ram[53619] = {-9'd96,-10'd296};
ram[53620] = {-9'd92,-10'd293};
ram[53621] = {-9'd89,-10'd290};
ram[53622] = {-9'd86,-10'd286};
ram[53623] = {-9'd83,-10'd283};
ram[53624] = {-9'd80,-10'd280};
ram[53625] = {-9'd77,-10'd277};
ram[53626] = {-9'd74,-10'd274};
ram[53627] = {-9'd70,-10'd271};
ram[53628] = {-9'd67,-10'd268};
ram[53629] = {-9'd64,-10'd264};
ram[53630] = {-9'd61,-10'd261};
ram[53631] = {-9'd58,-10'd258};
ram[53632] = {-9'd58,-10'd258};
ram[53633] = {-9'd55,-10'd255};
ram[53634] = {-9'd52,-10'd252};
ram[53635] = {-9'd48,-10'd249};
ram[53636] = {-9'd45,-10'd246};
ram[53637] = {-9'd42,-10'd242};
ram[53638] = {-9'd39,-10'd239};
ram[53639] = {-9'd36,-10'd236};
ram[53640] = {-9'd33,-10'd233};
ram[53641] = {-9'd30,-10'd230};
ram[53642] = {-9'd26,-10'd227};
ram[53643] = {-9'd23,-10'd224};
ram[53644] = {-9'd20,-10'd220};
ram[53645] = {-9'd17,-10'd217};
ram[53646] = {-9'd14,-10'd214};
ram[53647] = {-9'd11,-10'd211};
ram[53648] = {-9'd8,-10'd208};
ram[53649] = {-9'd4,-10'd205};
ram[53650] = {-9'd1,-10'd202};
ram[53651] = {9'd2,-10'd198};
ram[53652] = {9'd5,-10'd195};
ram[53653] = {9'd8,-10'd192};
ram[53654] = {9'd11,-10'd189};
ram[53655] = {9'd14,-10'd186};
ram[53656] = {9'd18,-10'd183};
ram[53657] = {9'd21,-10'd180};
ram[53658] = {9'd24,-10'd176};
ram[53659] = {9'd27,-10'd173};
ram[53660] = {9'd30,-10'd170};
ram[53661] = {9'd33,-10'd167};
ram[53662] = {9'd36,-10'd164};
ram[53663] = {9'd40,-10'd161};
ram[53664] = {9'd43,-10'd158};
ram[53665] = {9'd46,-10'd154};
ram[53666] = {9'd49,-10'd151};
ram[53667] = {9'd52,-10'd148};
ram[53668] = {9'd55,-10'd145};
ram[53669] = {9'd58,-10'd142};
ram[53670] = {9'd62,-10'd139};
ram[53671] = {9'd65,-10'd136};
ram[53672] = {9'd68,-10'd132};
ram[53673] = {9'd71,-10'd129};
ram[53674] = {9'd74,-10'd126};
ram[53675] = {9'd77,-10'd123};
ram[53676] = {9'd80,-10'd120};
ram[53677] = {9'd84,-10'd117};
ram[53678] = {9'd87,-10'd114};
ram[53679] = {9'd90,-10'd110};
ram[53680] = {9'd93,-10'd107};
ram[53681] = {9'd96,-10'd104};
ram[53682] = {9'd99,-10'd101};
ram[53683] = {-9'd98,-10'd98};
ram[53684] = {-9'd95,-10'd95};
ram[53685] = {-9'd92,-10'd92};
ram[53686] = {-9'd88,-10'd88};
ram[53687] = {-9'd85,-10'd85};
ram[53688] = {-9'd82,-10'd82};
ram[53689] = {-9'd79,-10'd79};
ram[53690] = {-9'd76,-10'd76};
ram[53691] = {-9'd73,-10'd73};
ram[53692] = {-9'd70,-10'd70};
ram[53693] = {-9'd66,-10'd66};
ram[53694] = {-9'd63,-10'd63};
ram[53695] = {-9'd60,-10'd60};
ram[53696] = {-9'd57,-10'd57};
ram[53697] = {-9'd54,-10'd54};
ram[53698] = {-9'd51,-10'd51};
ram[53699] = {-9'd48,-10'd48};
ram[53700] = {-9'd44,-10'd44};
ram[53701] = {-9'd41,-10'd41};
ram[53702] = {-9'd38,-10'd38};
ram[53703] = {-9'd35,-10'd35};
ram[53704] = {-9'd32,-10'd32};
ram[53705] = {-9'd29,-10'd29};
ram[53706] = {-9'd26,-10'd26};
ram[53707] = {-9'd22,-10'd22};
ram[53708] = {-9'd19,-10'd19};
ram[53709] = {-9'd16,-10'd16};
ram[53710] = {-9'd13,-10'd13};
ram[53711] = {-9'd10,-10'd10};
ram[53712] = {-9'd7,-10'd7};
ram[53713] = {-9'd4,-10'd4};
ram[53714] = {9'd0,10'd0};
ram[53715] = {9'd3,10'd3};
ram[53716] = {9'd6,10'd6};
ram[53717] = {9'd9,10'd9};
ram[53718] = {9'd12,10'd12};
ram[53719] = {9'd15,10'd15};
ram[53720] = {9'd18,10'd18};
ram[53721] = {9'd21,10'd21};
ram[53722] = {9'd25,10'd25};
ram[53723] = {9'd28,10'd28};
ram[53724] = {9'd31,10'd31};
ram[53725] = {9'd34,10'd34};
ram[53726] = {9'd37,10'd37};
ram[53727] = {9'd40,10'd40};
ram[53728] = {9'd43,10'd43};
ram[53729] = {9'd47,10'd47};
ram[53730] = {9'd50,10'd50};
ram[53731] = {9'd53,10'd53};
ram[53732] = {9'd56,10'd56};
ram[53733] = {9'd59,10'd59};
ram[53734] = {9'd62,10'd62};
ram[53735] = {9'd65,10'd65};
ram[53736] = {9'd69,10'd69};
ram[53737] = {9'd72,10'd72};
ram[53738] = {9'd75,10'd75};
ram[53739] = {9'd78,10'd78};
ram[53740] = {9'd81,10'd81};
ram[53741] = {9'd84,10'd84};
ram[53742] = {9'd87,10'd87};
ram[53743] = {9'd91,10'd91};
ram[53744] = {9'd94,10'd94};
ram[53745] = {9'd97,10'd97};
ram[53746] = {-9'd100,10'd100};
ram[53747] = {-9'd97,10'd103};
ram[53748] = {-9'd94,10'd106};
ram[53749] = {-9'd91,10'd109};
ram[53750] = {-9'd88,10'd113};
ram[53751] = {-9'd85,10'd116};
ram[53752] = {-9'd81,10'd119};
ram[53753] = {-9'd78,10'd122};
ram[53754] = {-9'd75,10'd125};
ram[53755] = {-9'd72,10'd128};
ram[53756] = {-9'd69,10'd131};
ram[53757] = {-9'd66,10'd135};
ram[53758] = {-9'd63,10'd138};
ram[53759] = {-9'd59,10'd141};
ram[53760] = {-9'd59,10'd141};
ram[53761] = {-9'd56,10'd144};
ram[53762] = {-9'd53,10'd147};
ram[53763] = {-9'd50,10'd150};
ram[53764] = {-9'd47,10'd153};
ram[53765] = {-9'd44,10'd157};
ram[53766] = {-9'd41,10'd160};
ram[53767] = {-9'd37,10'd163};
ram[53768] = {-9'd34,10'd166};
ram[53769] = {-9'd31,10'd169};
ram[53770] = {-9'd28,10'd172};
ram[53771] = {-9'd25,10'd175};
ram[53772] = {-9'd22,10'd179};
ram[53773] = {-9'd19,10'd182};
ram[53774] = {-9'd15,10'd185};
ram[53775] = {-9'd12,10'd188};
ram[53776] = {-9'd9,10'd191};
ram[53777] = {-9'd6,10'd194};
ram[53778] = {-9'd3,10'd197};
ram[53779] = {9'd0,10'd201};
ram[53780] = {9'd3,10'd204};
ram[53781] = {9'd7,10'd207};
ram[53782] = {9'd10,10'd210};
ram[53783] = {9'd13,10'd213};
ram[53784] = {9'd16,10'd216};
ram[53785] = {9'd19,10'd219};
ram[53786] = {9'd22,10'd223};
ram[53787] = {9'd25,10'd226};
ram[53788] = {9'd29,10'd229};
ram[53789] = {9'd32,10'd232};
ram[53790] = {9'd35,10'd235};
ram[53791] = {9'd38,10'd238};
ram[53792] = {9'd41,10'd241};
ram[53793] = {9'd44,10'd245};
ram[53794] = {9'd47,10'd248};
ram[53795] = {9'd51,10'd251};
ram[53796] = {9'd54,10'd254};
ram[53797] = {9'd57,10'd257};
ram[53798] = {9'd60,10'd260};
ram[53799] = {9'd63,10'd263};
ram[53800] = {9'd66,10'd267};
ram[53801] = {9'd69,10'd270};
ram[53802] = {9'd73,10'd273};
ram[53803] = {9'd76,10'd276};
ram[53804] = {9'd79,10'd279};
ram[53805] = {9'd82,10'd282};
ram[53806] = {9'd85,10'd285};
ram[53807] = {9'd88,10'd289};
ram[53808] = {9'd91,10'd292};
ram[53809] = {9'd95,10'd295};
ram[53810] = {9'd98,10'd298};
ram[53811] = {-9'd99,10'd301};
ram[53812] = {-9'd96,10'd304};
ram[53813] = {-9'd93,10'd307};
ram[53814] = {-9'd90,10'd311};
ram[53815] = {-9'd87,10'd314};
ram[53816] = {-9'd84,10'd317};
ram[53817] = {-9'd81,10'd320};
ram[53818] = {-9'd77,10'd323};
ram[53819] = {-9'd74,10'd326};
ram[53820] = {-9'd71,10'd329};
ram[53821] = {-9'd68,10'd333};
ram[53822] = {-9'd65,10'd336};
ram[53823] = {-9'd62,10'd339};
ram[53824] = {-9'd59,10'd342};
ram[53825] = {-9'd55,10'd345};
ram[53826] = {-9'd52,10'd348};
ram[53827] = {-9'd49,10'd351};
ram[53828] = {-9'd46,10'd354};
ram[53829] = {-9'd43,10'd358};
ram[53830] = {-9'd40,10'd361};
ram[53831] = {-9'd37,10'd364};
ram[53832] = {-9'd33,10'd367};
ram[53833] = {-9'd30,10'd370};
ram[53834] = {-9'd27,10'd373};
ram[53835] = {-9'd24,10'd376};
ram[53836] = {-9'd21,10'd380};
ram[53837] = {-9'd18,10'd383};
ram[53838] = {-9'd15,10'd386};
ram[53839] = {-9'd11,10'd389};
ram[53840] = {-9'd8,10'd392};
ram[53841] = {-9'd5,10'd395};
ram[53842] = {-9'd2,10'd398};
ram[53843] = {9'd1,-10'd399};
ram[53844] = {9'd4,-10'd396};
ram[53845] = {9'd7,-10'd393};
ram[53846] = {9'd10,-10'd390};
ram[53847] = {9'd14,-10'd387};
ram[53848] = {9'd17,-10'd384};
ram[53849] = {9'd20,-10'd381};
ram[53850] = {9'd23,-10'd377};
ram[53851] = {9'd26,-10'd374};
ram[53852] = {9'd29,-10'd371};
ram[53853] = {9'd32,-10'd368};
ram[53854] = {9'd36,-10'd365};
ram[53855] = {9'd39,-10'd362};
ram[53856] = {9'd42,-10'd359};
ram[53857] = {9'd45,-10'd355};
ram[53858] = {9'd48,-10'd352};
ram[53859] = {9'd51,-10'd349};
ram[53860] = {9'd54,-10'd346};
ram[53861] = {9'd58,-10'd343};
ram[53862] = {9'd61,-10'd340};
ram[53863] = {9'd64,-10'd337};
ram[53864] = {9'd67,-10'd334};
ram[53865] = {9'd70,-10'd330};
ram[53866] = {9'd73,-10'd327};
ram[53867] = {9'd76,-10'd324};
ram[53868] = {9'd80,-10'd321};
ram[53869] = {9'd83,-10'd318};
ram[53870] = {9'd86,-10'd315};
ram[53871] = {9'd89,-10'd312};
ram[53872] = {9'd92,-10'd308};
ram[53873] = {9'd95,-10'd305};
ram[53874] = {9'd98,-10'd302};
ram[53875] = {-9'd99,-10'd299};
ram[53876] = {-9'd96,-10'd296};
ram[53877] = {-9'd92,-10'd293};
ram[53878] = {-9'd89,-10'd290};
ram[53879] = {-9'd86,-10'd286};
ram[53880] = {-9'd83,-10'd283};
ram[53881] = {-9'd80,-10'd280};
ram[53882] = {-9'd77,-10'd277};
ram[53883] = {-9'd74,-10'd274};
ram[53884] = {-9'd70,-10'd271};
ram[53885] = {-9'd67,-10'd268};
ram[53886] = {-9'd64,-10'd264};
ram[53887] = {-9'd61,-10'd261};
ram[53888] = {-9'd61,-10'd261};
ram[53889] = {-9'd58,-10'd258};
ram[53890] = {-9'd55,-10'd255};
ram[53891] = {-9'd52,-10'd252};
ram[53892] = {-9'd48,-10'd249};
ram[53893] = {-9'd45,-10'd246};
ram[53894] = {-9'd42,-10'd242};
ram[53895] = {-9'd39,-10'd239};
ram[53896] = {-9'd36,-10'd236};
ram[53897] = {-9'd33,-10'd233};
ram[53898] = {-9'd30,-10'd230};
ram[53899] = {-9'd26,-10'd227};
ram[53900] = {-9'd23,-10'd224};
ram[53901] = {-9'd20,-10'd220};
ram[53902] = {-9'd17,-10'd217};
ram[53903] = {-9'd14,-10'd214};
ram[53904] = {-9'd11,-10'd211};
ram[53905] = {-9'd8,-10'd208};
ram[53906] = {-9'd4,-10'd205};
ram[53907] = {-9'd1,-10'd202};
ram[53908] = {9'd2,-10'd198};
ram[53909] = {9'd5,-10'd195};
ram[53910] = {9'd8,-10'd192};
ram[53911] = {9'd11,-10'd189};
ram[53912] = {9'd14,-10'd186};
ram[53913] = {9'd18,-10'd183};
ram[53914] = {9'd21,-10'd180};
ram[53915] = {9'd24,-10'd176};
ram[53916] = {9'd27,-10'd173};
ram[53917] = {9'd30,-10'd170};
ram[53918] = {9'd33,-10'd167};
ram[53919] = {9'd36,-10'd164};
ram[53920] = {9'd40,-10'd161};
ram[53921] = {9'd43,-10'd158};
ram[53922] = {9'd46,-10'd154};
ram[53923] = {9'd49,-10'd151};
ram[53924] = {9'd52,-10'd148};
ram[53925] = {9'd55,-10'd145};
ram[53926] = {9'd58,-10'd142};
ram[53927] = {9'd62,-10'd139};
ram[53928] = {9'd65,-10'd136};
ram[53929] = {9'd68,-10'd132};
ram[53930] = {9'd71,-10'd129};
ram[53931] = {9'd74,-10'd126};
ram[53932] = {9'd77,-10'd123};
ram[53933] = {9'd80,-10'd120};
ram[53934] = {9'd84,-10'd117};
ram[53935] = {9'd87,-10'd114};
ram[53936] = {9'd90,-10'd110};
ram[53937] = {9'd93,-10'd107};
ram[53938] = {9'd96,-10'd104};
ram[53939] = {9'd99,-10'd101};
ram[53940] = {-9'd98,-10'd98};
ram[53941] = {-9'd95,-10'd95};
ram[53942] = {-9'd92,-10'd92};
ram[53943] = {-9'd88,-10'd88};
ram[53944] = {-9'd85,-10'd85};
ram[53945] = {-9'd82,-10'd82};
ram[53946] = {-9'd79,-10'd79};
ram[53947] = {-9'd76,-10'd76};
ram[53948] = {-9'd73,-10'd73};
ram[53949] = {-9'd70,-10'd70};
ram[53950] = {-9'd66,-10'd66};
ram[53951] = {-9'd63,-10'd63};
ram[53952] = {-9'd60,-10'd60};
ram[53953] = {-9'd57,-10'd57};
ram[53954] = {-9'd54,-10'd54};
ram[53955] = {-9'd51,-10'd51};
ram[53956] = {-9'd48,-10'd48};
ram[53957] = {-9'd44,-10'd44};
ram[53958] = {-9'd41,-10'd41};
ram[53959] = {-9'd38,-10'd38};
ram[53960] = {-9'd35,-10'd35};
ram[53961] = {-9'd32,-10'd32};
ram[53962] = {-9'd29,-10'd29};
ram[53963] = {-9'd26,-10'd26};
ram[53964] = {-9'd22,-10'd22};
ram[53965] = {-9'd19,-10'd19};
ram[53966] = {-9'd16,-10'd16};
ram[53967] = {-9'd13,-10'd13};
ram[53968] = {-9'd10,-10'd10};
ram[53969] = {-9'd7,-10'd7};
ram[53970] = {-9'd4,-10'd4};
ram[53971] = {9'd0,10'd0};
ram[53972] = {9'd3,10'd3};
ram[53973] = {9'd6,10'd6};
ram[53974] = {9'd9,10'd9};
ram[53975] = {9'd12,10'd12};
ram[53976] = {9'd15,10'd15};
ram[53977] = {9'd18,10'd18};
ram[53978] = {9'd21,10'd21};
ram[53979] = {9'd25,10'd25};
ram[53980] = {9'd28,10'd28};
ram[53981] = {9'd31,10'd31};
ram[53982] = {9'd34,10'd34};
ram[53983] = {9'd37,10'd37};
ram[53984] = {9'd40,10'd40};
ram[53985] = {9'd43,10'd43};
ram[53986] = {9'd47,10'd47};
ram[53987] = {9'd50,10'd50};
ram[53988] = {9'd53,10'd53};
ram[53989] = {9'd56,10'd56};
ram[53990] = {9'd59,10'd59};
ram[53991] = {9'd62,10'd62};
ram[53992] = {9'd65,10'd65};
ram[53993] = {9'd69,10'd69};
ram[53994] = {9'd72,10'd72};
ram[53995] = {9'd75,10'd75};
ram[53996] = {9'd78,10'd78};
ram[53997] = {9'd81,10'd81};
ram[53998] = {9'd84,10'd84};
ram[53999] = {9'd87,10'd87};
ram[54000] = {9'd91,10'd91};
ram[54001] = {9'd94,10'd94};
ram[54002] = {9'd97,10'd97};
ram[54003] = {-9'd100,10'd100};
ram[54004] = {-9'd97,10'd103};
ram[54005] = {-9'd94,10'd106};
ram[54006] = {-9'd91,10'd109};
ram[54007] = {-9'd88,10'd113};
ram[54008] = {-9'd85,10'd116};
ram[54009] = {-9'd81,10'd119};
ram[54010] = {-9'd78,10'd122};
ram[54011] = {-9'd75,10'd125};
ram[54012] = {-9'd72,10'd128};
ram[54013] = {-9'd69,10'd131};
ram[54014] = {-9'd66,10'd135};
ram[54015] = {-9'd63,10'd138};
ram[54016] = {-9'd63,10'd138};
ram[54017] = {-9'd59,10'd141};
ram[54018] = {-9'd56,10'd144};
ram[54019] = {-9'd53,10'd147};
ram[54020] = {-9'd50,10'd150};
ram[54021] = {-9'd47,10'd153};
ram[54022] = {-9'd44,10'd157};
ram[54023] = {-9'd41,10'd160};
ram[54024] = {-9'd37,10'd163};
ram[54025] = {-9'd34,10'd166};
ram[54026] = {-9'd31,10'd169};
ram[54027] = {-9'd28,10'd172};
ram[54028] = {-9'd25,10'd175};
ram[54029] = {-9'd22,10'd179};
ram[54030] = {-9'd19,10'd182};
ram[54031] = {-9'd15,10'd185};
ram[54032] = {-9'd12,10'd188};
ram[54033] = {-9'd9,10'd191};
ram[54034] = {-9'd6,10'd194};
ram[54035] = {-9'd3,10'd197};
ram[54036] = {9'd0,10'd201};
ram[54037] = {9'd3,10'd204};
ram[54038] = {9'd7,10'd207};
ram[54039] = {9'd10,10'd210};
ram[54040] = {9'd13,10'd213};
ram[54041] = {9'd16,10'd216};
ram[54042] = {9'd19,10'd219};
ram[54043] = {9'd22,10'd223};
ram[54044] = {9'd25,10'd226};
ram[54045] = {9'd29,10'd229};
ram[54046] = {9'd32,10'd232};
ram[54047] = {9'd35,10'd235};
ram[54048] = {9'd38,10'd238};
ram[54049] = {9'd41,10'd241};
ram[54050] = {9'd44,10'd245};
ram[54051] = {9'd47,10'd248};
ram[54052] = {9'd51,10'd251};
ram[54053] = {9'd54,10'd254};
ram[54054] = {9'd57,10'd257};
ram[54055] = {9'd60,10'd260};
ram[54056] = {9'd63,10'd263};
ram[54057] = {9'd66,10'd267};
ram[54058] = {9'd69,10'd270};
ram[54059] = {9'd73,10'd273};
ram[54060] = {9'd76,10'd276};
ram[54061] = {9'd79,10'd279};
ram[54062] = {9'd82,10'd282};
ram[54063] = {9'd85,10'd285};
ram[54064] = {9'd88,10'd289};
ram[54065] = {9'd91,10'd292};
ram[54066] = {9'd95,10'd295};
ram[54067] = {9'd98,10'd298};
ram[54068] = {-9'd99,10'd301};
ram[54069] = {-9'd96,10'd304};
ram[54070] = {-9'd93,10'd307};
ram[54071] = {-9'd90,10'd311};
ram[54072] = {-9'd87,10'd314};
ram[54073] = {-9'd84,10'd317};
ram[54074] = {-9'd81,10'd320};
ram[54075] = {-9'd77,10'd323};
ram[54076] = {-9'd74,10'd326};
ram[54077] = {-9'd71,10'd329};
ram[54078] = {-9'd68,10'd333};
ram[54079] = {-9'd65,10'd336};
ram[54080] = {-9'd62,10'd339};
ram[54081] = {-9'd59,10'd342};
ram[54082] = {-9'd55,10'd345};
ram[54083] = {-9'd52,10'd348};
ram[54084] = {-9'd49,10'd351};
ram[54085] = {-9'd46,10'd354};
ram[54086] = {-9'd43,10'd358};
ram[54087] = {-9'd40,10'd361};
ram[54088] = {-9'd37,10'd364};
ram[54089] = {-9'd33,10'd367};
ram[54090] = {-9'd30,10'd370};
ram[54091] = {-9'd27,10'd373};
ram[54092] = {-9'd24,10'd376};
ram[54093] = {-9'd21,10'd380};
ram[54094] = {-9'd18,10'd383};
ram[54095] = {-9'd15,10'd386};
ram[54096] = {-9'd11,10'd389};
ram[54097] = {-9'd8,10'd392};
ram[54098] = {-9'd5,10'd395};
ram[54099] = {-9'd2,10'd398};
ram[54100] = {9'd1,-10'd399};
ram[54101] = {9'd4,-10'd396};
ram[54102] = {9'd7,-10'd393};
ram[54103] = {9'd10,-10'd390};
ram[54104] = {9'd14,-10'd387};
ram[54105] = {9'd17,-10'd384};
ram[54106] = {9'd20,-10'd381};
ram[54107] = {9'd23,-10'd377};
ram[54108] = {9'd26,-10'd374};
ram[54109] = {9'd29,-10'd371};
ram[54110] = {9'd32,-10'd368};
ram[54111] = {9'd36,-10'd365};
ram[54112] = {9'd39,-10'd362};
ram[54113] = {9'd42,-10'd359};
ram[54114] = {9'd45,-10'd355};
ram[54115] = {9'd48,-10'd352};
ram[54116] = {9'd51,-10'd349};
ram[54117] = {9'd54,-10'd346};
ram[54118] = {9'd58,-10'd343};
ram[54119] = {9'd61,-10'd340};
ram[54120] = {9'd64,-10'd337};
ram[54121] = {9'd67,-10'd334};
ram[54122] = {9'd70,-10'd330};
ram[54123] = {9'd73,-10'd327};
ram[54124] = {9'd76,-10'd324};
ram[54125] = {9'd80,-10'd321};
ram[54126] = {9'd83,-10'd318};
ram[54127] = {9'd86,-10'd315};
ram[54128] = {9'd89,-10'd312};
ram[54129] = {9'd92,-10'd308};
ram[54130] = {9'd95,-10'd305};
ram[54131] = {9'd98,-10'd302};
ram[54132] = {-9'd99,-10'd299};
ram[54133] = {-9'd96,-10'd296};
ram[54134] = {-9'd92,-10'd293};
ram[54135] = {-9'd89,-10'd290};
ram[54136] = {-9'd86,-10'd286};
ram[54137] = {-9'd83,-10'd283};
ram[54138] = {-9'd80,-10'd280};
ram[54139] = {-9'd77,-10'd277};
ram[54140] = {-9'd74,-10'd274};
ram[54141] = {-9'd70,-10'd271};
ram[54142] = {-9'd67,-10'd268};
ram[54143] = {-9'd64,-10'd264};
ram[54144] = {-9'd64,-10'd264};
ram[54145] = {-9'd61,-10'd261};
ram[54146] = {-9'd58,-10'd258};
ram[54147] = {-9'd55,-10'd255};
ram[54148] = {-9'd52,-10'd252};
ram[54149] = {-9'd48,-10'd249};
ram[54150] = {-9'd45,-10'd246};
ram[54151] = {-9'd42,-10'd242};
ram[54152] = {-9'd39,-10'd239};
ram[54153] = {-9'd36,-10'd236};
ram[54154] = {-9'd33,-10'd233};
ram[54155] = {-9'd30,-10'd230};
ram[54156] = {-9'd26,-10'd227};
ram[54157] = {-9'd23,-10'd224};
ram[54158] = {-9'd20,-10'd220};
ram[54159] = {-9'd17,-10'd217};
ram[54160] = {-9'd14,-10'd214};
ram[54161] = {-9'd11,-10'd211};
ram[54162] = {-9'd8,-10'd208};
ram[54163] = {-9'd4,-10'd205};
ram[54164] = {-9'd1,-10'd202};
ram[54165] = {9'd2,-10'd198};
ram[54166] = {9'd5,-10'd195};
ram[54167] = {9'd8,-10'd192};
ram[54168] = {9'd11,-10'd189};
ram[54169] = {9'd14,-10'd186};
ram[54170] = {9'd18,-10'd183};
ram[54171] = {9'd21,-10'd180};
ram[54172] = {9'd24,-10'd176};
ram[54173] = {9'd27,-10'd173};
ram[54174] = {9'd30,-10'd170};
ram[54175] = {9'd33,-10'd167};
ram[54176] = {9'd36,-10'd164};
ram[54177] = {9'd40,-10'd161};
ram[54178] = {9'd43,-10'd158};
ram[54179] = {9'd46,-10'd154};
ram[54180] = {9'd49,-10'd151};
ram[54181] = {9'd52,-10'd148};
ram[54182] = {9'd55,-10'd145};
ram[54183] = {9'd58,-10'd142};
ram[54184] = {9'd62,-10'd139};
ram[54185] = {9'd65,-10'd136};
ram[54186] = {9'd68,-10'd132};
ram[54187] = {9'd71,-10'd129};
ram[54188] = {9'd74,-10'd126};
ram[54189] = {9'd77,-10'd123};
ram[54190] = {9'd80,-10'd120};
ram[54191] = {9'd84,-10'd117};
ram[54192] = {9'd87,-10'd114};
ram[54193] = {9'd90,-10'd110};
ram[54194] = {9'd93,-10'd107};
ram[54195] = {9'd96,-10'd104};
ram[54196] = {9'd99,-10'd101};
ram[54197] = {-9'd98,-10'd98};
ram[54198] = {-9'd95,-10'd95};
ram[54199] = {-9'd92,-10'd92};
ram[54200] = {-9'd88,-10'd88};
ram[54201] = {-9'd85,-10'd85};
ram[54202] = {-9'd82,-10'd82};
ram[54203] = {-9'd79,-10'd79};
ram[54204] = {-9'd76,-10'd76};
ram[54205] = {-9'd73,-10'd73};
ram[54206] = {-9'd70,-10'd70};
ram[54207] = {-9'd66,-10'd66};
ram[54208] = {-9'd63,-10'd63};
ram[54209] = {-9'd60,-10'd60};
ram[54210] = {-9'd57,-10'd57};
ram[54211] = {-9'd54,-10'd54};
ram[54212] = {-9'd51,-10'd51};
ram[54213] = {-9'd48,-10'd48};
ram[54214] = {-9'd44,-10'd44};
ram[54215] = {-9'd41,-10'd41};
ram[54216] = {-9'd38,-10'd38};
ram[54217] = {-9'd35,-10'd35};
ram[54218] = {-9'd32,-10'd32};
ram[54219] = {-9'd29,-10'd29};
ram[54220] = {-9'd26,-10'd26};
ram[54221] = {-9'd22,-10'd22};
ram[54222] = {-9'd19,-10'd19};
ram[54223] = {-9'd16,-10'd16};
ram[54224] = {-9'd13,-10'd13};
ram[54225] = {-9'd10,-10'd10};
ram[54226] = {-9'd7,-10'd7};
ram[54227] = {-9'd4,-10'd4};
ram[54228] = {9'd0,10'd0};
ram[54229] = {9'd3,10'd3};
ram[54230] = {9'd6,10'd6};
ram[54231] = {9'd9,10'd9};
ram[54232] = {9'd12,10'd12};
ram[54233] = {9'd15,10'd15};
ram[54234] = {9'd18,10'd18};
ram[54235] = {9'd21,10'd21};
ram[54236] = {9'd25,10'd25};
ram[54237] = {9'd28,10'd28};
ram[54238] = {9'd31,10'd31};
ram[54239] = {9'd34,10'd34};
ram[54240] = {9'd37,10'd37};
ram[54241] = {9'd40,10'd40};
ram[54242] = {9'd43,10'd43};
ram[54243] = {9'd47,10'd47};
ram[54244] = {9'd50,10'd50};
ram[54245] = {9'd53,10'd53};
ram[54246] = {9'd56,10'd56};
ram[54247] = {9'd59,10'd59};
ram[54248] = {9'd62,10'd62};
ram[54249] = {9'd65,10'd65};
ram[54250] = {9'd69,10'd69};
ram[54251] = {9'd72,10'd72};
ram[54252] = {9'd75,10'd75};
ram[54253] = {9'd78,10'd78};
ram[54254] = {9'd81,10'd81};
ram[54255] = {9'd84,10'd84};
ram[54256] = {9'd87,10'd87};
ram[54257] = {9'd91,10'd91};
ram[54258] = {9'd94,10'd94};
ram[54259] = {9'd97,10'd97};
ram[54260] = {-9'd100,10'd100};
ram[54261] = {-9'd97,10'd103};
ram[54262] = {-9'd94,10'd106};
ram[54263] = {-9'd91,10'd109};
ram[54264] = {-9'd88,10'd113};
ram[54265] = {-9'd85,10'd116};
ram[54266] = {-9'd81,10'd119};
ram[54267] = {-9'd78,10'd122};
ram[54268] = {-9'd75,10'd125};
ram[54269] = {-9'd72,10'd128};
ram[54270] = {-9'd69,10'd131};
ram[54271] = {-9'd66,10'd135};
ram[54272] = {-9'd66,10'd135};
ram[54273] = {-9'd63,10'd138};
ram[54274] = {-9'd59,10'd141};
ram[54275] = {-9'd56,10'd144};
ram[54276] = {-9'd53,10'd147};
ram[54277] = {-9'd50,10'd150};
ram[54278] = {-9'd47,10'd153};
ram[54279] = {-9'd44,10'd157};
ram[54280] = {-9'd41,10'd160};
ram[54281] = {-9'd37,10'd163};
ram[54282] = {-9'd34,10'd166};
ram[54283] = {-9'd31,10'd169};
ram[54284] = {-9'd28,10'd172};
ram[54285] = {-9'd25,10'd175};
ram[54286] = {-9'd22,10'd179};
ram[54287] = {-9'd19,10'd182};
ram[54288] = {-9'd15,10'd185};
ram[54289] = {-9'd12,10'd188};
ram[54290] = {-9'd9,10'd191};
ram[54291] = {-9'd6,10'd194};
ram[54292] = {-9'd3,10'd197};
ram[54293] = {9'd0,10'd201};
ram[54294] = {9'd3,10'd204};
ram[54295] = {9'd7,10'd207};
ram[54296] = {9'd10,10'd210};
ram[54297] = {9'd13,10'd213};
ram[54298] = {9'd16,10'd216};
ram[54299] = {9'd19,10'd219};
ram[54300] = {9'd22,10'd223};
ram[54301] = {9'd25,10'd226};
ram[54302] = {9'd29,10'd229};
ram[54303] = {9'd32,10'd232};
ram[54304] = {9'd35,10'd235};
ram[54305] = {9'd38,10'd238};
ram[54306] = {9'd41,10'd241};
ram[54307] = {9'd44,10'd245};
ram[54308] = {9'd47,10'd248};
ram[54309] = {9'd51,10'd251};
ram[54310] = {9'd54,10'd254};
ram[54311] = {9'd57,10'd257};
ram[54312] = {9'd60,10'd260};
ram[54313] = {9'd63,10'd263};
ram[54314] = {9'd66,10'd267};
ram[54315] = {9'd69,10'd270};
ram[54316] = {9'd73,10'd273};
ram[54317] = {9'd76,10'd276};
ram[54318] = {9'd79,10'd279};
ram[54319] = {9'd82,10'd282};
ram[54320] = {9'd85,10'd285};
ram[54321] = {9'd88,10'd289};
ram[54322] = {9'd91,10'd292};
ram[54323] = {9'd95,10'd295};
ram[54324] = {9'd98,10'd298};
ram[54325] = {-9'd99,10'd301};
ram[54326] = {-9'd96,10'd304};
ram[54327] = {-9'd93,10'd307};
ram[54328] = {-9'd90,10'd311};
ram[54329] = {-9'd87,10'd314};
ram[54330] = {-9'd84,10'd317};
ram[54331] = {-9'd81,10'd320};
ram[54332] = {-9'd77,10'd323};
ram[54333] = {-9'd74,10'd326};
ram[54334] = {-9'd71,10'd329};
ram[54335] = {-9'd68,10'd333};
ram[54336] = {-9'd65,10'd336};
ram[54337] = {-9'd62,10'd339};
ram[54338] = {-9'd59,10'd342};
ram[54339] = {-9'd55,10'd345};
ram[54340] = {-9'd52,10'd348};
ram[54341] = {-9'd49,10'd351};
ram[54342] = {-9'd46,10'd354};
ram[54343] = {-9'd43,10'd358};
ram[54344] = {-9'd40,10'd361};
ram[54345] = {-9'd37,10'd364};
ram[54346] = {-9'd33,10'd367};
ram[54347] = {-9'd30,10'd370};
ram[54348] = {-9'd27,10'd373};
ram[54349] = {-9'd24,10'd376};
ram[54350] = {-9'd21,10'd380};
ram[54351] = {-9'd18,10'd383};
ram[54352] = {-9'd15,10'd386};
ram[54353] = {-9'd11,10'd389};
ram[54354] = {-9'd8,10'd392};
ram[54355] = {-9'd5,10'd395};
ram[54356] = {-9'd2,10'd398};
ram[54357] = {9'd1,-10'd399};
ram[54358] = {9'd4,-10'd396};
ram[54359] = {9'd7,-10'd393};
ram[54360] = {9'd10,-10'd390};
ram[54361] = {9'd14,-10'd387};
ram[54362] = {9'd17,-10'd384};
ram[54363] = {9'd20,-10'd381};
ram[54364] = {9'd23,-10'd377};
ram[54365] = {9'd26,-10'd374};
ram[54366] = {9'd29,-10'd371};
ram[54367] = {9'd32,-10'd368};
ram[54368] = {9'd36,-10'd365};
ram[54369] = {9'd39,-10'd362};
ram[54370] = {9'd42,-10'd359};
ram[54371] = {9'd45,-10'd355};
ram[54372] = {9'd48,-10'd352};
ram[54373] = {9'd51,-10'd349};
ram[54374] = {9'd54,-10'd346};
ram[54375] = {9'd58,-10'd343};
ram[54376] = {9'd61,-10'd340};
ram[54377] = {9'd64,-10'd337};
ram[54378] = {9'd67,-10'd334};
ram[54379] = {9'd70,-10'd330};
ram[54380] = {9'd73,-10'd327};
ram[54381] = {9'd76,-10'd324};
ram[54382] = {9'd80,-10'd321};
ram[54383] = {9'd83,-10'd318};
ram[54384] = {9'd86,-10'd315};
ram[54385] = {9'd89,-10'd312};
ram[54386] = {9'd92,-10'd308};
ram[54387] = {9'd95,-10'd305};
ram[54388] = {9'd98,-10'd302};
ram[54389] = {-9'd99,-10'd299};
ram[54390] = {-9'd96,-10'd296};
ram[54391] = {-9'd92,-10'd293};
ram[54392] = {-9'd89,-10'd290};
ram[54393] = {-9'd86,-10'd286};
ram[54394] = {-9'd83,-10'd283};
ram[54395] = {-9'd80,-10'd280};
ram[54396] = {-9'd77,-10'd277};
ram[54397] = {-9'd74,-10'd274};
ram[54398] = {-9'd70,-10'd271};
ram[54399] = {-9'd67,-10'd268};
ram[54400] = {-9'd67,-10'd268};
ram[54401] = {-9'd64,-10'd264};
ram[54402] = {-9'd61,-10'd261};
ram[54403] = {-9'd58,-10'd258};
ram[54404] = {-9'd55,-10'd255};
ram[54405] = {-9'd52,-10'd252};
ram[54406] = {-9'd48,-10'd249};
ram[54407] = {-9'd45,-10'd246};
ram[54408] = {-9'd42,-10'd242};
ram[54409] = {-9'd39,-10'd239};
ram[54410] = {-9'd36,-10'd236};
ram[54411] = {-9'd33,-10'd233};
ram[54412] = {-9'd30,-10'd230};
ram[54413] = {-9'd26,-10'd227};
ram[54414] = {-9'd23,-10'd224};
ram[54415] = {-9'd20,-10'd220};
ram[54416] = {-9'd17,-10'd217};
ram[54417] = {-9'd14,-10'd214};
ram[54418] = {-9'd11,-10'd211};
ram[54419] = {-9'd8,-10'd208};
ram[54420] = {-9'd4,-10'd205};
ram[54421] = {-9'd1,-10'd202};
ram[54422] = {9'd2,-10'd198};
ram[54423] = {9'd5,-10'd195};
ram[54424] = {9'd8,-10'd192};
ram[54425] = {9'd11,-10'd189};
ram[54426] = {9'd14,-10'd186};
ram[54427] = {9'd18,-10'd183};
ram[54428] = {9'd21,-10'd180};
ram[54429] = {9'd24,-10'd176};
ram[54430] = {9'd27,-10'd173};
ram[54431] = {9'd30,-10'd170};
ram[54432] = {9'd33,-10'd167};
ram[54433] = {9'd36,-10'd164};
ram[54434] = {9'd40,-10'd161};
ram[54435] = {9'd43,-10'd158};
ram[54436] = {9'd46,-10'd154};
ram[54437] = {9'd49,-10'd151};
ram[54438] = {9'd52,-10'd148};
ram[54439] = {9'd55,-10'd145};
ram[54440] = {9'd58,-10'd142};
ram[54441] = {9'd62,-10'd139};
ram[54442] = {9'd65,-10'd136};
ram[54443] = {9'd68,-10'd132};
ram[54444] = {9'd71,-10'd129};
ram[54445] = {9'd74,-10'd126};
ram[54446] = {9'd77,-10'd123};
ram[54447] = {9'd80,-10'd120};
ram[54448] = {9'd84,-10'd117};
ram[54449] = {9'd87,-10'd114};
ram[54450] = {9'd90,-10'd110};
ram[54451] = {9'd93,-10'd107};
ram[54452] = {9'd96,-10'd104};
ram[54453] = {9'd99,-10'd101};
ram[54454] = {-9'd98,-10'd98};
ram[54455] = {-9'd95,-10'd95};
ram[54456] = {-9'd92,-10'd92};
ram[54457] = {-9'd88,-10'd88};
ram[54458] = {-9'd85,-10'd85};
ram[54459] = {-9'd82,-10'd82};
ram[54460] = {-9'd79,-10'd79};
ram[54461] = {-9'd76,-10'd76};
ram[54462] = {-9'd73,-10'd73};
ram[54463] = {-9'd70,-10'd70};
ram[54464] = {-9'd66,-10'd66};
ram[54465] = {-9'd63,-10'd63};
ram[54466] = {-9'd60,-10'd60};
ram[54467] = {-9'd57,-10'd57};
ram[54468] = {-9'd54,-10'd54};
ram[54469] = {-9'd51,-10'd51};
ram[54470] = {-9'd48,-10'd48};
ram[54471] = {-9'd44,-10'd44};
ram[54472] = {-9'd41,-10'd41};
ram[54473] = {-9'd38,-10'd38};
ram[54474] = {-9'd35,-10'd35};
ram[54475] = {-9'd32,-10'd32};
ram[54476] = {-9'd29,-10'd29};
ram[54477] = {-9'd26,-10'd26};
ram[54478] = {-9'd22,-10'd22};
ram[54479] = {-9'd19,-10'd19};
ram[54480] = {-9'd16,-10'd16};
ram[54481] = {-9'd13,-10'd13};
ram[54482] = {-9'd10,-10'd10};
ram[54483] = {-9'd7,-10'd7};
ram[54484] = {-9'd4,-10'd4};
ram[54485] = {9'd0,10'd0};
ram[54486] = {9'd3,10'd3};
ram[54487] = {9'd6,10'd6};
ram[54488] = {9'd9,10'd9};
ram[54489] = {9'd12,10'd12};
ram[54490] = {9'd15,10'd15};
ram[54491] = {9'd18,10'd18};
ram[54492] = {9'd21,10'd21};
ram[54493] = {9'd25,10'd25};
ram[54494] = {9'd28,10'd28};
ram[54495] = {9'd31,10'd31};
ram[54496] = {9'd34,10'd34};
ram[54497] = {9'd37,10'd37};
ram[54498] = {9'd40,10'd40};
ram[54499] = {9'd43,10'd43};
ram[54500] = {9'd47,10'd47};
ram[54501] = {9'd50,10'd50};
ram[54502] = {9'd53,10'd53};
ram[54503] = {9'd56,10'd56};
ram[54504] = {9'd59,10'd59};
ram[54505] = {9'd62,10'd62};
ram[54506] = {9'd65,10'd65};
ram[54507] = {9'd69,10'd69};
ram[54508] = {9'd72,10'd72};
ram[54509] = {9'd75,10'd75};
ram[54510] = {9'd78,10'd78};
ram[54511] = {9'd81,10'd81};
ram[54512] = {9'd84,10'd84};
ram[54513] = {9'd87,10'd87};
ram[54514] = {9'd91,10'd91};
ram[54515] = {9'd94,10'd94};
ram[54516] = {9'd97,10'd97};
ram[54517] = {-9'd100,10'd100};
ram[54518] = {-9'd97,10'd103};
ram[54519] = {-9'd94,10'd106};
ram[54520] = {-9'd91,10'd109};
ram[54521] = {-9'd88,10'd113};
ram[54522] = {-9'd85,10'd116};
ram[54523] = {-9'd81,10'd119};
ram[54524] = {-9'd78,10'd122};
ram[54525] = {-9'd75,10'd125};
ram[54526] = {-9'd72,10'd128};
ram[54527] = {-9'd69,10'd131};
ram[54528] = {-9'd69,10'd131};
ram[54529] = {-9'd66,10'd135};
ram[54530] = {-9'd63,10'd138};
ram[54531] = {-9'd59,10'd141};
ram[54532] = {-9'd56,10'd144};
ram[54533] = {-9'd53,10'd147};
ram[54534] = {-9'd50,10'd150};
ram[54535] = {-9'd47,10'd153};
ram[54536] = {-9'd44,10'd157};
ram[54537] = {-9'd41,10'd160};
ram[54538] = {-9'd37,10'd163};
ram[54539] = {-9'd34,10'd166};
ram[54540] = {-9'd31,10'd169};
ram[54541] = {-9'd28,10'd172};
ram[54542] = {-9'd25,10'd175};
ram[54543] = {-9'd22,10'd179};
ram[54544] = {-9'd19,10'd182};
ram[54545] = {-9'd15,10'd185};
ram[54546] = {-9'd12,10'd188};
ram[54547] = {-9'd9,10'd191};
ram[54548] = {-9'd6,10'd194};
ram[54549] = {-9'd3,10'd197};
ram[54550] = {9'd0,10'd201};
ram[54551] = {9'd3,10'd204};
ram[54552] = {9'd7,10'd207};
ram[54553] = {9'd10,10'd210};
ram[54554] = {9'd13,10'd213};
ram[54555] = {9'd16,10'd216};
ram[54556] = {9'd19,10'd219};
ram[54557] = {9'd22,10'd223};
ram[54558] = {9'd25,10'd226};
ram[54559] = {9'd29,10'd229};
ram[54560] = {9'd32,10'd232};
ram[54561] = {9'd35,10'd235};
ram[54562] = {9'd38,10'd238};
ram[54563] = {9'd41,10'd241};
ram[54564] = {9'd44,10'd245};
ram[54565] = {9'd47,10'd248};
ram[54566] = {9'd51,10'd251};
ram[54567] = {9'd54,10'd254};
ram[54568] = {9'd57,10'd257};
ram[54569] = {9'd60,10'd260};
ram[54570] = {9'd63,10'd263};
ram[54571] = {9'd66,10'd267};
ram[54572] = {9'd69,10'd270};
ram[54573] = {9'd73,10'd273};
ram[54574] = {9'd76,10'd276};
ram[54575] = {9'd79,10'd279};
ram[54576] = {9'd82,10'd282};
ram[54577] = {9'd85,10'd285};
ram[54578] = {9'd88,10'd289};
ram[54579] = {9'd91,10'd292};
ram[54580] = {9'd95,10'd295};
ram[54581] = {9'd98,10'd298};
ram[54582] = {-9'd99,10'd301};
ram[54583] = {-9'd96,10'd304};
ram[54584] = {-9'd93,10'd307};
ram[54585] = {-9'd90,10'd311};
ram[54586] = {-9'd87,10'd314};
ram[54587] = {-9'd84,10'd317};
ram[54588] = {-9'd81,10'd320};
ram[54589] = {-9'd77,10'd323};
ram[54590] = {-9'd74,10'd326};
ram[54591] = {-9'd71,10'd329};
ram[54592] = {-9'd68,10'd333};
ram[54593] = {-9'd65,10'd336};
ram[54594] = {-9'd62,10'd339};
ram[54595] = {-9'd59,10'd342};
ram[54596] = {-9'd55,10'd345};
ram[54597] = {-9'd52,10'd348};
ram[54598] = {-9'd49,10'd351};
ram[54599] = {-9'd46,10'd354};
ram[54600] = {-9'd43,10'd358};
ram[54601] = {-9'd40,10'd361};
ram[54602] = {-9'd37,10'd364};
ram[54603] = {-9'd33,10'd367};
ram[54604] = {-9'd30,10'd370};
ram[54605] = {-9'd27,10'd373};
ram[54606] = {-9'd24,10'd376};
ram[54607] = {-9'd21,10'd380};
ram[54608] = {-9'd18,10'd383};
ram[54609] = {-9'd15,10'd386};
ram[54610] = {-9'd11,10'd389};
ram[54611] = {-9'd8,10'd392};
ram[54612] = {-9'd5,10'd395};
ram[54613] = {-9'd2,10'd398};
ram[54614] = {9'd1,-10'd399};
ram[54615] = {9'd4,-10'd396};
ram[54616] = {9'd7,-10'd393};
ram[54617] = {9'd10,-10'd390};
ram[54618] = {9'd14,-10'd387};
ram[54619] = {9'd17,-10'd384};
ram[54620] = {9'd20,-10'd381};
ram[54621] = {9'd23,-10'd377};
ram[54622] = {9'd26,-10'd374};
ram[54623] = {9'd29,-10'd371};
ram[54624] = {9'd32,-10'd368};
ram[54625] = {9'd36,-10'd365};
ram[54626] = {9'd39,-10'd362};
ram[54627] = {9'd42,-10'd359};
ram[54628] = {9'd45,-10'd355};
ram[54629] = {9'd48,-10'd352};
ram[54630] = {9'd51,-10'd349};
ram[54631] = {9'd54,-10'd346};
ram[54632] = {9'd58,-10'd343};
ram[54633] = {9'd61,-10'd340};
ram[54634] = {9'd64,-10'd337};
ram[54635] = {9'd67,-10'd334};
ram[54636] = {9'd70,-10'd330};
ram[54637] = {9'd73,-10'd327};
ram[54638] = {9'd76,-10'd324};
ram[54639] = {9'd80,-10'd321};
ram[54640] = {9'd83,-10'd318};
ram[54641] = {9'd86,-10'd315};
ram[54642] = {9'd89,-10'd312};
ram[54643] = {9'd92,-10'd308};
ram[54644] = {9'd95,-10'd305};
ram[54645] = {9'd98,-10'd302};
ram[54646] = {-9'd99,-10'd299};
ram[54647] = {-9'd96,-10'd296};
ram[54648] = {-9'd92,-10'd293};
ram[54649] = {-9'd89,-10'd290};
ram[54650] = {-9'd86,-10'd286};
ram[54651] = {-9'd83,-10'd283};
ram[54652] = {-9'd80,-10'd280};
ram[54653] = {-9'd77,-10'd277};
ram[54654] = {-9'd74,-10'd274};
ram[54655] = {-9'd70,-10'd271};
ram[54656] = {-9'd70,-10'd271};
ram[54657] = {-9'd67,-10'd268};
ram[54658] = {-9'd64,-10'd264};
ram[54659] = {-9'd61,-10'd261};
ram[54660] = {-9'd58,-10'd258};
ram[54661] = {-9'd55,-10'd255};
ram[54662] = {-9'd52,-10'd252};
ram[54663] = {-9'd48,-10'd249};
ram[54664] = {-9'd45,-10'd246};
ram[54665] = {-9'd42,-10'd242};
ram[54666] = {-9'd39,-10'd239};
ram[54667] = {-9'd36,-10'd236};
ram[54668] = {-9'd33,-10'd233};
ram[54669] = {-9'd30,-10'd230};
ram[54670] = {-9'd26,-10'd227};
ram[54671] = {-9'd23,-10'd224};
ram[54672] = {-9'd20,-10'd220};
ram[54673] = {-9'd17,-10'd217};
ram[54674] = {-9'd14,-10'd214};
ram[54675] = {-9'd11,-10'd211};
ram[54676] = {-9'd8,-10'd208};
ram[54677] = {-9'd4,-10'd205};
ram[54678] = {-9'd1,-10'd202};
ram[54679] = {9'd2,-10'd198};
ram[54680] = {9'd5,-10'd195};
ram[54681] = {9'd8,-10'd192};
ram[54682] = {9'd11,-10'd189};
ram[54683] = {9'd14,-10'd186};
ram[54684] = {9'd18,-10'd183};
ram[54685] = {9'd21,-10'd180};
ram[54686] = {9'd24,-10'd176};
ram[54687] = {9'd27,-10'd173};
ram[54688] = {9'd30,-10'd170};
ram[54689] = {9'd33,-10'd167};
ram[54690] = {9'd36,-10'd164};
ram[54691] = {9'd40,-10'd161};
ram[54692] = {9'd43,-10'd158};
ram[54693] = {9'd46,-10'd154};
ram[54694] = {9'd49,-10'd151};
ram[54695] = {9'd52,-10'd148};
ram[54696] = {9'd55,-10'd145};
ram[54697] = {9'd58,-10'd142};
ram[54698] = {9'd62,-10'd139};
ram[54699] = {9'd65,-10'd136};
ram[54700] = {9'd68,-10'd132};
ram[54701] = {9'd71,-10'd129};
ram[54702] = {9'd74,-10'd126};
ram[54703] = {9'd77,-10'd123};
ram[54704] = {9'd80,-10'd120};
ram[54705] = {9'd84,-10'd117};
ram[54706] = {9'd87,-10'd114};
ram[54707] = {9'd90,-10'd110};
ram[54708] = {9'd93,-10'd107};
ram[54709] = {9'd96,-10'd104};
ram[54710] = {9'd99,-10'd101};
ram[54711] = {-9'd98,-10'd98};
ram[54712] = {-9'd95,-10'd95};
ram[54713] = {-9'd92,-10'd92};
ram[54714] = {-9'd88,-10'd88};
ram[54715] = {-9'd85,-10'd85};
ram[54716] = {-9'd82,-10'd82};
ram[54717] = {-9'd79,-10'd79};
ram[54718] = {-9'd76,-10'd76};
ram[54719] = {-9'd73,-10'd73};
ram[54720] = {-9'd70,-10'd70};
ram[54721] = {-9'd66,-10'd66};
ram[54722] = {-9'd63,-10'd63};
ram[54723] = {-9'd60,-10'd60};
ram[54724] = {-9'd57,-10'd57};
ram[54725] = {-9'd54,-10'd54};
ram[54726] = {-9'd51,-10'd51};
ram[54727] = {-9'd48,-10'd48};
ram[54728] = {-9'd44,-10'd44};
ram[54729] = {-9'd41,-10'd41};
ram[54730] = {-9'd38,-10'd38};
ram[54731] = {-9'd35,-10'd35};
ram[54732] = {-9'd32,-10'd32};
ram[54733] = {-9'd29,-10'd29};
ram[54734] = {-9'd26,-10'd26};
ram[54735] = {-9'd22,-10'd22};
ram[54736] = {-9'd19,-10'd19};
ram[54737] = {-9'd16,-10'd16};
ram[54738] = {-9'd13,-10'd13};
ram[54739] = {-9'd10,-10'd10};
ram[54740] = {-9'd7,-10'd7};
ram[54741] = {-9'd4,-10'd4};
ram[54742] = {9'd0,10'd0};
ram[54743] = {9'd3,10'd3};
ram[54744] = {9'd6,10'd6};
ram[54745] = {9'd9,10'd9};
ram[54746] = {9'd12,10'd12};
ram[54747] = {9'd15,10'd15};
ram[54748] = {9'd18,10'd18};
ram[54749] = {9'd21,10'd21};
ram[54750] = {9'd25,10'd25};
ram[54751] = {9'd28,10'd28};
ram[54752] = {9'd31,10'd31};
ram[54753] = {9'd34,10'd34};
ram[54754] = {9'd37,10'd37};
ram[54755] = {9'd40,10'd40};
ram[54756] = {9'd43,10'd43};
ram[54757] = {9'd47,10'd47};
ram[54758] = {9'd50,10'd50};
ram[54759] = {9'd53,10'd53};
ram[54760] = {9'd56,10'd56};
ram[54761] = {9'd59,10'd59};
ram[54762] = {9'd62,10'd62};
ram[54763] = {9'd65,10'd65};
ram[54764] = {9'd69,10'd69};
ram[54765] = {9'd72,10'd72};
ram[54766] = {9'd75,10'd75};
ram[54767] = {9'd78,10'd78};
ram[54768] = {9'd81,10'd81};
ram[54769] = {9'd84,10'd84};
ram[54770] = {9'd87,10'd87};
ram[54771] = {9'd91,10'd91};
ram[54772] = {9'd94,10'd94};
ram[54773] = {9'd97,10'd97};
ram[54774] = {-9'd100,10'd100};
ram[54775] = {-9'd97,10'd103};
ram[54776] = {-9'd94,10'd106};
ram[54777] = {-9'd91,10'd109};
ram[54778] = {-9'd88,10'd113};
ram[54779] = {-9'd85,10'd116};
ram[54780] = {-9'd81,10'd119};
ram[54781] = {-9'd78,10'd122};
ram[54782] = {-9'd75,10'd125};
ram[54783] = {-9'd72,10'd128};
ram[54784] = {-9'd72,10'd128};
ram[54785] = {-9'd69,10'd131};
ram[54786] = {-9'd66,10'd135};
ram[54787] = {-9'd63,10'd138};
ram[54788] = {-9'd59,10'd141};
ram[54789] = {-9'd56,10'd144};
ram[54790] = {-9'd53,10'd147};
ram[54791] = {-9'd50,10'd150};
ram[54792] = {-9'd47,10'd153};
ram[54793] = {-9'd44,10'd157};
ram[54794] = {-9'd41,10'd160};
ram[54795] = {-9'd37,10'd163};
ram[54796] = {-9'd34,10'd166};
ram[54797] = {-9'd31,10'd169};
ram[54798] = {-9'd28,10'd172};
ram[54799] = {-9'd25,10'd175};
ram[54800] = {-9'd22,10'd179};
ram[54801] = {-9'd19,10'd182};
ram[54802] = {-9'd15,10'd185};
ram[54803] = {-9'd12,10'd188};
ram[54804] = {-9'd9,10'd191};
ram[54805] = {-9'd6,10'd194};
ram[54806] = {-9'd3,10'd197};
ram[54807] = {9'd0,10'd201};
ram[54808] = {9'd3,10'd204};
ram[54809] = {9'd7,10'd207};
ram[54810] = {9'd10,10'd210};
ram[54811] = {9'd13,10'd213};
ram[54812] = {9'd16,10'd216};
ram[54813] = {9'd19,10'd219};
ram[54814] = {9'd22,10'd223};
ram[54815] = {9'd25,10'd226};
ram[54816] = {9'd29,10'd229};
ram[54817] = {9'd32,10'd232};
ram[54818] = {9'd35,10'd235};
ram[54819] = {9'd38,10'd238};
ram[54820] = {9'd41,10'd241};
ram[54821] = {9'd44,10'd245};
ram[54822] = {9'd47,10'd248};
ram[54823] = {9'd51,10'd251};
ram[54824] = {9'd54,10'd254};
ram[54825] = {9'd57,10'd257};
ram[54826] = {9'd60,10'd260};
ram[54827] = {9'd63,10'd263};
ram[54828] = {9'd66,10'd267};
ram[54829] = {9'd69,10'd270};
ram[54830] = {9'd73,10'd273};
ram[54831] = {9'd76,10'd276};
ram[54832] = {9'd79,10'd279};
ram[54833] = {9'd82,10'd282};
ram[54834] = {9'd85,10'd285};
ram[54835] = {9'd88,10'd289};
ram[54836] = {9'd91,10'd292};
ram[54837] = {9'd95,10'd295};
ram[54838] = {9'd98,10'd298};
ram[54839] = {-9'd99,10'd301};
ram[54840] = {-9'd96,10'd304};
ram[54841] = {-9'd93,10'd307};
ram[54842] = {-9'd90,10'd311};
ram[54843] = {-9'd87,10'd314};
ram[54844] = {-9'd84,10'd317};
ram[54845] = {-9'd81,10'd320};
ram[54846] = {-9'd77,10'd323};
ram[54847] = {-9'd74,10'd326};
ram[54848] = {-9'd71,10'd329};
ram[54849] = {-9'd68,10'd333};
ram[54850] = {-9'd65,10'd336};
ram[54851] = {-9'd62,10'd339};
ram[54852] = {-9'd59,10'd342};
ram[54853] = {-9'd55,10'd345};
ram[54854] = {-9'd52,10'd348};
ram[54855] = {-9'd49,10'd351};
ram[54856] = {-9'd46,10'd354};
ram[54857] = {-9'd43,10'd358};
ram[54858] = {-9'd40,10'd361};
ram[54859] = {-9'd37,10'd364};
ram[54860] = {-9'd33,10'd367};
ram[54861] = {-9'd30,10'd370};
ram[54862] = {-9'd27,10'd373};
ram[54863] = {-9'd24,10'd376};
ram[54864] = {-9'd21,10'd380};
ram[54865] = {-9'd18,10'd383};
ram[54866] = {-9'd15,10'd386};
ram[54867] = {-9'd11,10'd389};
ram[54868] = {-9'd8,10'd392};
ram[54869] = {-9'd5,10'd395};
ram[54870] = {-9'd2,10'd398};
ram[54871] = {9'd1,-10'd399};
ram[54872] = {9'd4,-10'd396};
ram[54873] = {9'd7,-10'd393};
ram[54874] = {9'd10,-10'd390};
ram[54875] = {9'd14,-10'd387};
ram[54876] = {9'd17,-10'd384};
ram[54877] = {9'd20,-10'd381};
ram[54878] = {9'd23,-10'd377};
ram[54879] = {9'd26,-10'd374};
ram[54880] = {9'd29,-10'd371};
ram[54881] = {9'd32,-10'd368};
ram[54882] = {9'd36,-10'd365};
ram[54883] = {9'd39,-10'd362};
ram[54884] = {9'd42,-10'd359};
ram[54885] = {9'd45,-10'd355};
ram[54886] = {9'd48,-10'd352};
ram[54887] = {9'd51,-10'd349};
ram[54888] = {9'd54,-10'd346};
ram[54889] = {9'd58,-10'd343};
ram[54890] = {9'd61,-10'd340};
ram[54891] = {9'd64,-10'd337};
ram[54892] = {9'd67,-10'd334};
ram[54893] = {9'd70,-10'd330};
ram[54894] = {9'd73,-10'd327};
ram[54895] = {9'd76,-10'd324};
ram[54896] = {9'd80,-10'd321};
ram[54897] = {9'd83,-10'd318};
ram[54898] = {9'd86,-10'd315};
ram[54899] = {9'd89,-10'd312};
ram[54900] = {9'd92,-10'd308};
ram[54901] = {9'd95,-10'd305};
ram[54902] = {9'd98,-10'd302};
ram[54903] = {-9'd99,-10'd299};
ram[54904] = {-9'd96,-10'd296};
ram[54905] = {-9'd92,-10'd293};
ram[54906] = {-9'd89,-10'd290};
ram[54907] = {-9'd86,-10'd286};
ram[54908] = {-9'd83,-10'd283};
ram[54909] = {-9'd80,-10'd280};
ram[54910] = {-9'd77,-10'd277};
ram[54911] = {-9'd74,-10'd274};
ram[54912] = {-9'd74,-10'd274};
ram[54913] = {-9'd70,-10'd271};
ram[54914] = {-9'd67,-10'd268};
ram[54915] = {-9'd64,-10'd264};
ram[54916] = {-9'd61,-10'd261};
ram[54917] = {-9'd58,-10'd258};
ram[54918] = {-9'd55,-10'd255};
ram[54919] = {-9'd52,-10'd252};
ram[54920] = {-9'd48,-10'd249};
ram[54921] = {-9'd45,-10'd246};
ram[54922] = {-9'd42,-10'd242};
ram[54923] = {-9'd39,-10'd239};
ram[54924] = {-9'd36,-10'd236};
ram[54925] = {-9'd33,-10'd233};
ram[54926] = {-9'd30,-10'd230};
ram[54927] = {-9'd26,-10'd227};
ram[54928] = {-9'd23,-10'd224};
ram[54929] = {-9'd20,-10'd220};
ram[54930] = {-9'd17,-10'd217};
ram[54931] = {-9'd14,-10'd214};
ram[54932] = {-9'd11,-10'd211};
ram[54933] = {-9'd8,-10'd208};
ram[54934] = {-9'd4,-10'd205};
ram[54935] = {-9'd1,-10'd202};
ram[54936] = {9'd2,-10'd198};
ram[54937] = {9'd5,-10'd195};
ram[54938] = {9'd8,-10'd192};
ram[54939] = {9'd11,-10'd189};
ram[54940] = {9'd14,-10'd186};
ram[54941] = {9'd18,-10'd183};
ram[54942] = {9'd21,-10'd180};
ram[54943] = {9'd24,-10'd176};
ram[54944] = {9'd27,-10'd173};
ram[54945] = {9'd30,-10'd170};
ram[54946] = {9'd33,-10'd167};
ram[54947] = {9'd36,-10'd164};
ram[54948] = {9'd40,-10'd161};
ram[54949] = {9'd43,-10'd158};
ram[54950] = {9'd46,-10'd154};
ram[54951] = {9'd49,-10'd151};
ram[54952] = {9'd52,-10'd148};
ram[54953] = {9'd55,-10'd145};
ram[54954] = {9'd58,-10'd142};
ram[54955] = {9'd62,-10'd139};
ram[54956] = {9'd65,-10'd136};
ram[54957] = {9'd68,-10'd132};
ram[54958] = {9'd71,-10'd129};
ram[54959] = {9'd74,-10'd126};
ram[54960] = {9'd77,-10'd123};
ram[54961] = {9'd80,-10'd120};
ram[54962] = {9'd84,-10'd117};
ram[54963] = {9'd87,-10'd114};
ram[54964] = {9'd90,-10'd110};
ram[54965] = {9'd93,-10'd107};
ram[54966] = {9'd96,-10'd104};
ram[54967] = {9'd99,-10'd101};
ram[54968] = {-9'd98,-10'd98};
ram[54969] = {-9'd95,-10'd95};
ram[54970] = {-9'd92,-10'd92};
ram[54971] = {-9'd88,-10'd88};
ram[54972] = {-9'd85,-10'd85};
ram[54973] = {-9'd82,-10'd82};
ram[54974] = {-9'd79,-10'd79};
ram[54975] = {-9'd76,-10'd76};
ram[54976] = {-9'd73,-10'd73};
ram[54977] = {-9'd70,-10'd70};
ram[54978] = {-9'd66,-10'd66};
ram[54979] = {-9'd63,-10'd63};
ram[54980] = {-9'd60,-10'd60};
ram[54981] = {-9'd57,-10'd57};
ram[54982] = {-9'd54,-10'd54};
ram[54983] = {-9'd51,-10'd51};
ram[54984] = {-9'd48,-10'd48};
ram[54985] = {-9'd44,-10'd44};
ram[54986] = {-9'd41,-10'd41};
ram[54987] = {-9'd38,-10'd38};
ram[54988] = {-9'd35,-10'd35};
ram[54989] = {-9'd32,-10'd32};
ram[54990] = {-9'd29,-10'd29};
ram[54991] = {-9'd26,-10'd26};
ram[54992] = {-9'd22,-10'd22};
ram[54993] = {-9'd19,-10'd19};
ram[54994] = {-9'd16,-10'd16};
ram[54995] = {-9'd13,-10'd13};
ram[54996] = {-9'd10,-10'd10};
ram[54997] = {-9'd7,-10'd7};
ram[54998] = {-9'd4,-10'd4};
ram[54999] = {9'd0,10'd0};
ram[55000] = {9'd3,10'd3};
ram[55001] = {9'd6,10'd6};
ram[55002] = {9'd9,10'd9};
ram[55003] = {9'd12,10'd12};
ram[55004] = {9'd15,10'd15};
ram[55005] = {9'd18,10'd18};
ram[55006] = {9'd21,10'd21};
ram[55007] = {9'd25,10'd25};
ram[55008] = {9'd28,10'd28};
ram[55009] = {9'd31,10'd31};
ram[55010] = {9'd34,10'd34};
ram[55011] = {9'd37,10'd37};
ram[55012] = {9'd40,10'd40};
ram[55013] = {9'd43,10'd43};
ram[55014] = {9'd47,10'd47};
ram[55015] = {9'd50,10'd50};
ram[55016] = {9'd53,10'd53};
ram[55017] = {9'd56,10'd56};
ram[55018] = {9'd59,10'd59};
ram[55019] = {9'd62,10'd62};
ram[55020] = {9'd65,10'd65};
ram[55021] = {9'd69,10'd69};
ram[55022] = {9'd72,10'd72};
ram[55023] = {9'd75,10'd75};
ram[55024] = {9'd78,10'd78};
ram[55025] = {9'd81,10'd81};
ram[55026] = {9'd84,10'd84};
ram[55027] = {9'd87,10'd87};
ram[55028] = {9'd91,10'd91};
ram[55029] = {9'd94,10'd94};
ram[55030] = {9'd97,10'd97};
ram[55031] = {-9'd100,10'd100};
ram[55032] = {-9'd97,10'd103};
ram[55033] = {-9'd94,10'd106};
ram[55034] = {-9'd91,10'd109};
ram[55035] = {-9'd88,10'd113};
ram[55036] = {-9'd85,10'd116};
ram[55037] = {-9'd81,10'd119};
ram[55038] = {-9'd78,10'd122};
ram[55039] = {-9'd75,10'd125};
ram[55040] = {-9'd75,10'd125};
ram[55041] = {-9'd72,10'd128};
ram[55042] = {-9'd69,10'd131};
ram[55043] = {-9'd66,10'd135};
ram[55044] = {-9'd63,10'd138};
ram[55045] = {-9'd59,10'd141};
ram[55046] = {-9'd56,10'd144};
ram[55047] = {-9'd53,10'd147};
ram[55048] = {-9'd50,10'd150};
ram[55049] = {-9'd47,10'd153};
ram[55050] = {-9'd44,10'd157};
ram[55051] = {-9'd41,10'd160};
ram[55052] = {-9'd37,10'd163};
ram[55053] = {-9'd34,10'd166};
ram[55054] = {-9'd31,10'd169};
ram[55055] = {-9'd28,10'd172};
ram[55056] = {-9'd25,10'd175};
ram[55057] = {-9'd22,10'd179};
ram[55058] = {-9'd19,10'd182};
ram[55059] = {-9'd15,10'd185};
ram[55060] = {-9'd12,10'd188};
ram[55061] = {-9'd9,10'd191};
ram[55062] = {-9'd6,10'd194};
ram[55063] = {-9'd3,10'd197};
ram[55064] = {9'd0,10'd201};
ram[55065] = {9'd3,10'd204};
ram[55066] = {9'd7,10'd207};
ram[55067] = {9'd10,10'd210};
ram[55068] = {9'd13,10'd213};
ram[55069] = {9'd16,10'd216};
ram[55070] = {9'd19,10'd219};
ram[55071] = {9'd22,10'd223};
ram[55072] = {9'd25,10'd226};
ram[55073] = {9'd29,10'd229};
ram[55074] = {9'd32,10'd232};
ram[55075] = {9'd35,10'd235};
ram[55076] = {9'd38,10'd238};
ram[55077] = {9'd41,10'd241};
ram[55078] = {9'd44,10'd245};
ram[55079] = {9'd47,10'd248};
ram[55080] = {9'd51,10'd251};
ram[55081] = {9'd54,10'd254};
ram[55082] = {9'd57,10'd257};
ram[55083] = {9'd60,10'd260};
ram[55084] = {9'd63,10'd263};
ram[55085] = {9'd66,10'd267};
ram[55086] = {9'd69,10'd270};
ram[55087] = {9'd73,10'd273};
ram[55088] = {9'd76,10'd276};
ram[55089] = {9'd79,10'd279};
ram[55090] = {9'd82,10'd282};
ram[55091] = {9'd85,10'd285};
ram[55092] = {9'd88,10'd289};
ram[55093] = {9'd91,10'd292};
ram[55094] = {9'd95,10'd295};
ram[55095] = {9'd98,10'd298};
ram[55096] = {-9'd99,10'd301};
ram[55097] = {-9'd96,10'd304};
ram[55098] = {-9'd93,10'd307};
ram[55099] = {-9'd90,10'd311};
ram[55100] = {-9'd87,10'd314};
ram[55101] = {-9'd84,10'd317};
ram[55102] = {-9'd81,10'd320};
ram[55103] = {-9'd77,10'd323};
ram[55104] = {-9'd74,10'd326};
ram[55105] = {-9'd71,10'd329};
ram[55106] = {-9'd68,10'd333};
ram[55107] = {-9'd65,10'd336};
ram[55108] = {-9'd62,10'd339};
ram[55109] = {-9'd59,10'd342};
ram[55110] = {-9'd55,10'd345};
ram[55111] = {-9'd52,10'd348};
ram[55112] = {-9'd49,10'd351};
ram[55113] = {-9'd46,10'd354};
ram[55114] = {-9'd43,10'd358};
ram[55115] = {-9'd40,10'd361};
ram[55116] = {-9'd37,10'd364};
ram[55117] = {-9'd33,10'd367};
ram[55118] = {-9'd30,10'd370};
ram[55119] = {-9'd27,10'd373};
ram[55120] = {-9'd24,10'd376};
ram[55121] = {-9'd21,10'd380};
ram[55122] = {-9'd18,10'd383};
ram[55123] = {-9'd15,10'd386};
ram[55124] = {-9'd11,10'd389};
ram[55125] = {-9'd8,10'd392};
ram[55126] = {-9'd5,10'd395};
ram[55127] = {-9'd2,10'd398};
ram[55128] = {9'd1,-10'd399};
ram[55129] = {9'd4,-10'd396};
ram[55130] = {9'd7,-10'd393};
ram[55131] = {9'd10,-10'd390};
ram[55132] = {9'd14,-10'd387};
ram[55133] = {9'd17,-10'd384};
ram[55134] = {9'd20,-10'd381};
ram[55135] = {9'd23,-10'd377};
ram[55136] = {9'd26,-10'd374};
ram[55137] = {9'd29,-10'd371};
ram[55138] = {9'd32,-10'd368};
ram[55139] = {9'd36,-10'd365};
ram[55140] = {9'd39,-10'd362};
ram[55141] = {9'd42,-10'd359};
ram[55142] = {9'd45,-10'd355};
ram[55143] = {9'd48,-10'd352};
ram[55144] = {9'd51,-10'd349};
ram[55145] = {9'd54,-10'd346};
ram[55146] = {9'd58,-10'd343};
ram[55147] = {9'd61,-10'd340};
ram[55148] = {9'd64,-10'd337};
ram[55149] = {9'd67,-10'd334};
ram[55150] = {9'd70,-10'd330};
ram[55151] = {9'd73,-10'd327};
ram[55152] = {9'd76,-10'd324};
ram[55153] = {9'd80,-10'd321};
ram[55154] = {9'd83,-10'd318};
ram[55155] = {9'd86,-10'd315};
ram[55156] = {9'd89,-10'd312};
ram[55157] = {9'd92,-10'd308};
ram[55158] = {9'd95,-10'd305};
ram[55159] = {9'd98,-10'd302};
ram[55160] = {-9'd99,-10'd299};
ram[55161] = {-9'd96,-10'd296};
ram[55162] = {-9'd92,-10'd293};
ram[55163] = {-9'd89,-10'd290};
ram[55164] = {-9'd86,-10'd286};
ram[55165] = {-9'd83,-10'd283};
ram[55166] = {-9'd80,-10'd280};
ram[55167] = {-9'd77,-10'd277};
ram[55168] = {-9'd77,-10'd277};
ram[55169] = {-9'd74,-10'd274};
ram[55170] = {-9'd70,-10'd271};
ram[55171] = {-9'd67,-10'd268};
ram[55172] = {-9'd64,-10'd264};
ram[55173] = {-9'd61,-10'd261};
ram[55174] = {-9'd58,-10'd258};
ram[55175] = {-9'd55,-10'd255};
ram[55176] = {-9'd52,-10'd252};
ram[55177] = {-9'd48,-10'd249};
ram[55178] = {-9'd45,-10'd246};
ram[55179] = {-9'd42,-10'd242};
ram[55180] = {-9'd39,-10'd239};
ram[55181] = {-9'd36,-10'd236};
ram[55182] = {-9'd33,-10'd233};
ram[55183] = {-9'd30,-10'd230};
ram[55184] = {-9'd26,-10'd227};
ram[55185] = {-9'd23,-10'd224};
ram[55186] = {-9'd20,-10'd220};
ram[55187] = {-9'd17,-10'd217};
ram[55188] = {-9'd14,-10'd214};
ram[55189] = {-9'd11,-10'd211};
ram[55190] = {-9'd8,-10'd208};
ram[55191] = {-9'd4,-10'd205};
ram[55192] = {-9'd1,-10'd202};
ram[55193] = {9'd2,-10'd198};
ram[55194] = {9'd5,-10'd195};
ram[55195] = {9'd8,-10'd192};
ram[55196] = {9'd11,-10'd189};
ram[55197] = {9'd14,-10'd186};
ram[55198] = {9'd18,-10'd183};
ram[55199] = {9'd21,-10'd180};
ram[55200] = {9'd24,-10'd176};
ram[55201] = {9'd27,-10'd173};
ram[55202] = {9'd30,-10'd170};
ram[55203] = {9'd33,-10'd167};
ram[55204] = {9'd36,-10'd164};
ram[55205] = {9'd40,-10'd161};
ram[55206] = {9'd43,-10'd158};
ram[55207] = {9'd46,-10'd154};
ram[55208] = {9'd49,-10'd151};
ram[55209] = {9'd52,-10'd148};
ram[55210] = {9'd55,-10'd145};
ram[55211] = {9'd58,-10'd142};
ram[55212] = {9'd62,-10'd139};
ram[55213] = {9'd65,-10'd136};
ram[55214] = {9'd68,-10'd132};
ram[55215] = {9'd71,-10'd129};
ram[55216] = {9'd74,-10'd126};
ram[55217] = {9'd77,-10'd123};
ram[55218] = {9'd80,-10'd120};
ram[55219] = {9'd84,-10'd117};
ram[55220] = {9'd87,-10'd114};
ram[55221] = {9'd90,-10'd110};
ram[55222] = {9'd93,-10'd107};
ram[55223] = {9'd96,-10'd104};
ram[55224] = {9'd99,-10'd101};
ram[55225] = {-9'd98,-10'd98};
ram[55226] = {-9'd95,-10'd95};
ram[55227] = {-9'd92,-10'd92};
ram[55228] = {-9'd88,-10'd88};
ram[55229] = {-9'd85,-10'd85};
ram[55230] = {-9'd82,-10'd82};
ram[55231] = {-9'd79,-10'd79};
ram[55232] = {-9'd76,-10'd76};
ram[55233] = {-9'd73,-10'd73};
ram[55234] = {-9'd70,-10'd70};
ram[55235] = {-9'd66,-10'd66};
ram[55236] = {-9'd63,-10'd63};
ram[55237] = {-9'd60,-10'd60};
ram[55238] = {-9'd57,-10'd57};
ram[55239] = {-9'd54,-10'd54};
ram[55240] = {-9'd51,-10'd51};
ram[55241] = {-9'd48,-10'd48};
ram[55242] = {-9'd44,-10'd44};
ram[55243] = {-9'd41,-10'd41};
ram[55244] = {-9'd38,-10'd38};
ram[55245] = {-9'd35,-10'd35};
ram[55246] = {-9'd32,-10'd32};
ram[55247] = {-9'd29,-10'd29};
ram[55248] = {-9'd26,-10'd26};
ram[55249] = {-9'd22,-10'd22};
ram[55250] = {-9'd19,-10'd19};
ram[55251] = {-9'd16,-10'd16};
ram[55252] = {-9'd13,-10'd13};
ram[55253] = {-9'd10,-10'd10};
ram[55254] = {-9'd7,-10'd7};
ram[55255] = {-9'd4,-10'd4};
ram[55256] = {9'd0,10'd0};
ram[55257] = {9'd3,10'd3};
ram[55258] = {9'd6,10'd6};
ram[55259] = {9'd9,10'd9};
ram[55260] = {9'd12,10'd12};
ram[55261] = {9'd15,10'd15};
ram[55262] = {9'd18,10'd18};
ram[55263] = {9'd21,10'd21};
ram[55264] = {9'd25,10'd25};
ram[55265] = {9'd28,10'd28};
ram[55266] = {9'd31,10'd31};
ram[55267] = {9'd34,10'd34};
ram[55268] = {9'd37,10'd37};
ram[55269] = {9'd40,10'd40};
ram[55270] = {9'd43,10'd43};
ram[55271] = {9'd47,10'd47};
ram[55272] = {9'd50,10'd50};
ram[55273] = {9'd53,10'd53};
ram[55274] = {9'd56,10'd56};
ram[55275] = {9'd59,10'd59};
ram[55276] = {9'd62,10'd62};
ram[55277] = {9'd65,10'd65};
ram[55278] = {9'd69,10'd69};
ram[55279] = {9'd72,10'd72};
ram[55280] = {9'd75,10'd75};
ram[55281] = {9'd78,10'd78};
ram[55282] = {9'd81,10'd81};
ram[55283] = {9'd84,10'd84};
ram[55284] = {9'd87,10'd87};
ram[55285] = {9'd91,10'd91};
ram[55286] = {9'd94,10'd94};
ram[55287] = {9'd97,10'd97};
ram[55288] = {-9'd100,10'd100};
ram[55289] = {-9'd97,10'd103};
ram[55290] = {-9'd94,10'd106};
ram[55291] = {-9'd91,10'd109};
ram[55292] = {-9'd88,10'd113};
ram[55293] = {-9'd85,10'd116};
ram[55294] = {-9'd81,10'd119};
ram[55295] = {-9'd78,10'd122};
ram[55296] = {-9'd78,10'd122};
ram[55297] = {-9'd75,10'd125};
ram[55298] = {-9'd72,10'd128};
ram[55299] = {-9'd69,10'd131};
ram[55300] = {-9'd66,10'd135};
ram[55301] = {-9'd63,10'd138};
ram[55302] = {-9'd59,10'd141};
ram[55303] = {-9'd56,10'd144};
ram[55304] = {-9'd53,10'd147};
ram[55305] = {-9'd50,10'd150};
ram[55306] = {-9'd47,10'd153};
ram[55307] = {-9'd44,10'd157};
ram[55308] = {-9'd41,10'd160};
ram[55309] = {-9'd37,10'd163};
ram[55310] = {-9'd34,10'd166};
ram[55311] = {-9'd31,10'd169};
ram[55312] = {-9'd28,10'd172};
ram[55313] = {-9'd25,10'd175};
ram[55314] = {-9'd22,10'd179};
ram[55315] = {-9'd19,10'd182};
ram[55316] = {-9'd15,10'd185};
ram[55317] = {-9'd12,10'd188};
ram[55318] = {-9'd9,10'd191};
ram[55319] = {-9'd6,10'd194};
ram[55320] = {-9'd3,10'd197};
ram[55321] = {9'd0,10'd201};
ram[55322] = {9'd3,10'd204};
ram[55323] = {9'd7,10'd207};
ram[55324] = {9'd10,10'd210};
ram[55325] = {9'd13,10'd213};
ram[55326] = {9'd16,10'd216};
ram[55327] = {9'd19,10'd219};
ram[55328] = {9'd22,10'd223};
ram[55329] = {9'd25,10'd226};
ram[55330] = {9'd29,10'd229};
ram[55331] = {9'd32,10'd232};
ram[55332] = {9'd35,10'd235};
ram[55333] = {9'd38,10'd238};
ram[55334] = {9'd41,10'd241};
ram[55335] = {9'd44,10'd245};
ram[55336] = {9'd47,10'd248};
ram[55337] = {9'd51,10'd251};
ram[55338] = {9'd54,10'd254};
ram[55339] = {9'd57,10'd257};
ram[55340] = {9'd60,10'd260};
ram[55341] = {9'd63,10'd263};
ram[55342] = {9'd66,10'd267};
ram[55343] = {9'd69,10'd270};
ram[55344] = {9'd73,10'd273};
ram[55345] = {9'd76,10'd276};
ram[55346] = {9'd79,10'd279};
ram[55347] = {9'd82,10'd282};
ram[55348] = {9'd85,10'd285};
ram[55349] = {9'd88,10'd289};
ram[55350] = {9'd91,10'd292};
ram[55351] = {9'd95,10'd295};
ram[55352] = {9'd98,10'd298};
ram[55353] = {-9'd99,10'd301};
ram[55354] = {-9'd96,10'd304};
ram[55355] = {-9'd93,10'd307};
ram[55356] = {-9'd90,10'd311};
ram[55357] = {-9'd87,10'd314};
ram[55358] = {-9'd84,10'd317};
ram[55359] = {-9'd81,10'd320};
ram[55360] = {-9'd77,10'd323};
ram[55361] = {-9'd74,10'd326};
ram[55362] = {-9'd71,10'd329};
ram[55363] = {-9'd68,10'd333};
ram[55364] = {-9'd65,10'd336};
ram[55365] = {-9'd62,10'd339};
ram[55366] = {-9'd59,10'd342};
ram[55367] = {-9'd55,10'd345};
ram[55368] = {-9'd52,10'd348};
ram[55369] = {-9'd49,10'd351};
ram[55370] = {-9'd46,10'd354};
ram[55371] = {-9'd43,10'd358};
ram[55372] = {-9'd40,10'd361};
ram[55373] = {-9'd37,10'd364};
ram[55374] = {-9'd33,10'd367};
ram[55375] = {-9'd30,10'd370};
ram[55376] = {-9'd27,10'd373};
ram[55377] = {-9'd24,10'd376};
ram[55378] = {-9'd21,10'd380};
ram[55379] = {-9'd18,10'd383};
ram[55380] = {-9'd15,10'd386};
ram[55381] = {-9'd11,10'd389};
ram[55382] = {-9'd8,10'd392};
ram[55383] = {-9'd5,10'd395};
ram[55384] = {-9'd2,10'd398};
ram[55385] = {9'd1,-10'd399};
ram[55386] = {9'd4,-10'd396};
ram[55387] = {9'd7,-10'd393};
ram[55388] = {9'd10,-10'd390};
ram[55389] = {9'd14,-10'd387};
ram[55390] = {9'd17,-10'd384};
ram[55391] = {9'd20,-10'd381};
ram[55392] = {9'd23,-10'd377};
ram[55393] = {9'd26,-10'd374};
ram[55394] = {9'd29,-10'd371};
ram[55395] = {9'd32,-10'd368};
ram[55396] = {9'd36,-10'd365};
ram[55397] = {9'd39,-10'd362};
ram[55398] = {9'd42,-10'd359};
ram[55399] = {9'd45,-10'd355};
ram[55400] = {9'd48,-10'd352};
ram[55401] = {9'd51,-10'd349};
ram[55402] = {9'd54,-10'd346};
ram[55403] = {9'd58,-10'd343};
ram[55404] = {9'd61,-10'd340};
ram[55405] = {9'd64,-10'd337};
ram[55406] = {9'd67,-10'd334};
ram[55407] = {9'd70,-10'd330};
ram[55408] = {9'd73,-10'd327};
ram[55409] = {9'd76,-10'd324};
ram[55410] = {9'd80,-10'd321};
ram[55411] = {9'd83,-10'd318};
ram[55412] = {9'd86,-10'd315};
ram[55413] = {9'd89,-10'd312};
ram[55414] = {9'd92,-10'd308};
ram[55415] = {9'd95,-10'd305};
ram[55416] = {9'd98,-10'd302};
ram[55417] = {-9'd99,-10'd299};
ram[55418] = {-9'd96,-10'd296};
ram[55419] = {-9'd92,-10'd293};
ram[55420] = {-9'd89,-10'd290};
ram[55421] = {-9'd86,-10'd286};
ram[55422] = {-9'd83,-10'd283};
ram[55423] = {-9'd80,-10'd280};
ram[55424] = {-9'd80,-10'd280};
ram[55425] = {-9'd77,-10'd277};
ram[55426] = {-9'd74,-10'd274};
ram[55427] = {-9'd70,-10'd271};
ram[55428] = {-9'd67,-10'd268};
ram[55429] = {-9'd64,-10'd264};
ram[55430] = {-9'd61,-10'd261};
ram[55431] = {-9'd58,-10'd258};
ram[55432] = {-9'd55,-10'd255};
ram[55433] = {-9'd52,-10'd252};
ram[55434] = {-9'd48,-10'd249};
ram[55435] = {-9'd45,-10'd246};
ram[55436] = {-9'd42,-10'd242};
ram[55437] = {-9'd39,-10'd239};
ram[55438] = {-9'd36,-10'd236};
ram[55439] = {-9'd33,-10'd233};
ram[55440] = {-9'd30,-10'd230};
ram[55441] = {-9'd26,-10'd227};
ram[55442] = {-9'd23,-10'd224};
ram[55443] = {-9'd20,-10'd220};
ram[55444] = {-9'd17,-10'd217};
ram[55445] = {-9'd14,-10'd214};
ram[55446] = {-9'd11,-10'd211};
ram[55447] = {-9'd8,-10'd208};
ram[55448] = {-9'd4,-10'd205};
ram[55449] = {-9'd1,-10'd202};
ram[55450] = {9'd2,-10'd198};
ram[55451] = {9'd5,-10'd195};
ram[55452] = {9'd8,-10'd192};
ram[55453] = {9'd11,-10'd189};
ram[55454] = {9'd14,-10'd186};
ram[55455] = {9'd18,-10'd183};
ram[55456] = {9'd21,-10'd180};
ram[55457] = {9'd24,-10'd176};
ram[55458] = {9'd27,-10'd173};
ram[55459] = {9'd30,-10'd170};
ram[55460] = {9'd33,-10'd167};
ram[55461] = {9'd36,-10'd164};
ram[55462] = {9'd40,-10'd161};
ram[55463] = {9'd43,-10'd158};
ram[55464] = {9'd46,-10'd154};
ram[55465] = {9'd49,-10'd151};
ram[55466] = {9'd52,-10'd148};
ram[55467] = {9'd55,-10'd145};
ram[55468] = {9'd58,-10'd142};
ram[55469] = {9'd62,-10'd139};
ram[55470] = {9'd65,-10'd136};
ram[55471] = {9'd68,-10'd132};
ram[55472] = {9'd71,-10'd129};
ram[55473] = {9'd74,-10'd126};
ram[55474] = {9'd77,-10'd123};
ram[55475] = {9'd80,-10'd120};
ram[55476] = {9'd84,-10'd117};
ram[55477] = {9'd87,-10'd114};
ram[55478] = {9'd90,-10'd110};
ram[55479] = {9'd93,-10'd107};
ram[55480] = {9'd96,-10'd104};
ram[55481] = {9'd99,-10'd101};
ram[55482] = {-9'd98,-10'd98};
ram[55483] = {-9'd95,-10'd95};
ram[55484] = {-9'd92,-10'd92};
ram[55485] = {-9'd88,-10'd88};
ram[55486] = {-9'd85,-10'd85};
ram[55487] = {-9'd82,-10'd82};
ram[55488] = {-9'd79,-10'd79};
ram[55489] = {-9'd76,-10'd76};
ram[55490] = {-9'd73,-10'd73};
ram[55491] = {-9'd70,-10'd70};
ram[55492] = {-9'd66,-10'd66};
ram[55493] = {-9'd63,-10'd63};
ram[55494] = {-9'd60,-10'd60};
ram[55495] = {-9'd57,-10'd57};
ram[55496] = {-9'd54,-10'd54};
ram[55497] = {-9'd51,-10'd51};
ram[55498] = {-9'd48,-10'd48};
ram[55499] = {-9'd44,-10'd44};
ram[55500] = {-9'd41,-10'd41};
ram[55501] = {-9'd38,-10'd38};
ram[55502] = {-9'd35,-10'd35};
ram[55503] = {-9'd32,-10'd32};
ram[55504] = {-9'd29,-10'd29};
ram[55505] = {-9'd26,-10'd26};
ram[55506] = {-9'd22,-10'd22};
ram[55507] = {-9'd19,-10'd19};
ram[55508] = {-9'd16,-10'd16};
ram[55509] = {-9'd13,-10'd13};
ram[55510] = {-9'd10,-10'd10};
ram[55511] = {-9'd7,-10'd7};
ram[55512] = {-9'd4,-10'd4};
ram[55513] = {9'd0,10'd0};
ram[55514] = {9'd3,10'd3};
ram[55515] = {9'd6,10'd6};
ram[55516] = {9'd9,10'd9};
ram[55517] = {9'd12,10'd12};
ram[55518] = {9'd15,10'd15};
ram[55519] = {9'd18,10'd18};
ram[55520] = {9'd21,10'd21};
ram[55521] = {9'd25,10'd25};
ram[55522] = {9'd28,10'd28};
ram[55523] = {9'd31,10'd31};
ram[55524] = {9'd34,10'd34};
ram[55525] = {9'd37,10'd37};
ram[55526] = {9'd40,10'd40};
ram[55527] = {9'd43,10'd43};
ram[55528] = {9'd47,10'd47};
ram[55529] = {9'd50,10'd50};
ram[55530] = {9'd53,10'd53};
ram[55531] = {9'd56,10'd56};
ram[55532] = {9'd59,10'd59};
ram[55533] = {9'd62,10'd62};
ram[55534] = {9'd65,10'd65};
ram[55535] = {9'd69,10'd69};
ram[55536] = {9'd72,10'd72};
ram[55537] = {9'd75,10'd75};
ram[55538] = {9'd78,10'd78};
ram[55539] = {9'd81,10'd81};
ram[55540] = {9'd84,10'd84};
ram[55541] = {9'd87,10'd87};
ram[55542] = {9'd91,10'd91};
ram[55543] = {9'd94,10'd94};
ram[55544] = {9'd97,10'd97};
ram[55545] = {-9'd100,10'd100};
ram[55546] = {-9'd97,10'd103};
ram[55547] = {-9'd94,10'd106};
ram[55548] = {-9'd91,10'd109};
ram[55549] = {-9'd88,10'd113};
ram[55550] = {-9'd85,10'd116};
ram[55551] = {-9'd81,10'd119};
ram[55552] = {-9'd81,10'd119};
ram[55553] = {-9'd78,10'd122};
ram[55554] = {-9'd75,10'd125};
ram[55555] = {-9'd72,10'd128};
ram[55556] = {-9'd69,10'd131};
ram[55557] = {-9'd66,10'd135};
ram[55558] = {-9'd63,10'd138};
ram[55559] = {-9'd59,10'd141};
ram[55560] = {-9'd56,10'd144};
ram[55561] = {-9'd53,10'd147};
ram[55562] = {-9'd50,10'd150};
ram[55563] = {-9'd47,10'd153};
ram[55564] = {-9'd44,10'd157};
ram[55565] = {-9'd41,10'd160};
ram[55566] = {-9'd37,10'd163};
ram[55567] = {-9'd34,10'd166};
ram[55568] = {-9'd31,10'd169};
ram[55569] = {-9'd28,10'd172};
ram[55570] = {-9'd25,10'd175};
ram[55571] = {-9'd22,10'd179};
ram[55572] = {-9'd19,10'd182};
ram[55573] = {-9'd15,10'd185};
ram[55574] = {-9'd12,10'd188};
ram[55575] = {-9'd9,10'd191};
ram[55576] = {-9'd6,10'd194};
ram[55577] = {-9'd3,10'd197};
ram[55578] = {9'd0,10'd201};
ram[55579] = {9'd3,10'd204};
ram[55580] = {9'd7,10'd207};
ram[55581] = {9'd10,10'd210};
ram[55582] = {9'd13,10'd213};
ram[55583] = {9'd16,10'd216};
ram[55584] = {9'd19,10'd219};
ram[55585] = {9'd22,10'd223};
ram[55586] = {9'd25,10'd226};
ram[55587] = {9'd29,10'd229};
ram[55588] = {9'd32,10'd232};
ram[55589] = {9'd35,10'd235};
ram[55590] = {9'd38,10'd238};
ram[55591] = {9'd41,10'd241};
ram[55592] = {9'd44,10'd245};
ram[55593] = {9'd47,10'd248};
ram[55594] = {9'd51,10'd251};
ram[55595] = {9'd54,10'd254};
ram[55596] = {9'd57,10'd257};
ram[55597] = {9'd60,10'd260};
ram[55598] = {9'd63,10'd263};
ram[55599] = {9'd66,10'd267};
ram[55600] = {9'd69,10'd270};
ram[55601] = {9'd73,10'd273};
ram[55602] = {9'd76,10'd276};
ram[55603] = {9'd79,10'd279};
ram[55604] = {9'd82,10'd282};
ram[55605] = {9'd85,10'd285};
ram[55606] = {9'd88,10'd289};
ram[55607] = {9'd91,10'd292};
ram[55608] = {9'd95,10'd295};
ram[55609] = {9'd98,10'd298};
ram[55610] = {-9'd99,10'd301};
ram[55611] = {-9'd96,10'd304};
ram[55612] = {-9'd93,10'd307};
ram[55613] = {-9'd90,10'd311};
ram[55614] = {-9'd87,10'd314};
ram[55615] = {-9'd84,10'd317};
ram[55616] = {-9'd81,10'd320};
ram[55617] = {-9'd77,10'd323};
ram[55618] = {-9'd74,10'd326};
ram[55619] = {-9'd71,10'd329};
ram[55620] = {-9'd68,10'd333};
ram[55621] = {-9'd65,10'd336};
ram[55622] = {-9'd62,10'd339};
ram[55623] = {-9'd59,10'd342};
ram[55624] = {-9'd55,10'd345};
ram[55625] = {-9'd52,10'd348};
ram[55626] = {-9'd49,10'd351};
ram[55627] = {-9'd46,10'd354};
ram[55628] = {-9'd43,10'd358};
ram[55629] = {-9'd40,10'd361};
ram[55630] = {-9'd37,10'd364};
ram[55631] = {-9'd33,10'd367};
ram[55632] = {-9'd30,10'd370};
ram[55633] = {-9'd27,10'd373};
ram[55634] = {-9'd24,10'd376};
ram[55635] = {-9'd21,10'd380};
ram[55636] = {-9'd18,10'd383};
ram[55637] = {-9'd15,10'd386};
ram[55638] = {-9'd11,10'd389};
ram[55639] = {-9'd8,10'd392};
ram[55640] = {-9'd5,10'd395};
ram[55641] = {-9'd2,10'd398};
ram[55642] = {9'd1,-10'd399};
ram[55643] = {9'd4,-10'd396};
ram[55644] = {9'd7,-10'd393};
ram[55645] = {9'd10,-10'd390};
ram[55646] = {9'd14,-10'd387};
ram[55647] = {9'd17,-10'd384};
ram[55648] = {9'd20,-10'd381};
ram[55649] = {9'd23,-10'd377};
ram[55650] = {9'd26,-10'd374};
ram[55651] = {9'd29,-10'd371};
ram[55652] = {9'd32,-10'd368};
ram[55653] = {9'd36,-10'd365};
ram[55654] = {9'd39,-10'd362};
ram[55655] = {9'd42,-10'd359};
ram[55656] = {9'd45,-10'd355};
ram[55657] = {9'd48,-10'd352};
ram[55658] = {9'd51,-10'd349};
ram[55659] = {9'd54,-10'd346};
ram[55660] = {9'd58,-10'd343};
ram[55661] = {9'd61,-10'd340};
ram[55662] = {9'd64,-10'd337};
ram[55663] = {9'd67,-10'd334};
ram[55664] = {9'd70,-10'd330};
ram[55665] = {9'd73,-10'd327};
ram[55666] = {9'd76,-10'd324};
ram[55667] = {9'd80,-10'd321};
ram[55668] = {9'd83,-10'd318};
ram[55669] = {9'd86,-10'd315};
ram[55670] = {9'd89,-10'd312};
ram[55671] = {9'd92,-10'd308};
ram[55672] = {9'd95,-10'd305};
ram[55673] = {9'd98,-10'd302};
ram[55674] = {-9'd99,-10'd299};
ram[55675] = {-9'd96,-10'd296};
ram[55676] = {-9'd92,-10'd293};
ram[55677] = {-9'd89,-10'd290};
ram[55678] = {-9'd86,-10'd286};
ram[55679] = {-9'd83,-10'd283};
ram[55680] = {-9'd83,-10'd283};
ram[55681] = {-9'd80,-10'd280};
ram[55682] = {-9'd77,-10'd277};
ram[55683] = {-9'd74,-10'd274};
ram[55684] = {-9'd70,-10'd271};
ram[55685] = {-9'd67,-10'd268};
ram[55686] = {-9'd64,-10'd264};
ram[55687] = {-9'd61,-10'd261};
ram[55688] = {-9'd58,-10'd258};
ram[55689] = {-9'd55,-10'd255};
ram[55690] = {-9'd52,-10'd252};
ram[55691] = {-9'd48,-10'd249};
ram[55692] = {-9'd45,-10'd246};
ram[55693] = {-9'd42,-10'd242};
ram[55694] = {-9'd39,-10'd239};
ram[55695] = {-9'd36,-10'd236};
ram[55696] = {-9'd33,-10'd233};
ram[55697] = {-9'd30,-10'd230};
ram[55698] = {-9'd26,-10'd227};
ram[55699] = {-9'd23,-10'd224};
ram[55700] = {-9'd20,-10'd220};
ram[55701] = {-9'd17,-10'd217};
ram[55702] = {-9'd14,-10'd214};
ram[55703] = {-9'd11,-10'd211};
ram[55704] = {-9'd8,-10'd208};
ram[55705] = {-9'd4,-10'd205};
ram[55706] = {-9'd1,-10'd202};
ram[55707] = {9'd2,-10'd198};
ram[55708] = {9'd5,-10'd195};
ram[55709] = {9'd8,-10'd192};
ram[55710] = {9'd11,-10'd189};
ram[55711] = {9'd14,-10'd186};
ram[55712] = {9'd18,-10'd183};
ram[55713] = {9'd21,-10'd180};
ram[55714] = {9'd24,-10'd176};
ram[55715] = {9'd27,-10'd173};
ram[55716] = {9'd30,-10'd170};
ram[55717] = {9'd33,-10'd167};
ram[55718] = {9'd36,-10'd164};
ram[55719] = {9'd40,-10'd161};
ram[55720] = {9'd43,-10'd158};
ram[55721] = {9'd46,-10'd154};
ram[55722] = {9'd49,-10'd151};
ram[55723] = {9'd52,-10'd148};
ram[55724] = {9'd55,-10'd145};
ram[55725] = {9'd58,-10'd142};
ram[55726] = {9'd62,-10'd139};
ram[55727] = {9'd65,-10'd136};
ram[55728] = {9'd68,-10'd132};
ram[55729] = {9'd71,-10'd129};
ram[55730] = {9'd74,-10'd126};
ram[55731] = {9'd77,-10'd123};
ram[55732] = {9'd80,-10'd120};
ram[55733] = {9'd84,-10'd117};
ram[55734] = {9'd87,-10'd114};
ram[55735] = {9'd90,-10'd110};
ram[55736] = {9'd93,-10'd107};
ram[55737] = {9'd96,-10'd104};
ram[55738] = {9'd99,-10'd101};
ram[55739] = {-9'd98,-10'd98};
ram[55740] = {-9'd95,-10'd95};
ram[55741] = {-9'd92,-10'd92};
ram[55742] = {-9'd88,-10'd88};
ram[55743] = {-9'd85,-10'd85};
ram[55744] = {-9'd82,-10'd82};
ram[55745] = {-9'd79,-10'd79};
ram[55746] = {-9'd76,-10'd76};
ram[55747] = {-9'd73,-10'd73};
ram[55748] = {-9'd70,-10'd70};
ram[55749] = {-9'd66,-10'd66};
ram[55750] = {-9'd63,-10'd63};
ram[55751] = {-9'd60,-10'd60};
ram[55752] = {-9'd57,-10'd57};
ram[55753] = {-9'd54,-10'd54};
ram[55754] = {-9'd51,-10'd51};
ram[55755] = {-9'd48,-10'd48};
ram[55756] = {-9'd44,-10'd44};
ram[55757] = {-9'd41,-10'd41};
ram[55758] = {-9'd38,-10'd38};
ram[55759] = {-9'd35,-10'd35};
ram[55760] = {-9'd32,-10'd32};
ram[55761] = {-9'd29,-10'd29};
ram[55762] = {-9'd26,-10'd26};
ram[55763] = {-9'd22,-10'd22};
ram[55764] = {-9'd19,-10'd19};
ram[55765] = {-9'd16,-10'd16};
ram[55766] = {-9'd13,-10'd13};
ram[55767] = {-9'd10,-10'd10};
ram[55768] = {-9'd7,-10'd7};
ram[55769] = {-9'd4,-10'd4};
ram[55770] = {9'd0,10'd0};
ram[55771] = {9'd3,10'd3};
ram[55772] = {9'd6,10'd6};
ram[55773] = {9'd9,10'd9};
ram[55774] = {9'd12,10'd12};
ram[55775] = {9'd15,10'd15};
ram[55776] = {9'd18,10'd18};
ram[55777] = {9'd21,10'd21};
ram[55778] = {9'd25,10'd25};
ram[55779] = {9'd28,10'd28};
ram[55780] = {9'd31,10'd31};
ram[55781] = {9'd34,10'd34};
ram[55782] = {9'd37,10'd37};
ram[55783] = {9'd40,10'd40};
ram[55784] = {9'd43,10'd43};
ram[55785] = {9'd47,10'd47};
ram[55786] = {9'd50,10'd50};
ram[55787] = {9'd53,10'd53};
ram[55788] = {9'd56,10'd56};
ram[55789] = {9'd59,10'd59};
ram[55790] = {9'd62,10'd62};
ram[55791] = {9'd65,10'd65};
ram[55792] = {9'd69,10'd69};
ram[55793] = {9'd72,10'd72};
ram[55794] = {9'd75,10'd75};
ram[55795] = {9'd78,10'd78};
ram[55796] = {9'd81,10'd81};
ram[55797] = {9'd84,10'd84};
ram[55798] = {9'd87,10'd87};
ram[55799] = {9'd91,10'd91};
ram[55800] = {9'd94,10'd94};
ram[55801] = {9'd97,10'd97};
ram[55802] = {-9'd100,10'd100};
ram[55803] = {-9'd97,10'd103};
ram[55804] = {-9'd94,10'd106};
ram[55805] = {-9'd91,10'd109};
ram[55806] = {-9'd88,10'd113};
ram[55807] = {-9'd85,10'd116};
ram[55808] = {-9'd85,10'd116};
ram[55809] = {-9'd81,10'd119};
ram[55810] = {-9'd78,10'd122};
ram[55811] = {-9'd75,10'd125};
ram[55812] = {-9'd72,10'd128};
ram[55813] = {-9'd69,10'd131};
ram[55814] = {-9'd66,10'd135};
ram[55815] = {-9'd63,10'd138};
ram[55816] = {-9'd59,10'd141};
ram[55817] = {-9'd56,10'd144};
ram[55818] = {-9'd53,10'd147};
ram[55819] = {-9'd50,10'd150};
ram[55820] = {-9'd47,10'd153};
ram[55821] = {-9'd44,10'd157};
ram[55822] = {-9'd41,10'd160};
ram[55823] = {-9'd37,10'd163};
ram[55824] = {-9'd34,10'd166};
ram[55825] = {-9'd31,10'd169};
ram[55826] = {-9'd28,10'd172};
ram[55827] = {-9'd25,10'd175};
ram[55828] = {-9'd22,10'd179};
ram[55829] = {-9'd19,10'd182};
ram[55830] = {-9'd15,10'd185};
ram[55831] = {-9'd12,10'd188};
ram[55832] = {-9'd9,10'd191};
ram[55833] = {-9'd6,10'd194};
ram[55834] = {-9'd3,10'd197};
ram[55835] = {9'd0,10'd201};
ram[55836] = {9'd3,10'd204};
ram[55837] = {9'd7,10'd207};
ram[55838] = {9'd10,10'd210};
ram[55839] = {9'd13,10'd213};
ram[55840] = {9'd16,10'd216};
ram[55841] = {9'd19,10'd219};
ram[55842] = {9'd22,10'd223};
ram[55843] = {9'd25,10'd226};
ram[55844] = {9'd29,10'd229};
ram[55845] = {9'd32,10'd232};
ram[55846] = {9'd35,10'd235};
ram[55847] = {9'd38,10'd238};
ram[55848] = {9'd41,10'd241};
ram[55849] = {9'd44,10'd245};
ram[55850] = {9'd47,10'd248};
ram[55851] = {9'd51,10'd251};
ram[55852] = {9'd54,10'd254};
ram[55853] = {9'd57,10'd257};
ram[55854] = {9'd60,10'd260};
ram[55855] = {9'd63,10'd263};
ram[55856] = {9'd66,10'd267};
ram[55857] = {9'd69,10'd270};
ram[55858] = {9'd73,10'd273};
ram[55859] = {9'd76,10'd276};
ram[55860] = {9'd79,10'd279};
ram[55861] = {9'd82,10'd282};
ram[55862] = {9'd85,10'd285};
ram[55863] = {9'd88,10'd289};
ram[55864] = {9'd91,10'd292};
ram[55865] = {9'd95,10'd295};
ram[55866] = {9'd98,10'd298};
ram[55867] = {-9'd99,10'd301};
ram[55868] = {-9'd96,10'd304};
ram[55869] = {-9'd93,10'd307};
ram[55870] = {-9'd90,10'd311};
ram[55871] = {-9'd87,10'd314};
ram[55872] = {-9'd84,10'd317};
ram[55873] = {-9'd81,10'd320};
ram[55874] = {-9'd77,10'd323};
ram[55875] = {-9'd74,10'd326};
ram[55876] = {-9'd71,10'd329};
ram[55877] = {-9'd68,10'd333};
ram[55878] = {-9'd65,10'd336};
ram[55879] = {-9'd62,10'd339};
ram[55880] = {-9'd59,10'd342};
ram[55881] = {-9'd55,10'd345};
ram[55882] = {-9'd52,10'd348};
ram[55883] = {-9'd49,10'd351};
ram[55884] = {-9'd46,10'd354};
ram[55885] = {-9'd43,10'd358};
ram[55886] = {-9'd40,10'd361};
ram[55887] = {-9'd37,10'd364};
ram[55888] = {-9'd33,10'd367};
ram[55889] = {-9'd30,10'd370};
ram[55890] = {-9'd27,10'd373};
ram[55891] = {-9'd24,10'd376};
ram[55892] = {-9'd21,10'd380};
ram[55893] = {-9'd18,10'd383};
ram[55894] = {-9'd15,10'd386};
ram[55895] = {-9'd11,10'd389};
ram[55896] = {-9'd8,10'd392};
ram[55897] = {-9'd5,10'd395};
ram[55898] = {-9'd2,10'd398};
ram[55899] = {9'd1,-10'd399};
ram[55900] = {9'd4,-10'd396};
ram[55901] = {9'd7,-10'd393};
ram[55902] = {9'd10,-10'd390};
ram[55903] = {9'd14,-10'd387};
ram[55904] = {9'd17,-10'd384};
ram[55905] = {9'd20,-10'd381};
ram[55906] = {9'd23,-10'd377};
ram[55907] = {9'd26,-10'd374};
ram[55908] = {9'd29,-10'd371};
ram[55909] = {9'd32,-10'd368};
ram[55910] = {9'd36,-10'd365};
ram[55911] = {9'd39,-10'd362};
ram[55912] = {9'd42,-10'd359};
ram[55913] = {9'd45,-10'd355};
ram[55914] = {9'd48,-10'd352};
ram[55915] = {9'd51,-10'd349};
ram[55916] = {9'd54,-10'd346};
ram[55917] = {9'd58,-10'd343};
ram[55918] = {9'd61,-10'd340};
ram[55919] = {9'd64,-10'd337};
ram[55920] = {9'd67,-10'd334};
ram[55921] = {9'd70,-10'd330};
ram[55922] = {9'd73,-10'd327};
ram[55923] = {9'd76,-10'd324};
ram[55924] = {9'd80,-10'd321};
ram[55925] = {9'd83,-10'd318};
ram[55926] = {9'd86,-10'd315};
ram[55927] = {9'd89,-10'd312};
ram[55928] = {9'd92,-10'd308};
ram[55929] = {9'd95,-10'd305};
ram[55930] = {9'd98,-10'd302};
ram[55931] = {-9'd99,-10'd299};
ram[55932] = {-9'd96,-10'd296};
ram[55933] = {-9'd92,-10'd293};
ram[55934] = {-9'd89,-10'd290};
ram[55935] = {-9'd86,-10'd286};
ram[55936] = {-9'd86,-10'd286};
ram[55937] = {-9'd83,-10'd283};
ram[55938] = {-9'd80,-10'd280};
ram[55939] = {-9'd77,-10'd277};
ram[55940] = {-9'd74,-10'd274};
ram[55941] = {-9'd70,-10'd271};
ram[55942] = {-9'd67,-10'd268};
ram[55943] = {-9'd64,-10'd264};
ram[55944] = {-9'd61,-10'd261};
ram[55945] = {-9'd58,-10'd258};
ram[55946] = {-9'd55,-10'd255};
ram[55947] = {-9'd52,-10'd252};
ram[55948] = {-9'd48,-10'd249};
ram[55949] = {-9'd45,-10'd246};
ram[55950] = {-9'd42,-10'd242};
ram[55951] = {-9'd39,-10'd239};
ram[55952] = {-9'd36,-10'd236};
ram[55953] = {-9'd33,-10'd233};
ram[55954] = {-9'd30,-10'd230};
ram[55955] = {-9'd26,-10'd227};
ram[55956] = {-9'd23,-10'd224};
ram[55957] = {-9'd20,-10'd220};
ram[55958] = {-9'd17,-10'd217};
ram[55959] = {-9'd14,-10'd214};
ram[55960] = {-9'd11,-10'd211};
ram[55961] = {-9'd8,-10'd208};
ram[55962] = {-9'd4,-10'd205};
ram[55963] = {-9'd1,-10'd202};
ram[55964] = {9'd2,-10'd198};
ram[55965] = {9'd5,-10'd195};
ram[55966] = {9'd8,-10'd192};
ram[55967] = {9'd11,-10'd189};
ram[55968] = {9'd14,-10'd186};
ram[55969] = {9'd18,-10'd183};
ram[55970] = {9'd21,-10'd180};
ram[55971] = {9'd24,-10'd176};
ram[55972] = {9'd27,-10'd173};
ram[55973] = {9'd30,-10'd170};
ram[55974] = {9'd33,-10'd167};
ram[55975] = {9'd36,-10'd164};
ram[55976] = {9'd40,-10'd161};
ram[55977] = {9'd43,-10'd158};
ram[55978] = {9'd46,-10'd154};
ram[55979] = {9'd49,-10'd151};
ram[55980] = {9'd52,-10'd148};
ram[55981] = {9'd55,-10'd145};
ram[55982] = {9'd58,-10'd142};
ram[55983] = {9'd62,-10'd139};
ram[55984] = {9'd65,-10'd136};
ram[55985] = {9'd68,-10'd132};
ram[55986] = {9'd71,-10'd129};
ram[55987] = {9'd74,-10'd126};
ram[55988] = {9'd77,-10'd123};
ram[55989] = {9'd80,-10'd120};
ram[55990] = {9'd84,-10'd117};
ram[55991] = {9'd87,-10'd114};
ram[55992] = {9'd90,-10'd110};
ram[55993] = {9'd93,-10'd107};
ram[55994] = {9'd96,-10'd104};
ram[55995] = {9'd99,-10'd101};
ram[55996] = {-9'd98,-10'd98};
ram[55997] = {-9'd95,-10'd95};
ram[55998] = {-9'd92,-10'd92};
ram[55999] = {-9'd88,-10'd88};
ram[56000] = {-9'd85,-10'd85};
ram[56001] = {-9'd82,-10'd82};
ram[56002] = {-9'd79,-10'd79};
ram[56003] = {-9'd76,-10'd76};
ram[56004] = {-9'd73,-10'd73};
ram[56005] = {-9'd70,-10'd70};
ram[56006] = {-9'd66,-10'd66};
ram[56007] = {-9'd63,-10'd63};
ram[56008] = {-9'd60,-10'd60};
ram[56009] = {-9'd57,-10'd57};
ram[56010] = {-9'd54,-10'd54};
ram[56011] = {-9'd51,-10'd51};
ram[56012] = {-9'd48,-10'd48};
ram[56013] = {-9'd44,-10'd44};
ram[56014] = {-9'd41,-10'd41};
ram[56015] = {-9'd38,-10'd38};
ram[56016] = {-9'd35,-10'd35};
ram[56017] = {-9'd32,-10'd32};
ram[56018] = {-9'd29,-10'd29};
ram[56019] = {-9'd26,-10'd26};
ram[56020] = {-9'd22,-10'd22};
ram[56021] = {-9'd19,-10'd19};
ram[56022] = {-9'd16,-10'd16};
ram[56023] = {-9'd13,-10'd13};
ram[56024] = {-9'd10,-10'd10};
ram[56025] = {-9'd7,-10'd7};
ram[56026] = {-9'd4,-10'd4};
ram[56027] = {9'd0,10'd0};
ram[56028] = {9'd3,10'd3};
ram[56029] = {9'd6,10'd6};
ram[56030] = {9'd9,10'd9};
ram[56031] = {9'd12,10'd12};
ram[56032] = {9'd15,10'd15};
ram[56033] = {9'd18,10'd18};
ram[56034] = {9'd21,10'd21};
ram[56035] = {9'd25,10'd25};
ram[56036] = {9'd28,10'd28};
ram[56037] = {9'd31,10'd31};
ram[56038] = {9'd34,10'd34};
ram[56039] = {9'd37,10'd37};
ram[56040] = {9'd40,10'd40};
ram[56041] = {9'd43,10'd43};
ram[56042] = {9'd47,10'd47};
ram[56043] = {9'd50,10'd50};
ram[56044] = {9'd53,10'd53};
ram[56045] = {9'd56,10'd56};
ram[56046] = {9'd59,10'd59};
ram[56047] = {9'd62,10'd62};
ram[56048] = {9'd65,10'd65};
ram[56049] = {9'd69,10'd69};
ram[56050] = {9'd72,10'd72};
ram[56051] = {9'd75,10'd75};
ram[56052] = {9'd78,10'd78};
ram[56053] = {9'd81,10'd81};
ram[56054] = {9'd84,10'd84};
ram[56055] = {9'd87,10'd87};
ram[56056] = {9'd91,10'd91};
ram[56057] = {9'd94,10'd94};
ram[56058] = {9'd97,10'd97};
ram[56059] = {-9'd100,10'd100};
ram[56060] = {-9'd97,10'd103};
ram[56061] = {-9'd94,10'd106};
ram[56062] = {-9'd91,10'd109};
ram[56063] = {-9'd88,10'd113};
ram[56064] = {-9'd88,10'd113};
ram[56065] = {-9'd85,10'd116};
ram[56066] = {-9'd81,10'd119};
ram[56067] = {-9'd78,10'd122};
ram[56068] = {-9'd75,10'd125};
ram[56069] = {-9'd72,10'd128};
ram[56070] = {-9'd69,10'd131};
ram[56071] = {-9'd66,10'd135};
ram[56072] = {-9'd63,10'd138};
ram[56073] = {-9'd59,10'd141};
ram[56074] = {-9'd56,10'd144};
ram[56075] = {-9'd53,10'd147};
ram[56076] = {-9'd50,10'd150};
ram[56077] = {-9'd47,10'd153};
ram[56078] = {-9'd44,10'd157};
ram[56079] = {-9'd41,10'd160};
ram[56080] = {-9'd37,10'd163};
ram[56081] = {-9'd34,10'd166};
ram[56082] = {-9'd31,10'd169};
ram[56083] = {-9'd28,10'd172};
ram[56084] = {-9'd25,10'd175};
ram[56085] = {-9'd22,10'd179};
ram[56086] = {-9'd19,10'd182};
ram[56087] = {-9'd15,10'd185};
ram[56088] = {-9'd12,10'd188};
ram[56089] = {-9'd9,10'd191};
ram[56090] = {-9'd6,10'd194};
ram[56091] = {-9'd3,10'd197};
ram[56092] = {9'd0,10'd201};
ram[56093] = {9'd3,10'd204};
ram[56094] = {9'd7,10'd207};
ram[56095] = {9'd10,10'd210};
ram[56096] = {9'd13,10'd213};
ram[56097] = {9'd16,10'd216};
ram[56098] = {9'd19,10'd219};
ram[56099] = {9'd22,10'd223};
ram[56100] = {9'd25,10'd226};
ram[56101] = {9'd29,10'd229};
ram[56102] = {9'd32,10'd232};
ram[56103] = {9'd35,10'd235};
ram[56104] = {9'd38,10'd238};
ram[56105] = {9'd41,10'd241};
ram[56106] = {9'd44,10'd245};
ram[56107] = {9'd47,10'd248};
ram[56108] = {9'd51,10'd251};
ram[56109] = {9'd54,10'd254};
ram[56110] = {9'd57,10'd257};
ram[56111] = {9'd60,10'd260};
ram[56112] = {9'd63,10'd263};
ram[56113] = {9'd66,10'd267};
ram[56114] = {9'd69,10'd270};
ram[56115] = {9'd73,10'd273};
ram[56116] = {9'd76,10'd276};
ram[56117] = {9'd79,10'd279};
ram[56118] = {9'd82,10'd282};
ram[56119] = {9'd85,10'd285};
ram[56120] = {9'd88,10'd289};
ram[56121] = {9'd91,10'd292};
ram[56122] = {9'd95,10'd295};
ram[56123] = {9'd98,10'd298};
ram[56124] = {-9'd99,10'd301};
ram[56125] = {-9'd96,10'd304};
ram[56126] = {-9'd93,10'd307};
ram[56127] = {-9'd90,10'd311};
ram[56128] = {-9'd87,10'd314};
ram[56129] = {-9'd84,10'd317};
ram[56130] = {-9'd81,10'd320};
ram[56131] = {-9'd77,10'd323};
ram[56132] = {-9'd74,10'd326};
ram[56133] = {-9'd71,10'd329};
ram[56134] = {-9'd68,10'd333};
ram[56135] = {-9'd65,10'd336};
ram[56136] = {-9'd62,10'd339};
ram[56137] = {-9'd59,10'd342};
ram[56138] = {-9'd55,10'd345};
ram[56139] = {-9'd52,10'd348};
ram[56140] = {-9'd49,10'd351};
ram[56141] = {-9'd46,10'd354};
ram[56142] = {-9'd43,10'd358};
ram[56143] = {-9'd40,10'd361};
ram[56144] = {-9'd37,10'd364};
ram[56145] = {-9'd33,10'd367};
ram[56146] = {-9'd30,10'd370};
ram[56147] = {-9'd27,10'd373};
ram[56148] = {-9'd24,10'd376};
ram[56149] = {-9'd21,10'd380};
ram[56150] = {-9'd18,10'd383};
ram[56151] = {-9'd15,10'd386};
ram[56152] = {-9'd11,10'd389};
ram[56153] = {-9'd8,10'd392};
ram[56154] = {-9'd5,10'd395};
ram[56155] = {-9'd2,10'd398};
ram[56156] = {9'd1,-10'd399};
ram[56157] = {9'd4,-10'd396};
ram[56158] = {9'd7,-10'd393};
ram[56159] = {9'd10,-10'd390};
ram[56160] = {9'd14,-10'd387};
ram[56161] = {9'd17,-10'd384};
ram[56162] = {9'd20,-10'd381};
ram[56163] = {9'd23,-10'd377};
ram[56164] = {9'd26,-10'd374};
ram[56165] = {9'd29,-10'd371};
ram[56166] = {9'd32,-10'd368};
ram[56167] = {9'd36,-10'd365};
ram[56168] = {9'd39,-10'd362};
ram[56169] = {9'd42,-10'd359};
ram[56170] = {9'd45,-10'd355};
ram[56171] = {9'd48,-10'd352};
ram[56172] = {9'd51,-10'd349};
ram[56173] = {9'd54,-10'd346};
ram[56174] = {9'd58,-10'd343};
ram[56175] = {9'd61,-10'd340};
ram[56176] = {9'd64,-10'd337};
ram[56177] = {9'd67,-10'd334};
ram[56178] = {9'd70,-10'd330};
ram[56179] = {9'd73,-10'd327};
ram[56180] = {9'd76,-10'd324};
ram[56181] = {9'd80,-10'd321};
ram[56182] = {9'd83,-10'd318};
ram[56183] = {9'd86,-10'd315};
ram[56184] = {9'd89,-10'd312};
ram[56185] = {9'd92,-10'd308};
ram[56186] = {9'd95,-10'd305};
ram[56187] = {9'd98,-10'd302};
ram[56188] = {-9'd99,-10'd299};
ram[56189] = {-9'd96,-10'd296};
ram[56190] = {-9'd92,-10'd293};
ram[56191] = {-9'd89,-10'd290};
ram[56192] = {-9'd89,-10'd290};
ram[56193] = {-9'd86,-10'd286};
ram[56194] = {-9'd83,-10'd283};
ram[56195] = {-9'd80,-10'd280};
ram[56196] = {-9'd77,-10'd277};
ram[56197] = {-9'd74,-10'd274};
ram[56198] = {-9'd70,-10'd271};
ram[56199] = {-9'd67,-10'd268};
ram[56200] = {-9'd64,-10'd264};
ram[56201] = {-9'd61,-10'd261};
ram[56202] = {-9'd58,-10'd258};
ram[56203] = {-9'd55,-10'd255};
ram[56204] = {-9'd52,-10'd252};
ram[56205] = {-9'd48,-10'd249};
ram[56206] = {-9'd45,-10'd246};
ram[56207] = {-9'd42,-10'd242};
ram[56208] = {-9'd39,-10'd239};
ram[56209] = {-9'd36,-10'd236};
ram[56210] = {-9'd33,-10'd233};
ram[56211] = {-9'd30,-10'd230};
ram[56212] = {-9'd26,-10'd227};
ram[56213] = {-9'd23,-10'd224};
ram[56214] = {-9'd20,-10'd220};
ram[56215] = {-9'd17,-10'd217};
ram[56216] = {-9'd14,-10'd214};
ram[56217] = {-9'd11,-10'd211};
ram[56218] = {-9'd8,-10'd208};
ram[56219] = {-9'd4,-10'd205};
ram[56220] = {-9'd1,-10'd202};
ram[56221] = {9'd2,-10'd198};
ram[56222] = {9'd5,-10'd195};
ram[56223] = {9'd8,-10'd192};
ram[56224] = {9'd11,-10'd189};
ram[56225] = {9'd14,-10'd186};
ram[56226] = {9'd18,-10'd183};
ram[56227] = {9'd21,-10'd180};
ram[56228] = {9'd24,-10'd176};
ram[56229] = {9'd27,-10'd173};
ram[56230] = {9'd30,-10'd170};
ram[56231] = {9'd33,-10'd167};
ram[56232] = {9'd36,-10'd164};
ram[56233] = {9'd40,-10'd161};
ram[56234] = {9'd43,-10'd158};
ram[56235] = {9'd46,-10'd154};
ram[56236] = {9'd49,-10'd151};
ram[56237] = {9'd52,-10'd148};
ram[56238] = {9'd55,-10'd145};
ram[56239] = {9'd58,-10'd142};
ram[56240] = {9'd62,-10'd139};
ram[56241] = {9'd65,-10'd136};
ram[56242] = {9'd68,-10'd132};
ram[56243] = {9'd71,-10'd129};
ram[56244] = {9'd74,-10'd126};
ram[56245] = {9'd77,-10'd123};
ram[56246] = {9'd80,-10'd120};
ram[56247] = {9'd84,-10'd117};
ram[56248] = {9'd87,-10'd114};
ram[56249] = {9'd90,-10'd110};
ram[56250] = {9'd93,-10'd107};
ram[56251] = {9'd96,-10'd104};
ram[56252] = {9'd99,-10'd101};
ram[56253] = {-9'd98,-10'd98};
ram[56254] = {-9'd95,-10'd95};
ram[56255] = {-9'd92,-10'd92};
ram[56256] = {-9'd88,-10'd88};
ram[56257] = {-9'd85,-10'd85};
ram[56258] = {-9'd82,-10'd82};
ram[56259] = {-9'd79,-10'd79};
ram[56260] = {-9'd76,-10'd76};
ram[56261] = {-9'd73,-10'd73};
ram[56262] = {-9'd70,-10'd70};
ram[56263] = {-9'd66,-10'd66};
ram[56264] = {-9'd63,-10'd63};
ram[56265] = {-9'd60,-10'd60};
ram[56266] = {-9'd57,-10'd57};
ram[56267] = {-9'd54,-10'd54};
ram[56268] = {-9'd51,-10'd51};
ram[56269] = {-9'd48,-10'd48};
ram[56270] = {-9'd44,-10'd44};
ram[56271] = {-9'd41,-10'd41};
ram[56272] = {-9'd38,-10'd38};
ram[56273] = {-9'd35,-10'd35};
ram[56274] = {-9'd32,-10'd32};
ram[56275] = {-9'd29,-10'd29};
ram[56276] = {-9'd26,-10'd26};
ram[56277] = {-9'd22,-10'd22};
ram[56278] = {-9'd19,-10'd19};
ram[56279] = {-9'd16,-10'd16};
ram[56280] = {-9'd13,-10'd13};
ram[56281] = {-9'd10,-10'd10};
ram[56282] = {-9'd7,-10'd7};
ram[56283] = {-9'd4,-10'd4};
ram[56284] = {-9'd1,-10'd1};
ram[56285] = {9'd3,10'd3};
ram[56286] = {9'd6,10'd6};
ram[56287] = {9'd9,10'd9};
ram[56288] = {9'd12,10'd12};
ram[56289] = {9'd15,10'd15};
ram[56290] = {9'd18,10'd18};
ram[56291] = {9'd21,10'd21};
ram[56292] = {9'd25,10'd25};
ram[56293] = {9'd28,10'd28};
ram[56294] = {9'd31,10'd31};
ram[56295] = {9'd34,10'd34};
ram[56296] = {9'd37,10'd37};
ram[56297] = {9'd40,10'd40};
ram[56298] = {9'd43,10'd43};
ram[56299] = {9'd47,10'd47};
ram[56300] = {9'd50,10'd50};
ram[56301] = {9'd53,10'd53};
ram[56302] = {9'd56,10'd56};
ram[56303] = {9'd59,10'd59};
ram[56304] = {9'd62,10'd62};
ram[56305] = {9'd65,10'd65};
ram[56306] = {9'd69,10'd69};
ram[56307] = {9'd72,10'd72};
ram[56308] = {9'd75,10'd75};
ram[56309] = {9'd78,10'd78};
ram[56310] = {9'd81,10'd81};
ram[56311] = {9'd84,10'd84};
ram[56312] = {9'd87,10'd87};
ram[56313] = {9'd91,10'd91};
ram[56314] = {9'd94,10'd94};
ram[56315] = {9'd97,10'd97};
ram[56316] = {-9'd100,10'd100};
ram[56317] = {-9'd97,10'd103};
ram[56318] = {-9'd94,10'd106};
ram[56319] = {-9'd91,10'd109};
ram[56320] = {-9'd91,10'd109};
ram[56321] = {-9'd88,10'd113};
ram[56322] = {-9'd85,10'd116};
ram[56323] = {-9'd81,10'd119};
ram[56324] = {-9'd78,10'd122};
ram[56325] = {-9'd75,10'd125};
ram[56326] = {-9'd72,10'd128};
ram[56327] = {-9'd69,10'd131};
ram[56328] = {-9'd66,10'd135};
ram[56329] = {-9'd63,10'd138};
ram[56330] = {-9'd59,10'd141};
ram[56331] = {-9'd56,10'd144};
ram[56332] = {-9'd53,10'd147};
ram[56333] = {-9'd50,10'd150};
ram[56334] = {-9'd47,10'd153};
ram[56335] = {-9'd44,10'd157};
ram[56336] = {-9'd41,10'd160};
ram[56337] = {-9'd37,10'd163};
ram[56338] = {-9'd34,10'd166};
ram[56339] = {-9'd31,10'd169};
ram[56340] = {-9'd28,10'd172};
ram[56341] = {-9'd25,10'd175};
ram[56342] = {-9'd22,10'd179};
ram[56343] = {-9'd19,10'd182};
ram[56344] = {-9'd15,10'd185};
ram[56345] = {-9'd12,10'd188};
ram[56346] = {-9'd9,10'd191};
ram[56347] = {-9'd6,10'd194};
ram[56348] = {-9'd3,10'd197};
ram[56349] = {9'd0,10'd201};
ram[56350] = {9'd3,10'd204};
ram[56351] = {9'd7,10'd207};
ram[56352] = {9'd10,10'd210};
ram[56353] = {9'd13,10'd213};
ram[56354] = {9'd16,10'd216};
ram[56355] = {9'd19,10'd219};
ram[56356] = {9'd22,10'd223};
ram[56357] = {9'd25,10'd226};
ram[56358] = {9'd29,10'd229};
ram[56359] = {9'd32,10'd232};
ram[56360] = {9'd35,10'd235};
ram[56361] = {9'd38,10'd238};
ram[56362] = {9'd41,10'd241};
ram[56363] = {9'd44,10'd245};
ram[56364] = {9'd47,10'd248};
ram[56365] = {9'd51,10'd251};
ram[56366] = {9'd54,10'd254};
ram[56367] = {9'd57,10'd257};
ram[56368] = {9'd60,10'd260};
ram[56369] = {9'd63,10'd263};
ram[56370] = {9'd66,10'd267};
ram[56371] = {9'd69,10'd270};
ram[56372] = {9'd73,10'd273};
ram[56373] = {9'd76,10'd276};
ram[56374] = {9'd79,10'd279};
ram[56375] = {9'd82,10'd282};
ram[56376] = {9'd85,10'd285};
ram[56377] = {9'd88,10'd289};
ram[56378] = {9'd91,10'd292};
ram[56379] = {9'd95,10'd295};
ram[56380] = {9'd98,10'd298};
ram[56381] = {-9'd99,10'd301};
ram[56382] = {-9'd96,10'd304};
ram[56383] = {-9'd93,10'd307};
ram[56384] = {-9'd90,10'd311};
ram[56385] = {-9'd87,10'd314};
ram[56386] = {-9'd84,10'd317};
ram[56387] = {-9'd81,10'd320};
ram[56388] = {-9'd77,10'd323};
ram[56389] = {-9'd74,10'd326};
ram[56390] = {-9'd71,10'd329};
ram[56391] = {-9'd68,10'd333};
ram[56392] = {-9'd65,10'd336};
ram[56393] = {-9'd62,10'd339};
ram[56394] = {-9'd59,10'd342};
ram[56395] = {-9'd55,10'd345};
ram[56396] = {-9'd52,10'd348};
ram[56397] = {-9'd49,10'd351};
ram[56398] = {-9'd46,10'd354};
ram[56399] = {-9'd43,10'd358};
ram[56400] = {-9'd40,10'd361};
ram[56401] = {-9'd37,10'd364};
ram[56402] = {-9'd33,10'd367};
ram[56403] = {-9'd30,10'd370};
ram[56404] = {-9'd27,10'd373};
ram[56405] = {-9'd24,10'd376};
ram[56406] = {-9'd21,10'd380};
ram[56407] = {-9'd18,10'd383};
ram[56408] = {-9'd15,10'd386};
ram[56409] = {-9'd11,10'd389};
ram[56410] = {-9'd8,10'd392};
ram[56411] = {-9'd5,10'd395};
ram[56412] = {-9'd2,10'd398};
ram[56413] = {9'd1,-10'd399};
ram[56414] = {9'd4,-10'd396};
ram[56415] = {9'd7,-10'd393};
ram[56416] = {9'd10,-10'd390};
ram[56417] = {9'd14,-10'd387};
ram[56418] = {9'd17,-10'd384};
ram[56419] = {9'd20,-10'd381};
ram[56420] = {9'd23,-10'd377};
ram[56421] = {9'd26,-10'd374};
ram[56422] = {9'd29,-10'd371};
ram[56423] = {9'd32,-10'd368};
ram[56424] = {9'd36,-10'd365};
ram[56425] = {9'd39,-10'd362};
ram[56426] = {9'd42,-10'd359};
ram[56427] = {9'd45,-10'd355};
ram[56428] = {9'd48,-10'd352};
ram[56429] = {9'd51,-10'd349};
ram[56430] = {9'd54,-10'd346};
ram[56431] = {9'd58,-10'd343};
ram[56432] = {9'd61,-10'd340};
ram[56433] = {9'd64,-10'd337};
ram[56434] = {9'd67,-10'd334};
ram[56435] = {9'd70,-10'd330};
ram[56436] = {9'd73,-10'd327};
ram[56437] = {9'd76,-10'd324};
ram[56438] = {9'd80,-10'd321};
ram[56439] = {9'd83,-10'd318};
ram[56440] = {9'd86,-10'd315};
ram[56441] = {9'd89,-10'd312};
ram[56442] = {9'd92,-10'd308};
ram[56443] = {9'd95,-10'd305};
ram[56444] = {9'd98,-10'd302};
ram[56445] = {-9'd99,-10'd299};
ram[56446] = {-9'd96,-10'd296};
ram[56447] = {-9'd92,-10'd293};
ram[56448] = {-9'd92,-10'd293};
ram[56449] = {-9'd89,-10'd290};
ram[56450] = {-9'd86,-10'd286};
ram[56451] = {-9'd83,-10'd283};
ram[56452] = {-9'd80,-10'd280};
ram[56453] = {-9'd77,-10'd277};
ram[56454] = {-9'd74,-10'd274};
ram[56455] = {-9'd70,-10'd271};
ram[56456] = {-9'd67,-10'd268};
ram[56457] = {-9'd64,-10'd264};
ram[56458] = {-9'd61,-10'd261};
ram[56459] = {-9'd58,-10'd258};
ram[56460] = {-9'd55,-10'd255};
ram[56461] = {-9'd52,-10'd252};
ram[56462] = {-9'd48,-10'd249};
ram[56463] = {-9'd45,-10'd246};
ram[56464] = {-9'd42,-10'd242};
ram[56465] = {-9'd39,-10'd239};
ram[56466] = {-9'd36,-10'd236};
ram[56467] = {-9'd33,-10'd233};
ram[56468] = {-9'd30,-10'd230};
ram[56469] = {-9'd26,-10'd227};
ram[56470] = {-9'd23,-10'd224};
ram[56471] = {-9'd20,-10'd220};
ram[56472] = {-9'd17,-10'd217};
ram[56473] = {-9'd14,-10'd214};
ram[56474] = {-9'd11,-10'd211};
ram[56475] = {-9'd8,-10'd208};
ram[56476] = {-9'd4,-10'd205};
ram[56477] = {-9'd1,-10'd202};
ram[56478] = {9'd2,-10'd198};
ram[56479] = {9'd5,-10'd195};
ram[56480] = {9'd8,-10'd192};
ram[56481] = {9'd11,-10'd189};
ram[56482] = {9'd14,-10'd186};
ram[56483] = {9'd18,-10'd183};
ram[56484] = {9'd21,-10'd180};
ram[56485] = {9'd24,-10'd176};
ram[56486] = {9'd27,-10'd173};
ram[56487] = {9'd30,-10'd170};
ram[56488] = {9'd33,-10'd167};
ram[56489] = {9'd36,-10'd164};
ram[56490] = {9'd40,-10'd161};
ram[56491] = {9'd43,-10'd158};
ram[56492] = {9'd46,-10'd154};
ram[56493] = {9'd49,-10'd151};
ram[56494] = {9'd52,-10'd148};
ram[56495] = {9'd55,-10'd145};
ram[56496] = {9'd58,-10'd142};
ram[56497] = {9'd62,-10'd139};
ram[56498] = {9'd65,-10'd136};
ram[56499] = {9'd68,-10'd132};
ram[56500] = {9'd71,-10'd129};
ram[56501] = {9'd74,-10'd126};
ram[56502] = {9'd77,-10'd123};
ram[56503] = {9'd80,-10'd120};
ram[56504] = {9'd84,-10'd117};
ram[56505] = {9'd87,-10'd114};
ram[56506] = {9'd90,-10'd110};
ram[56507] = {9'd93,-10'd107};
ram[56508] = {9'd96,-10'd104};
ram[56509] = {9'd99,-10'd101};
ram[56510] = {-9'd98,-10'd98};
ram[56511] = {-9'd95,-10'd95};
ram[56512] = {-9'd92,-10'd92};
ram[56513] = {-9'd88,-10'd88};
ram[56514] = {-9'd85,-10'd85};
ram[56515] = {-9'd82,-10'd82};
ram[56516] = {-9'd79,-10'd79};
ram[56517] = {-9'd76,-10'd76};
ram[56518] = {-9'd73,-10'd73};
ram[56519] = {-9'd70,-10'd70};
ram[56520] = {-9'd66,-10'd66};
ram[56521] = {-9'd63,-10'd63};
ram[56522] = {-9'd60,-10'd60};
ram[56523] = {-9'd57,-10'd57};
ram[56524] = {-9'd54,-10'd54};
ram[56525] = {-9'd51,-10'd51};
ram[56526] = {-9'd48,-10'd48};
ram[56527] = {-9'd44,-10'd44};
ram[56528] = {-9'd41,-10'd41};
ram[56529] = {-9'd38,-10'd38};
ram[56530] = {-9'd35,-10'd35};
ram[56531] = {-9'd32,-10'd32};
ram[56532] = {-9'd29,-10'd29};
ram[56533] = {-9'd26,-10'd26};
ram[56534] = {-9'd22,-10'd22};
ram[56535] = {-9'd19,-10'd19};
ram[56536] = {-9'd16,-10'd16};
ram[56537] = {-9'd13,-10'd13};
ram[56538] = {-9'd10,-10'd10};
ram[56539] = {-9'd7,-10'd7};
ram[56540] = {-9'd4,-10'd4};
ram[56541] = {-9'd1,-10'd1};
ram[56542] = {9'd3,10'd3};
ram[56543] = {9'd6,10'd6};
ram[56544] = {9'd9,10'd9};
ram[56545] = {9'd12,10'd12};
ram[56546] = {9'd15,10'd15};
ram[56547] = {9'd18,10'd18};
ram[56548] = {9'd21,10'd21};
ram[56549] = {9'd25,10'd25};
ram[56550] = {9'd28,10'd28};
ram[56551] = {9'd31,10'd31};
ram[56552] = {9'd34,10'd34};
ram[56553] = {9'd37,10'd37};
ram[56554] = {9'd40,10'd40};
ram[56555] = {9'd43,10'd43};
ram[56556] = {9'd47,10'd47};
ram[56557] = {9'd50,10'd50};
ram[56558] = {9'd53,10'd53};
ram[56559] = {9'd56,10'd56};
ram[56560] = {9'd59,10'd59};
ram[56561] = {9'd62,10'd62};
ram[56562] = {9'd65,10'd65};
ram[56563] = {9'd69,10'd69};
ram[56564] = {9'd72,10'd72};
ram[56565] = {9'd75,10'd75};
ram[56566] = {9'd78,10'd78};
ram[56567] = {9'd81,10'd81};
ram[56568] = {9'd84,10'd84};
ram[56569] = {9'd87,10'd87};
ram[56570] = {9'd91,10'd91};
ram[56571] = {9'd94,10'd94};
ram[56572] = {9'd97,10'd97};
ram[56573] = {-9'd100,10'd100};
ram[56574] = {-9'd97,10'd103};
ram[56575] = {-9'd94,10'd106};
ram[56576] = {-9'd94,10'd106};
ram[56577] = {-9'd91,10'd109};
ram[56578] = {-9'd88,10'd113};
ram[56579] = {-9'd85,10'd116};
ram[56580] = {-9'd81,10'd119};
ram[56581] = {-9'd78,10'd122};
ram[56582] = {-9'd75,10'd125};
ram[56583] = {-9'd72,10'd128};
ram[56584] = {-9'd69,10'd131};
ram[56585] = {-9'd66,10'd135};
ram[56586] = {-9'd63,10'd138};
ram[56587] = {-9'd59,10'd141};
ram[56588] = {-9'd56,10'd144};
ram[56589] = {-9'd53,10'd147};
ram[56590] = {-9'd50,10'd150};
ram[56591] = {-9'd47,10'd153};
ram[56592] = {-9'd44,10'd157};
ram[56593] = {-9'd41,10'd160};
ram[56594] = {-9'd37,10'd163};
ram[56595] = {-9'd34,10'd166};
ram[56596] = {-9'd31,10'd169};
ram[56597] = {-9'd28,10'd172};
ram[56598] = {-9'd25,10'd175};
ram[56599] = {-9'd22,10'd179};
ram[56600] = {-9'd19,10'd182};
ram[56601] = {-9'd15,10'd185};
ram[56602] = {-9'd12,10'd188};
ram[56603] = {-9'd9,10'd191};
ram[56604] = {-9'd6,10'd194};
ram[56605] = {-9'd3,10'd197};
ram[56606] = {9'd0,10'd201};
ram[56607] = {9'd3,10'd204};
ram[56608] = {9'd7,10'd207};
ram[56609] = {9'd10,10'd210};
ram[56610] = {9'd13,10'd213};
ram[56611] = {9'd16,10'd216};
ram[56612] = {9'd19,10'd219};
ram[56613] = {9'd22,10'd223};
ram[56614] = {9'd25,10'd226};
ram[56615] = {9'd29,10'd229};
ram[56616] = {9'd32,10'd232};
ram[56617] = {9'd35,10'd235};
ram[56618] = {9'd38,10'd238};
ram[56619] = {9'd41,10'd241};
ram[56620] = {9'd44,10'd245};
ram[56621] = {9'd47,10'd248};
ram[56622] = {9'd51,10'd251};
ram[56623] = {9'd54,10'd254};
ram[56624] = {9'd57,10'd257};
ram[56625] = {9'd60,10'd260};
ram[56626] = {9'd63,10'd263};
ram[56627] = {9'd66,10'd267};
ram[56628] = {9'd69,10'd270};
ram[56629] = {9'd73,10'd273};
ram[56630] = {9'd76,10'd276};
ram[56631] = {9'd79,10'd279};
ram[56632] = {9'd82,10'd282};
ram[56633] = {9'd85,10'd285};
ram[56634] = {9'd88,10'd289};
ram[56635] = {9'd91,10'd292};
ram[56636] = {9'd95,10'd295};
ram[56637] = {9'd98,10'd298};
ram[56638] = {-9'd99,10'd301};
ram[56639] = {-9'd96,10'd304};
ram[56640] = {-9'd93,10'd307};
ram[56641] = {-9'd90,10'd311};
ram[56642] = {-9'd87,10'd314};
ram[56643] = {-9'd84,10'd317};
ram[56644] = {-9'd81,10'd320};
ram[56645] = {-9'd77,10'd323};
ram[56646] = {-9'd74,10'd326};
ram[56647] = {-9'd71,10'd329};
ram[56648] = {-9'd68,10'd333};
ram[56649] = {-9'd65,10'd336};
ram[56650] = {-9'd62,10'd339};
ram[56651] = {-9'd59,10'd342};
ram[56652] = {-9'd55,10'd345};
ram[56653] = {-9'd52,10'd348};
ram[56654] = {-9'd49,10'd351};
ram[56655] = {-9'd46,10'd354};
ram[56656] = {-9'd43,10'd358};
ram[56657] = {-9'd40,10'd361};
ram[56658] = {-9'd37,10'd364};
ram[56659] = {-9'd33,10'd367};
ram[56660] = {-9'd30,10'd370};
ram[56661] = {-9'd27,10'd373};
ram[56662] = {-9'd24,10'd376};
ram[56663] = {-9'd21,10'd380};
ram[56664] = {-9'd18,10'd383};
ram[56665] = {-9'd15,10'd386};
ram[56666] = {-9'd11,10'd389};
ram[56667] = {-9'd8,10'd392};
ram[56668] = {-9'd5,10'd395};
ram[56669] = {-9'd2,10'd398};
ram[56670] = {9'd1,-10'd399};
ram[56671] = {9'd4,-10'd396};
ram[56672] = {9'd7,-10'd393};
ram[56673] = {9'd10,-10'd390};
ram[56674] = {9'd14,-10'd387};
ram[56675] = {9'd17,-10'd384};
ram[56676] = {9'd20,-10'd381};
ram[56677] = {9'd23,-10'd377};
ram[56678] = {9'd26,-10'd374};
ram[56679] = {9'd29,-10'd371};
ram[56680] = {9'd32,-10'd368};
ram[56681] = {9'd36,-10'd365};
ram[56682] = {9'd39,-10'd362};
ram[56683] = {9'd42,-10'd359};
ram[56684] = {9'd45,-10'd355};
ram[56685] = {9'd48,-10'd352};
ram[56686] = {9'd51,-10'd349};
ram[56687] = {9'd54,-10'd346};
ram[56688] = {9'd58,-10'd343};
ram[56689] = {9'd61,-10'd340};
ram[56690] = {9'd64,-10'd337};
ram[56691] = {9'd67,-10'd334};
ram[56692] = {9'd70,-10'd330};
ram[56693] = {9'd73,-10'd327};
ram[56694] = {9'd76,-10'd324};
ram[56695] = {9'd80,-10'd321};
ram[56696] = {9'd83,-10'd318};
ram[56697] = {9'd86,-10'd315};
ram[56698] = {9'd89,-10'd312};
ram[56699] = {9'd92,-10'd308};
ram[56700] = {9'd95,-10'd305};
ram[56701] = {9'd98,-10'd302};
ram[56702] = {-9'd99,-10'd299};
ram[56703] = {-9'd96,-10'd296};
ram[56704] = {-9'd96,-10'd296};
ram[56705] = {-9'd92,-10'd293};
ram[56706] = {-9'd89,-10'd290};
ram[56707] = {-9'd86,-10'd286};
ram[56708] = {-9'd83,-10'd283};
ram[56709] = {-9'd80,-10'd280};
ram[56710] = {-9'd77,-10'd277};
ram[56711] = {-9'd74,-10'd274};
ram[56712] = {-9'd70,-10'd271};
ram[56713] = {-9'd67,-10'd268};
ram[56714] = {-9'd64,-10'd264};
ram[56715] = {-9'd61,-10'd261};
ram[56716] = {-9'd58,-10'd258};
ram[56717] = {-9'd55,-10'd255};
ram[56718] = {-9'd52,-10'd252};
ram[56719] = {-9'd48,-10'd249};
ram[56720] = {-9'd45,-10'd246};
ram[56721] = {-9'd42,-10'd242};
ram[56722] = {-9'd39,-10'd239};
ram[56723] = {-9'd36,-10'd236};
ram[56724] = {-9'd33,-10'd233};
ram[56725] = {-9'd30,-10'd230};
ram[56726] = {-9'd26,-10'd227};
ram[56727] = {-9'd23,-10'd224};
ram[56728] = {-9'd20,-10'd220};
ram[56729] = {-9'd17,-10'd217};
ram[56730] = {-9'd14,-10'd214};
ram[56731] = {-9'd11,-10'd211};
ram[56732] = {-9'd8,-10'd208};
ram[56733] = {-9'd4,-10'd205};
ram[56734] = {-9'd1,-10'd202};
ram[56735] = {9'd2,-10'd198};
ram[56736] = {9'd5,-10'd195};
ram[56737] = {9'd8,-10'd192};
ram[56738] = {9'd11,-10'd189};
ram[56739] = {9'd14,-10'd186};
ram[56740] = {9'd18,-10'd183};
ram[56741] = {9'd21,-10'd180};
ram[56742] = {9'd24,-10'd176};
ram[56743] = {9'd27,-10'd173};
ram[56744] = {9'd30,-10'd170};
ram[56745] = {9'd33,-10'd167};
ram[56746] = {9'd36,-10'd164};
ram[56747] = {9'd40,-10'd161};
ram[56748] = {9'd43,-10'd158};
ram[56749] = {9'd46,-10'd154};
ram[56750] = {9'd49,-10'd151};
ram[56751] = {9'd52,-10'd148};
ram[56752] = {9'd55,-10'd145};
ram[56753] = {9'd58,-10'd142};
ram[56754] = {9'd62,-10'd139};
ram[56755] = {9'd65,-10'd136};
ram[56756] = {9'd68,-10'd132};
ram[56757] = {9'd71,-10'd129};
ram[56758] = {9'd74,-10'd126};
ram[56759] = {9'd77,-10'd123};
ram[56760] = {9'd80,-10'd120};
ram[56761] = {9'd84,-10'd117};
ram[56762] = {9'd87,-10'd114};
ram[56763] = {9'd90,-10'd110};
ram[56764] = {9'd93,-10'd107};
ram[56765] = {9'd96,-10'd104};
ram[56766] = {9'd99,-10'd101};
ram[56767] = {-9'd98,-10'd98};
ram[56768] = {-9'd95,-10'd95};
ram[56769] = {-9'd92,-10'd92};
ram[56770] = {-9'd88,-10'd88};
ram[56771] = {-9'd85,-10'd85};
ram[56772] = {-9'd82,-10'd82};
ram[56773] = {-9'd79,-10'd79};
ram[56774] = {-9'd76,-10'd76};
ram[56775] = {-9'd73,-10'd73};
ram[56776] = {-9'd70,-10'd70};
ram[56777] = {-9'd66,-10'd66};
ram[56778] = {-9'd63,-10'd63};
ram[56779] = {-9'd60,-10'd60};
ram[56780] = {-9'd57,-10'd57};
ram[56781] = {-9'd54,-10'd54};
ram[56782] = {-9'd51,-10'd51};
ram[56783] = {-9'd48,-10'd48};
ram[56784] = {-9'd44,-10'd44};
ram[56785] = {-9'd41,-10'd41};
ram[56786] = {-9'd38,-10'd38};
ram[56787] = {-9'd35,-10'd35};
ram[56788] = {-9'd32,-10'd32};
ram[56789] = {-9'd29,-10'd29};
ram[56790] = {-9'd26,-10'd26};
ram[56791] = {-9'd22,-10'd22};
ram[56792] = {-9'd19,-10'd19};
ram[56793] = {-9'd16,-10'd16};
ram[56794] = {-9'd13,-10'd13};
ram[56795] = {-9'd10,-10'd10};
ram[56796] = {-9'd7,-10'd7};
ram[56797] = {-9'd4,-10'd4};
ram[56798] = {-9'd1,-10'd1};
ram[56799] = {9'd3,10'd3};
ram[56800] = {9'd6,10'd6};
ram[56801] = {9'd9,10'd9};
ram[56802] = {9'd12,10'd12};
ram[56803] = {9'd15,10'd15};
ram[56804] = {9'd18,10'd18};
ram[56805] = {9'd21,10'd21};
ram[56806] = {9'd25,10'd25};
ram[56807] = {9'd28,10'd28};
ram[56808] = {9'd31,10'd31};
ram[56809] = {9'd34,10'd34};
ram[56810] = {9'd37,10'd37};
ram[56811] = {9'd40,10'd40};
ram[56812] = {9'd43,10'd43};
ram[56813] = {9'd47,10'd47};
ram[56814] = {9'd50,10'd50};
ram[56815] = {9'd53,10'd53};
ram[56816] = {9'd56,10'd56};
ram[56817] = {9'd59,10'd59};
ram[56818] = {9'd62,10'd62};
ram[56819] = {9'd65,10'd65};
ram[56820] = {9'd69,10'd69};
ram[56821] = {9'd72,10'd72};
ram[56822] = {9'd75,10'd75};
ram[56823] = {9'd78,10'd78};
ram[56824] = {9'd81,10'd81};
ram[56825] = {9'd84,10'd84};
ram[56826] = {9'd87,10'd87};
ram[56827] = {9'd91,10'd91};
ram[56828] = {9'd94,10'd94};
ram[56829] = {9'd97,10'd97};
ram[56830] = {-9'd100,10'd100};
ram[56831] = {-9'd97,10'd103};
ram[56832] = {-9'd97,10'd103};
ram[56833] = {-9'd94,10'd106};
ram[56834] = {-9'd91,10'd109};
ram[56835] = {-9'd88,10'd113};
ram[56836] = {-9'd85,10'd116};
ram[56837] = {-9'd81,10'd119};
ram[56838] = {-9'd78,10'd122};
ram[56839] = {-9'd75,10'd125};
ram[56840] = {-9'd72,10'd128};
ram[56841] = {-9'd69,10'd131};
ram[56842] = {-9'd66,10'd135};
ram[56843] = {-9'd63,10'd138};
ram[56844] = {-9'd59,10'd141};
ram[56845] = {-9'd56,10'd144};
ram[56846] = {-9'd53,10'd147};
ram[56847] = {-9'd50,10'd150};
ram[56848] = {-9'd47,10'd153};
ram[56849] = {-9'd44,10'd157};
ram[56850] = {-9'd41,10'd160};
ram[56851] = {-9'd37,10'd163};
ram[56852] = {-9'd34,10'd166};
ram[56853] = {-9'd31,10'd169};
ram[56854] = {-9'd28,10'd172};
ram[56855] = {-9'd25,10'd175};
ram[56856] = {-9'd22,10'd179};
ram[56857] = {-9'd19,10'd182};
ram[56858] = {-9'd15,10'd185};
ram[56859] = {-9'd12,10'd188};
ram[56860] = {-9'd9,10'd191};
ram[56861] = {-9'd6,10'd194};
ram[56862] = {-9'd3,10'd197};
ram[56863] = {9'd0,10'd201};
ram[56864] = {9'd3,10'd204};
ram[56865] = {9'd7,10'd207};
ram[56866] = {9'd10,10'd210};
ram[56867] = {9'd13,10'd213};
ram[56868] = {9'd16,10'd216};
ram[56869] = {9'd19,10'd219};
ram[56870] = {9'd22,10'd223};
ram[56871] = {9'd25,10'd226};
ram[56872] = {9'd29,10'd229};
ram[56873] = {9'd32,10'd232};
ram[56874] = {9'd35,10'd235};
ram[56875] = {9'd38,10'd238};
ram[56876] = {9'd41,10'd241};
ram[56877] = {9'd44,10'd245};
ram[56878] = {9'd47,10'd248};
ram[56879] = {9'd51,10'd251};
ram[56880] = {9'd54,10'd254};
ram[56881] = {9'd57,10'd257};
ram[56882] = {9'd60,10'd260};
ram[56883] = {9'd63,10'd263};
ram[56884] = {9'd66,10'd267};
ram[56885] = {9'd69,10'd270};
ram[56886] = {9'd73,10'd273};
ram[56887] = {9'd76,10'd276};
ram[56888] = {9'd79,10'd279};
ram[56889] = {9'd82,10'd282};
ram[56890] = {9'd85,10'd285};
ram[56891] = {9'd88,10'd289};
ram[56892] = {9'd91,10'd292};
ram[56893] = {9'd95,10'd295};
ram[56894] = {9'd98,10'd298};
ram[56895] = {-9'd99,10'd301};
ram[56896] = {-9'd96,10'd304};
ram[56897] = {-9'd93,10'd307};
ram[56898] = {-9'd90,10'd311};
ram[56899] = {-9'd87,10'd314};
ram[56900] = {-9'd84,10'd317};
ram[56901] = {-9'd81,10'd320};
ram[56902] = {-9'd77,10'd323};
ram[56903] = {-9'd74,10'd326};
ram[56904] = {-9'd71,10'd329};
ram[56905] = {-9'd68,10'd333};
ram[56906] = {-9'd65,10'd336};
ram[56907] = {-9'd62,10'd339};
ram[56908] = {-9'd59,10'd342};
ram[56909] = {-9'd55,10'd345};
ram[56910] = {-9'd52,10'd348};
ram[56911] = {-9'd49,10'd351};
ram[56912] = {-9'd46,10'd354};
ram[56913] = {-9'd43,10'd358};
ram[56914] = {-9'd40,10'd361};
ram[56915] = {-9'd37,10'd364};
ram[56916] = {-9'd33,10'd367};
ram[56917] = {-9'd30,10'd370};
ram[56918] = {-9'd27,10'd373};
ram[56919] = {-9'd24,10'd376};
ram[56920] = {-9'd21,10'd380};
ram[56921] = {-9'd18,10'd383};
ram[56922] = {-9'd15,10'd386};
ram[56923] = {-9'd11,10'd389};
ram[56924] = {-9'd8,10'd392};
ram[56925] = {-9'd5,10'd395};
ram[56926] = {-9'd2,10'd398};
ram[56927] = {9'd1,-10'd399};
ram[56928] = {9'd4,-10'd396};
ram[56929] = {9'd7,-10'd393};
ram[56930] = {9'd10,-10'd390};
ram[56931] = {9'd14,-10'd387};
ram[56932] = {9'd17,-10'd384};
ram[56933] = {9'd20,-10'd381};
ram[56934] = {9'd23,-10'd377};
ram[56935] = {9'd26,-10'd374};
ram[56936] = {9'd29,-10'd371};
ram[56937] = {9'd32,-10'd368};
ram[56938] = {9'd36,-10'd365};
ram[56939] = {9'd39,-10'd362};
ram[56940] = {9'd42,-10'd359};
ram[56941] = {9'd45,-10'd355};
ram[56942] = {9'd48,-10'd352};
ram[56943] = {9'd51,-10'd349};
ram[56944] = {9'd54,-10'd346};
ram[56945] = {9'd58,-10'd343};
ram[56946] = {9'd61,-10'd340};
ram[56947] = {9'd64,-10'd337};
ram[56948] = {9'd67,-10'd334};
ram[56949] = {9'd70,-10'd330};
ram[56950] = {9'd73,-10'd327};
ram[56951] = {9'd76,-10'd324};
ram[56952] = {9'd80,-10'd321};
ram[56953] = {9'd83,-10'd318};
ram[56954] = {9'd86,-10'd315};
ram[56955] = {9'd89,-10'd312};
ram[56956] = {9'd92,-10'd308};
ram[56957] = {9'd95,-10'd305};
ram[56958] = {9'd98,-10'd302};
ram[56959] = {-9'd99,-10'd299};
ram[56960] = {-9'd99,-10'd299};
ram[56961] = {-9'd96,-10'd296};
ram[56962] = {-9'd92,-10'd293};
ram[56963] = {-9'd89,-10'd290};
ram[56964] = {-9'd86,-10'd286};
ram[56965] = {-9'd83,-10'd283};
ram[56966] = {-9'd80,-10'd280};
ram[56967] = {-9'd77,-10'd277};
ram[56968] = {-9'd74,-10'd274};
ram[56969] = {-9'd70,-10'd271};
ram[56970] = {-9'd67,-10'd268};
ram[56971] = {-9'd64,-10'd264};
ram[56972] = {-9'd61,-10'd261};
ram[56973] = {-9'd58,-10'd258};
ram[56974] = {-9'd55,-10'd255};
ram[56975] = {-9'd52,-10'd252};
ram[56976] = {-9'd48,-10'd249};
ram[56977] = {-9'd45,-10'd246};
ram[56978] = {-9'd42,-10'd242};
ram[56979] = {-9'd39,-10'd239};
ram[56980] = {-9'd36,-10'd236};
ram[56981] = {-9'd33,-10'd233};
ram[56982] = {-9'd30,-10'd230};
ram[56983] = {-9'd26,-10'd227};
ram[56984] = {-9'd23,-10'd224};
ram[56985] = {-9'd20,-10'd220};
ram[56986] = {-9'd17,-10'd217};
ram[56987] = {-9'd14,-10'd214};
ram[56988] = {-9'd11,-10'd211};
ram[56989] = {-9'd8,-10'd208};
ram[56990] = {-9'd4,-10'd205};
ram[56991] = {-9'd1,-10'd202};
ram[56992] = {9'd2,-10'd198};
ram[56993] = {9'd5,-10'd195};
ram[56994] = {9'd8,-10'd192};
ram[56995] = {9'd11,-10'd189};
ram[56996] = {9'd14,-10'd186};
ram[56997] = {9'd18,-10'd183};
ram[56998] = {9'd21,-10'd180};
ram[56999] = {9'd24,-10'd176};
ram[57000] = {9'd27,-10'd173};
ram[57001] = {9'd30,-10'd170};
ram[57002] = {9'd33,-10'd167};
ram[57003] = {9'd36,-10'd164};
ram[57004] = {9'd40,-10'd161};
ram[57005] = {9'd43,-10'd158};
ram[57006] = {9'd46,-10'd154};
ram[57007] = {9'd49,-10'd151};
ram[57008] = {9'd52,-10'd148};
ram[57009] = {9'd55,-10'd145};
ram[57010] = {9'd58,-10'd142};
ram[57011] = {9'd62,-10'd139};
ram[57012] = {9'd65,-10'd136};
ram[57013] = {9'd68,-10'd132};
ram[57014] = {9'd71,-10'd129};
ram[57015] = {9'd74,-10'd126};
ram[57016] = {9'd77,-10'd123};
ram[57017] = {9'd80,-10'd120};
ram[57018] = {9'd84,-10'd117};
ram[57019] = {9'd87,-10'd114};
ram[57020] = {9'd90,-10'd110};
ram[57021] = {9'd93,-10'd107};
ram[57022] = {9'd96,-10'd104};
ram[57023] = {9'd99,-10'd101};
ram[57024] = {-9'd98,-10'd98};
ram[57025] = {-9'd95,-10'd95};
ram[57026] = {-9'd92,-10'd92};
ram[57027] = {-9'd88,-10'd88};
ram[57028] = {-9'd85,-10'd85};
ram[57029] = {-9'd82,-10'd82};
ram[57030] = {-9'd79,-10'd79};
ram[57031] = {-9'd76,-10'd76};
ram[57032] = {-9'd73,-10'd73};
ram[57033] = {-9'd70,-10'd70};
ram[57034] = {-9'd66,-10'd66};
ram[57035] = {-9'd63,-10'd63};
ram[57036] = {-9'd60,-10'd60};
ram[57037] = {-9'd57,-10'd57};
ram[57038] = {-9'd54,-10'd54};
ram[57039] = {-9'd51,-10'd51};
ram[57040] = {-9'd48,-10'd48};
ram[57041] = {-9'd44,-10'd44};
ram[57042] = {-9'd41,-10'd41};
ram[57043] = {-9'd38,-10'd38};
ram[57044] = {-9'd35,-10'd35};
ram[57045] = {-9'd32,-10'd32};
ram[57046] = {-9'd29,-10'd29};
ram[57047] = {-9'd26,-10'd26};
ram[57048] = {-9'd22,-10'd22};
ram[57049] = {-9'd19,-10'd19};
ram[57050] = {-9'd16,-10'd16};
ram[57051] = {-9'd13,-10'd13};
ram[57052] = {-9'd10,-10'd10};
ram[57053] = {-9'd7,-10'd7};
ram[57054] = {-9'd4,-10'd4};
ram[57055] = {-9'd1,-10'd1};
ram[57056] = {9'd3,10'd3};
ram[57057] = {9'd6,10'd6};
ram[57058] = {9'd9,10'd9};
ram[57059] = {9'd12,10'd12};
ram[57060] = {9'd15,10'd15};
ram[57061] = {9'd18,10'd18};
ram[57062] = {9'd21,10'd21};
ram[57063] = {9'd25,10'd25};
ram[57064] = {9'd28,10'd28};
ram[57065] = {9'd31,10'd31};
ram[57066] = {9'd34,10'd34};
ram[57067] = {9'd37,10'd37};
ram[57068] = {9'd40,10'd40};
ram[57069] = {9'd43,10'd43};
ram[57070] = {9'd47,10'd47};
ram[57071] = {9'd50,10'd50};
ram[57072] = {9'd53,10'd53};
ram[57073] = {9'd56,10'd56};
ram[57074] = {9'd59,10'd59};
ram[57075] = {9'd62,10'd62};
ram[57076] = {9'd65,10'd65};
ram[57077] = {9'd69,10'd69};
ram[57078] = {9'd72,10'd72};
ram[57079] = {9'd75,10'd75};
ram[57080] = {9'd78,10'd78};
ram[57081] = {9'd81,10'd81};
ram[57082] = {9'd84,10'd84};
ram[57083] = {9'd87,10'd87};
ram[57084] = {9'd91,10'd91};
ram[57085] = {9'd94,10'd94};
ram[57086] = {9'd97,10'd97};
ram[57087] = {-9'd100,10'd100};
ram[57088] = {-9'd100,10'd100};
ram[57089] = {-9'd97,10'd103};
ram[57090] = {-9'd94,10'd106};
ram[57091] = {-9'd91,10'd109};
ram[57092] = {-9'd88,10'd113};
ram[57093] = {-9'd85,10'd116};
ram[57094] = {-9'd81,10'd119};
ram[57095] = {-9'd78,10'd122};
ram[57096] = {-9'd75,10'd125};
ram[57097] = {-9'd72,10'd128};
ram[57098] = {-9'd69,10'd131};
ram[57099] = {-9'd66,10'd135};
ram[57100] = {-9'd63,10'd138};
ram[57101] = {-9'd59,10'd141};
ram[57102] = {-9'd56,10'd144};
ram[57103] = {-9'd53,10'd147};
ram[57104] = {-9'd50,10'd150};
ram[57105] = {-9'd47,10'd153};
ram[57106] = {-9'd44,10'd157};
ram[57107] = {-9'd41,10'd160};
ram[57108] = {-9'd37,10'd163};
ram[57109] = {-9'd34,10'd166};
ram[57110] = {-9'd31,10'd169};
ram[57111] = {-9'd28,10'd172};
ram[57112] = {-9'd25,10'd175};
ram[57113] = {-9'd22,10'd179};
ram[57114] = {-9'd19,10'd182};
ram[57115] = {-9'd15,10'd185};
ram[57116] = {-9'd12,10'd188};
ram[57117] = {-9'd9,10'd191};
ram[57118] = {-9'd6,10'd194};
ram[57119] = {-9'd3,10'd197};
ram[57120] = {9'd0,10'd201};
ram[57121] = {9'd3,10'd204};
ram[57122] = {9'd7,10'd207};
ram[57123] = {9'd10,10'd210};
ram[57124] = {9'd13,10'd213};
ram[57125] = {9'd16,10'd216};
ram[57126] = {9'd19,10'd219};
ram[57127] = {9'd22,10'd223};
ram[57128] = {9'd25,10'd226};
ram[57129] = {9'd29,10'd229};
ram[57130] = {9'd32,10'd232};
ram[57131] = {9'd35,10'd235};
ram[57132] = {9'd38,10'd238};
ram[57133] = {9'd41,10'd241};
ram[57134] = {9'd44,10'd245};
ram[57135] = {9'd47,10'd248};
ram[57136] = {9'd51,10'd251};
ram[57137] = {9'd54,10'd254};
ram[57138] = {9'd57,10'd257};
ram[57139] = {9'd60,10'd260};
ram[57140] = {9'd63,10'd263};
ram[57141] = {9'd66,10'd267};
ram[57142] = {9'd69,10'd270};
ram[57143] = {9'd73,10'd273};
ram[57144] = {9'd76,10'd276};
ram[57145] = {9'd79,10'd279};
ram[57146] = {9'd82,10'd282};
ram[57147] = {9'd85,10'd285};
ram[57148] = {9'd88,10'd289};
ram[57149] = {9'd91,10'd292};
ram[57150] = {9'd95,10'd295};
ram[57151] = {9'd98,10'd298};
ram[57152] = {-9'd99,10'd301};
ram[57153] = {-9'd96,10'd304};
ram[57154] = {-9'd93,10'd307};
ram[57155] = {-9'd90,10'd311};
ram[57156] = {-9'd87,10'd314};
ram[57157] = {-9'd84,10'd317};
ram[57158] = {-9'd81,10'd320};
ram[57159] = {-9'd77,10'd323};
ram[57160] = {-9'd74,10'd326};
ram[57161] = {-9'd71,10'd329};
ram[57162] = {-9'd68,10'd333};
ram[57163] = {-9'd65,10'd336};
ram[57164] = {-9'd62,10'd339};
ram[57165] = {-9'd59,10'd342};
ram[57166] = {-9'd55,10'd345};
ram[57167] = {-9'd52,10'd348};
ram[57168] = {-9'd49,10'd351};
ram[57169] = {-9'd46,10'd354};
ram[57170] = {-9'd43,10'd358};
ram[57171] = {-9'd40,10'd361};
ram[57172] = {-9'd37,10'd364};
ram[57173] = {-9'd33,10'd367};
ram[57174] = {-9'd30,10'd370};
ram[57175] = {-9'd27,10'd373};
ram[57176] = {-9'd24,10'd376};
ram[57177] = {-9'd21,10'd380};
ram[57178] = {-9'd18,10'd383};
ram[57179] = {-9'd15,10'd386};
ram[57180] = {-9'd11,10'd389};
ram[57181] = {-9'd8,10'd392};
ram[57182] = {-9'd5,10'd395};
ram[57183] = {-9'd2,10'd398};
ram[57184] = {9'd1,-10'd399};
ram[57185] = {9'd4,-10'd396};
ram[57186] = {9'd7,-10'd393};
ram[57187] = {9'd10,-10'd390};
ram[57188] = {9'd14,-10'd387};
ram[57189] = {9'd17,-10'd384};
ram[57190] = {9'd20,-10'd381};
ram[57191] = {9'd23,-10'd377};
ram[57192] = {9'd26,-10'd374};
ram[57193] = {9'd29,-10'd371};
ram[57194] = {9'd32,-10'd368};
ram[57195] = {9'd36,-10'd365};
ram[57196] = {9'd39,-10'd362};
ram[57197] = {9'd42,-10'd359};
ram[57198] = {9'd45,-10'd355};
ram[57199] = {9'd48,-10'd352};
ram[57200] = {9'd51,-10'd349};
ram[57201] = {9'd54,-10'd346};
ram[57202] = {9'd58,-10'd343};
ram[57203] = {9'd61,-10'd340};
ram[57204] = {9'd64,-10'd337};
ram[57205] = {9'd67,-10'd334};
ram[57206] = {9'd70,-10'd330};
ram[57207] = {9'd73,-10'd327};
ram[57208] = {9'd76,-10'd324};
ram[57209] = {9'd80,-10'd321};
ram[57210] = {9'd83,-10'd318};
ram[57211] = {9'd86,-10'd315};
ram[57212] = {9'd89,-10'd312};
ram[57213] = {9'd92,-10'd308};
ram[57214] = {9'd95,-10'd305};
ram[57215] = {9'd98,-10'd302};
ram[57216] = {9'd98,-10'd302};
ram[57217] = {-9'd99,-10'd299};
ram[57218] = {-9'd96,-10'd296};
ram[57219] = {-9'd92,-10'd293};
ram[57220] = {-9'd89,-10'd290};
ram[57221] = {-9'd86,-10'd286};
ram[57222] = {-9'd83,-10'd283};
ram[57223] = {-9'd80,-10'd280};
ram[57224] = {-9'd77,-10'd277};
ram[57225] = {-9'd74,-10'd274};
ram[57226] = {-9'd70,-10'd271};
ram[57227] = {-9'd67,-10'd268};
ram[57228] = {-9'd64,-10'd264};
ram[57229] = {-9'd61,-10'd261};
ram[57230] = {-9'd58,-10'd258};
ram[57231] = {-9'd55,-10'd255};
ram[57232] = {-9'd52,-10'd252};
ram[57233] = {-9'd48,-10'd249};
ram[57234] = {-9'd45,-10'd246};
ram[57235] = {-9'd42,-10'd242};
ram[57236] = {-9'd39,-10'd239};
ram[57237] = {-9'd36,-10'd236};
ram[57238] = {-9'd33,-10'd233};
ram[57239] = {-9'd30,-10'd230};
ram[57240] = {-9'd26,-10'd227};
ram[57241] = {-9'd23,-10'd224};
ram[57242] = {-9'd20,-10'd220};
ram[57243] = {-9'd17,-10'd217};
ram[57244] = {-9'd14,-10'd214};
ram[57245] = {-9'd11,-10'd211};
ram[57246] = {-9'd8,-10'd208};
ram[57247] = {-9'd4,-10'd205};
ram[57248] = {-9'd1,-10'd202};
ram[57249] = {9'd2,-10'd198};
ram[57250] = {9'd5,-10'd195};
ram[57251] = {9'd8,-10'd192};
ram[57252] = {9'd11,-10'd189};
ram[57253] = {9'd14,-10'd186};
ram[57254] = {9'd18,-10'd183};
ram[57255] = {9'd21,-10'd180};
ram[57256] = {9'd24,-10'd176};
ram[57257] = {9'd27,-10'd173};
ram[57258] = {9'd30,-10'd170};
ram[57259] = {9'd33,-10'd167};
ram[57260] = {9'd36,-10'd164};
ram[57261] = {9'd40,-10'd161};
ram[57262] = {9'd43,-10'd158};
ram[57263] = {9'd46,-10'd154};
ram[57264] = {9'd49,-10'd151};
ram[57265] = {9'd52,-10'd148};
ram[57266] = {9'd55,-10'd145};
ram[57267] = {9'd58,-10'd142};
ram[57268] = {9'd62,-10'd139};
ram[57269] = {9'd65,-10'd136};
ram[57270] = {9'd68,-10'd132};
ram[57271] = {9'd71,-10'd129};
ram[57272] = {9'd74,-10'd126};
ram[57273] = {9'd77,-10'd123};
ram[57274] = {9'd80,-10'd120};
ram[57275] = {9'd84,-10'd117};
ram[57276] = {9'd87,-10'd114};
ram[57277] = {9'd90,-10'd110};
ram[57278] = {9'd93,-10'd107};
ram[57279] = {9'd96,-10'd104};
ram[57280] = {9'd99,-10'd101};
ram[57281] = {-9'd98,-10'd98};
ram[57282] = {-9'd95,-10'd95};
ram[57283] = {-9'd92,-10'd92};
ram[57284] = {-9'd88,-10'd88};
ram[57285] = {-9'd85,-10'd85};
ram[57286] = {-9'd82,-10'd82};
ram[57287] = {-9'd79,-10'd79};
ram[57288] = {-9'd76,-10'd76};
ram[57289] = {-9'd73,-10'd73};
ram[57290] = {-9'd70,-10'd70};
ram[57291] = {-9'd66,-10'd66};
ram[57292] = {-9'd63,-10'd63};
ram[57293] = {-9'd60,-10'd60};
ram[57294] = {-9'd57,-10'd57};
ram[57295] = {-9'd54,-10'd54};
ram[57296] = {-9'd51,-10'd51};
ram[57297] = {-9'd48,-10'd48};
ram[57298] = {-9'd44,-10'd44};
ram[57299] = {-9'd41,-10'd41};
ram[57300] = {-9'd38,-10'd38};
ram[57301] = {-9'd35,-10'd35};
ram[57302] = {-9'd32,-10'd32};
ram[57303] = {-9'd29,-10'd29};
ram[57304] = {-9'd26,-10'd26};
ram[57305] = {-9'd22,-10'd22};
ram[57306] = {-9'd19,-10'd19};
ram[57307] = {-9'd16,-10'd16};
ram[57308] = {-9'd13,-10'd13};
ram[57309] = {-9'd10,-10'd10};
ram[57310] = {-9'd7,-10'd7};
ram[57311] = {-9'd4,-10'd4};
ram[57312] = {9'd0,10'd0};
ram[57313] = {9'd3,10'd3};
ram[57314] = {9'd6,10'd6};
ram[57315] = {9'd9,10'd9};
ram[57316] = {9'd12,10'd12};
ram[57317] = {9'd15,10'd15};
ram[57318] = {9'd18,10'd18};
ram[57319] = {9'd21,10'd21};
ram[57320] = {9'd25,10'd25};
ram[57321] = {9'd28,10'd28};
ram[57322] = {9'd31,10'd31};
ram[57323] = {9'd34,10'd34};
ram[57324] = {9'd37,10'd37};
ram[57325] = {9'd40,10'd40};
ram[57326] = {9'd43,10'd43};
ram[57327] = {9'd47,10'd47};
ram[57328] = {9'd50,10'd50};
ram[57329] = {9'd53,10'd53};
ram[57330] = {9'd56,10'd56};
ram[57331] = {9'd59,10'd59};
ram[57332] = {9'd62,10'd62};
ram[57333] = {9'd65,10'd65};
ram[57334] = {9'd69,10'd69};
ram[57335] = {9'd72,10'd72};
ram[57336] = {9'd75,10'd75};
ram[57337] = {9'd78,10'd78};
ram[57338] = {9'd81,10'd81};
ram[57339] = {9'd84,10'd84};
ram[57340] = {9'd87,10'd87};
ram[57341] = {9'd91,10'd91};
ram[57342] = {9'd94,10'd94};
ram[57343] = {9'd97,10'd97};
ram[57344] = {9'd97,10'd97};
ram[57345] = {-9'd100,10'd100};
ram[57346] = {-9'd97,10'd103};
ram[57347] = {-9'd94,10'd106};
ram[57348] = {-9'd91,10'd109};
ram[57349] = {-9'd88,10'd113};
ram[57350] = {-9'd85,10'd116};
ram[57351] = {-9'd81,10'd119};
ram[57352] = {-9'd78,10'd122};
ram[57353] = {-9'd75,10'd125};
ram[57354] = {-9'd72,10'd128};
ram[57355] = {-9'd69,10'd131};
ram[57356] = {-9'd66,10'd135};
ram[57357] = {-9'd63,10'd138};
ram[57358] = {-9'd59,10'd141};
ram[57359] = {-9'd56,10'd144};
ram[57360] = {-9'd53,10'd147};
ram[57361] = {-9'd50,10'd150};
ram[57362] = {-9'd47,10'd153};
ram[57363] = {-9'd44,10'd157};
ram[57364] = {-9'd41,10'd160};
ram[57365] = {-9'd37,10'd163};
ram[57366] = {-9'd34,10'd166};
ram[57367] = {-9'd31,10'd169};
ram[57368] = {-9'd28,10'd172};
ram[57369] = {-9'd25,10'd175};
ram[57370] = {-9'd22,10'd179};
ram[57371] = {-9'd19,10'd182};
ram[57372] = {-9'd15,10'd185};
ram[57373] = {-9'd12,10'd188};
ram[57374] = {-9'd9,10'd191};
ram[57375] = {-9'd6,10'd194};
ram[57376] = {-9'd3,10'd197};
ram[57377] = {9'd0,10'd201};
ram[57378] = {9'd3,10'd204};
ram[57379] = {9'd7,10'd207};
ram[57380] = {9'd10,10'd210};
ram[57381] = {9'd13,10'd213};
ram[57382] = {9'd16,10'd216};
ram[57383] = {9'd19,10'd219};
ram[57384] = {9'd22,10'd223};
ram[57385] = {9'd25,10'd226};
ram[57386] = {9'd29,10'd229};
ram[57387] = {9'd32,10'd232};
ram[57388] = {9'd35,10'd235};
ram[57389] = {9'd38,10'd238};
ram[57390] = {9'd41,10'd241};
ram[57391] = {9'd44,10'd245};
ram[57392] = {9'd47,10'd248};
ram[57393] = {9'd51,10'd251};
ram[57394] = {9'd54,10'd254};
ram[57395] = {9'd57,10'd257};
ram[57396] = {9'd60,10'd260};
ram[57397] = {9'd63,10'd263};
ram[57398] = {9'd66,10'd267};
ram[57399] = {9'd69,10'd270};
ram[57400] = {9'd73,10'd273};
ram[57401] = {9'd76,10'd276};
ram[57402] = {9'd79,10'd279};
ram[57403] = {9'd82,10'd282};
ram[57404] = {9'd85,10'd285};
ram[57405] = {9'd88,10'd289};
ram[57406] = {9'd91,10'd292};
ram[57407] = {9'd95,10'd295};
ram[57408] = {9'd98,10'd298};
ram[57409] = {-9'd99,10'd301};
ram[57410] = {-9'd96,10'd304};
ram[57411] = {-9'd93,10'd307};
ram[57412] = {-9'd90,10'd311};
ram[57413] = {-9'd87,10'd314};
ram[57414] = {-9'd84,10'd317};
ram[57415] = {-9'd81,10'd320};
ram[57416] = {-9'd77,10'd323};
ram[57417] = {-9'd74,10'd326};
ram[57418] = {-9'd71,10'd329};
ram[57419] = {-9'd68,10'd333};
ram[57420] = {-9'd65,10'd336};
ram[57421] = {-9'd62,10'd339};
ram[57422] = {-9'd59,10'd342};
ram[57423] = {-9'd55,10'd345};
ram[57424] = {-9'd52,10'd348};
ram[57425] = {-9'd49,10'd351};
ram[57426] = {-9'd46,10'd354};
ram[57427] = {-9'd43,10'd358};
ram[57428] = {-9'd40,10'd361};
ram[57429] = {-9'd37,10'd364};
ram[57430] = {-9'd33,10'd367};
ram[57431] = {-9'd30,10'd370};
ram[57432] = {-9'd27,10'd373};
ram[57433] = {-9'd24,10'd376};
ram[57434] = {-9'd21,10'd380};
ram[57435] = {-9'd18,10'd383};
ram[57436] = {-9'd15,10'd386};
ram[57437] = {-9'd11,10'd389};
ram[57438] = {-9'd8,10'd392};
ram[57439] = {-9'd5,10'd395};
ram[57440] = {-9'd2,10'd398};
ram[57441] = {9'd1,-10'd399};
ram[57442] = {9'd4,-10'd396};
ram[57443] = {9'd7,-10'd393};
ram[57444] = {9'd10,-10'd390};
ram[57445] = {9'd14,-10'd387};
ram[57446] = {9'd17,-10'd384};
ram[57447] = {9'd20,-10'd381};
ram[57448] = {9'd23,-10'd377};
ram[57449] = {9'd26,-10'd374};
ram[57450] = {9'd29,-10'd371};
ram[57451] = {9'd32,-10'd368};
ram[57452] = {9'd36,-10'd365};
ram[57453] = {9'd39,-10'd362};
ram[57454] = {9'd42,-10'd359};
ram[57455] = {9'd45,-10'd355};
ram[57456] = {9'd48,-10'd352};
ram[57457] = {9'd51,-10'd349};
ram[57458] = {9'd54,-10'd346};
ram[57459] = {9'd58,-10'd343};
ram[57460] = {9'd61,-10'd340};
ram[57461] = {9'd64,-10'd337};
ram[57462] = {9'd67,-10'd334};
ram[57463] = {9'd70,-10'd330};
ram[57464] = {9'd73,-10'd327};
ram[57465] = {9'd76,-10'd324};
ram[57466] = {9'd80,-10'd321};
ram[57467] = {9'd83,-10'd318};
ram[57468] = {9'd86,-10'd315};
ram[57469] = {9'd89,-10'd312};
ram[57470] = {9'd92,-10'd308};
ram[57471] = {9'd95,-10'd305};
ram[57472] = {9'd95,-10'd305};
ram[57473] = {9'd98,-10'd302};
ram[57474] = {-9'd99,-10'd299};
ram[57475] = {-9'd96,-10'd296};
ram[57476] = {-9'd92,-10'd293};
ram[57477] = {-9'd89,-10'd290};
ram[57478] = {-9'd86,-10'd286};
ram[57479] = {-9'd83,-10'd283};
ram[57480] = {-9'd80,-10'd280};
ram[57481] = {-9'd77,-10'd277};
ram[57482] = {-9'd74,-10'd274};
ram[57483] = {-9'd70,-10'd271};
ram[57484] = {-9'd67,-10'd268};
ram[57485] = {-9'd64,-10'd264};
ram[57486] = {-9'd61,-10'd261};
ram[57487] = {-9'd58,-10'd258};
ram[57488] = {-9'd55,-10'd255};
ram[57489] = {-9'd52,-10'd252};
ram[57490] = {-9'd48,-10'd249};
ram[57491] = {-9'd45,-10'd246};
ram[57492] = {-9'd42,-10'd242};
ram[57493] = {-9'd39,-10'd239};
ram[57494] = {-9'd36,-10'd236};
ram[57495] = {-9'd33,-10'd233};
ram[57496] = {-9'd30,-10'd230};
ram[57497] = {-9'd26,-10'd227};
ram[57498] = {-9'd23,-10'd224};
ram[57499] = {-9'd20,-10'd220};
ram[57500] = {-9'd17,-10'd217};
ram[57501] = {-9'd14,-10'd214};
ram[57502] = {-9'd11,-10'd211};
ram[57503] = {-9'd8,-10'd208};
ram[57504] = {-9'd4,-10'd205};
ram[57505] = {-9'd1,-10'd202};
ram[57506] = {9'd2,-10'd198};
ram[57507] = {9'd5,-10'd195};
ram[57508] = {9'd8,-10'd192};
ram[57509] = {9'd11,-10'd189};
ram[57510] = {9'd14,-10'd186};
ram[57511] = {9'd18,-10'd183};
ram[57512] = {9'd21,-10'd180};
ram[57513] = {9'd24,-10'd176};
ram[57514] = {9'd27,-10'd173};
ram[57515] = {9'd30,-10'd170};
ram[57516] = {9'd33,-10'd167};
ram[57517] = {9'd36,-10'd164};
ram[57518] = {9'd40,-10'd161};
ram[57519] = {9'd43,-10'd158};
ram[57520] = {9'd46,-10'd154};
ram[57521] = {9'd49,-10'd151};
ram[57522] = {9'd52,-10'd148};
ram[57523] = {9'd55,-10'd145};
ram[57524] = {9'd58,-10'd142};
ram[57525] = {9'd62,-10'd139};
ram[57526] = {9'd65,-10'd136};
ram[57527] = {9'd68,-10'd132};
ram[57528] = {9'd71,-10'd129};
ram[57529] = {9'd74,-10'd126};
ram[57530] = {9'd77,-10'd123};
ram[57531] = {9'd80,-10'd120};
ram[57532] = {9'd84,-10'd117};
ram[57533] = {9'd87,-10'd114};
ram[57534] = {9'd90,-10'd110};
ram[57535] = {9'd93,-10'd107};
ram[57536] = {9'd96,-10'd104};
ram[57537] = {9'd99,-10'd101};
ram[57538] = {-9'd98,-10'd98};
ram[57539] = {-9'd95,-10'd95};
ram[57540] = {-9'd92,-10'd92};
ram[57541] = {-9'd88,-10'd88};
ram[57542] = {-9'd85,-10'd85};
ram[57543] = {-9'd82,-10'd82};
ram[57544] = {-9'd79,-10'd79};
ram[57545] = {-9'd76,-10'd76};
ram[57546] = {-9'd73,-10'd73};
ram[57547] = {-9'd70,-10'd70};
ram[57548] = {-9'd66,-10'd66};
ram[57549] = {-9'd63,-10'd63};
ram[57550] = {-9'd60,-10'd60};
ram[57551] = {-9'd57,-10'd57};
ram[57552] = {-9'd54,-10'd54};
ram[57553] = {-9'd51,-10'd51};
ram[57554] = {-9'd48,-10'd48};
ram[57555] = {-9'd44,-10'd44};
ram[57556] = {-9'd41,-10'd41};
ram[57557] = {-9'd38,-10'd38};
ram[57558] = {-9'd35,-10'd35};
ram[57559] = {-9'd32,-10'd32};
ram[57560] = {-9'd29,-10'd29};
ram[57561] = {-9'd26,-10'd26};
ram[57562] = {-9'd22,-10'd22};
ram[57563] = {-9'd19,-10'd19};
ram[57564] = {-9'd16,-10'd16};
ram[57565] = {-9'd13,-10'd13};
ram[57566] = {-9'd10,-10'd10};
ram[57567] = {-9'd7,-10'd7};
ram[57568] = {-9'd4,-10'd4};
ram[57569] = {9'd0,10'd0};
ram[57570] = {9'd3,10'd3};
ram[57571] = {9'd6,10'd6};
ram[57572] = {9'd9,10'd9};
ram[57573] = {9'd12,10'd12};
ram[57574] = {9'd15,10'd15};
ram[57575] = {9'd18,10'd18};
ram[57576] = {9'd21,10'd21};
ram[57577] = {9'd25,10'd25};
ram[57578] = {9'd28,10'd28};
ram[57579] = {9'd31,10'd31};
ram[57580] = {9'd34,10'd34};
ram[57581] = {9'd37,10'd37};
ram[57582] = {9'd40,10'd40};
ram[57583] = {9'd43,10'd43};
ram[57584] = {9'd47,10'd47};
ram[57585] = {9'd50,10'd50};
ram[57586] = {9'd53,10'd53};
ram[57587] = {9'd56,10'd56};
ram[57588] = {9'd59,10'd59};
ram[57589] = {9'd62,10'd62};
ram[57590] = {9'd65,10'd65};
ram[57591] = {9'd69,10'd69};
ram[57592] = {9'd72,10'd72};
ram[57593] = {9'd75,10'd75};
ram[57594] = {9'd78,10'd78};
ram[57595] = {9'd81,10'd81};
ram[57596] = {9'd84,10'd84};
ram[57597] = {9'd87,10'd87};
ram[57598] = {9'd91,10'd91};
ram[57599] = {9'd94,10'd94};
ram[57600] = {9'd94,10'd94};
ram[57601] = {9'd97,10'd97};
ram[57602] = {-9'd100,10'd100};
ram[57603] = {-9'd97,10'd103};
ram[57604] = {-9'd94,10'd106};
ram[57605] = {-9'd91,10'd109};
ram[57606] = {-9'd88,10'd113};
ram[57607] = {-9'd85,10'd116};
ram[57608] = {-9'd81,10'd119};
ram[57609] = {-9'd78,10'd122};
ram[57610] = {-9'd75,10'd125};
ram[57611] = {-9'd72,10'd128};
ram[57612] = {-9'd69,10'd131};
ram[57613] = {-9'd66,10'd135};
ram[57614] = {-9'd63,10'd138};
ram[57615] = {-9'd59,10'd141};
ram[57616] = {-9'd56,10'd144};
ram[57617] = {-9'd53,10'd147};
ram[57618] = {-9'd50,10'd150};
ram[57619] = {-9'd47,10'd153};
ram[57620] = {-9'd44,10'd157};
ram[57621] = {-9'd41,10'd160};
ram[57622] = {-9'd37,10'd163};
ram[57623] = {-9'd34,10'd166};
ram[57624] = {-9'd31,10'd169};
ram[57625] = {-9'd28,10'd172};
ram[57626] = {-9'd25,10'd175};
ram[57627] = {-9'd22,10'd179};
ram[57628] = {-9'd19,10'd182};
ram[57629] = {-9'd15,10'd185};
ram[57630] = {-9'd12,10'd188};
ram[57631] = {-9'd9,10'd191};
ram[57632] = {-9'd6,10'd194};
ram[57633] = {-9'd3,10'd197};
ram[57634] = {9'd0,10'd201};
ram[57635] = {9'd3,10'd204};
ram[57636] = {9'd7,10'd207};
ram[57637] = {9'd10,10'd210};
ram[57638] = {9'd13,10'd213};
ram[57639] = {9'd16,10'd216};
ram[57640] = {9'd19,10'd219};
ram[57641] = {9'd22,10'd223};
ram[57642] = {9'd25,10'd226};
ram[57643] = {9'd29,10'd229};
ram[57644] = {9'd32,10'd232};
ram[57645] = {9'd35,10'd235};
ram[57646] = {9'd38,10'd238};
ram[57647] = {9'd41,10'd241};
ram[57648] = {9'd44,10'd245};
ram[57649] = {9'd47,10'd248};
ram[57650] = {9'd51,10'd251};
ram[57651] = {9'd54,10'd254};
ram[57652] = {9'd57,10'd257};
ram[57653] = {9'd60,10'd260};
ram[57654] = {9'd63,10'd263};
ram[57655] = {9'd66,10'd267};
ram[57656] = {9'd69,10'd270};
ram[57657] = {9'd73,10'd273};
ram[57658] = {9'd76,10'd276};
ram[57659] = {9'd79,10'd279};
ram[57660] = {9'd82,10'd282};
ram[57661] = {9'd85,10'd285};
ram[57662] = {9'd88,10'd289};
ram[57663] = {9'd91,10'd292};
ram[57664] = {9'd95,10'd295};
ram[57665] = {9'd98,10'd298};
ram[57666] = {-9'd99,10'd301};
ram[57667] = {-9'd96,10'd304};
ram[57668] = {-9'd93,10'd307};
ram[57669] = {-9'd90,10'd311};
ram[57670] = {-9'd87,10'd314};
ram[57671] = {-9'd84,10'd317};
ram[57672] = {-9'd81,10'd320};
ram[57673] = {-9'd77,10'd323};
ram[57674] = {-9'd74,10'd326};
ram[57675] = {-9'd71,10'd329};
ram[57676] = {-9'd68,10'd333};
ram[57677] = {-9'd65,10'd336};
ram[57678] = {-9'd62,10'd339};
ram[57679] = {-9'd59,10'd342};
ram[57680] = {-9'd55,10'd345};
ram[57681] = {-9'd52,10'd348};
ram[57682] = {-9'd49,10'd351};
ram[57683] = {-9'd46,10'd354};
ram[57684] = {-9'd43,10'd358};
ram[57685] = {-9'd40,10'd361};
ram[57686] = {-9'd37,10'd364};
ram[57687] = {-9'd33,10'd367};
ram[57688] = {-9'd30,10'd370};
ram[57689] = {-9'd27,10'd373};
ram[57690] = {-9'd24,10'd376};
ram[57691] = {-9'd21,10'd380};
ram[57692] = {-9'd18,10'd383};
ram[57693] = {-9'd15,10'd386};
ram[57694] = {-9'd11,10'd389};
ram[57695] = {-9'd8,10'd392};
ram[57696] = {-9'd5,10'd395};
ram[57697] = {-9'd2,10'd398};
ram[57698] = {9'd1,-10'd399};
ram[57699] = {9'd4,-10'd396};
ram[57700] = {9'd7,-10'd393};
ram[57701] = {9'd10,-10'd390};
ram[57702] = {9'd14,-10'd387};
ram[57703] = {9'd17,-10'd384};
ram[57704] = {9'd20,-10'd381};
ram[57705] = {9'd23,-10'd377};
ram[57706] = {9'd26,-10'd374};
ram[57707] = {9'd29,-10'd371};
ram[57708] = {9'd32,-10'd368};
ram[57709] = {9'd36,-10'd365};
ram[57710] = {9'd39,-10'd362};
ram[57711] = {9'd42,-10'd359};
ram[57712] = {9'd45,-10'd355};
ram[57713] = {9'd48,-10'd352};
ram[57714] = {9'd51,-10'd349};
ram[57715] = {9'd54,-10'd346};
ram[57716] = {9'd58,-10'd343};
ram[57717] = {9'd61,-10'd340};
ram[57718] = {9'd64,-10'd337};
ram[57719] = {9'd67,-10'd334};
ram[57720] = {9'd70,-10'd330};
ram[57721] = {9'd73,-10'd327};
ram[57722] = {9'd76,-10'd324};
ram[57723] = {9'd80,-10'd321};
ram[57724] = {9'd83,-10'd318};
ram[57725] = {9'd86,-10'd315};
ram[57726] = {9'd89,-10'd312};
ram[57727] = {9'd92,-10'd308};
ram[57728] = {9'd92,-10'd308};
ram[57729] = {9'd95,-10'd305};
ram[57730] = {9'd98,-10'd302};
ram[57731] = {-9'd99,-10'd299};
ram[57732] = {-9'd96,-10'd296};
ram[57733] = {-9'd92,-10'd293};
ram[57734] = {-9'd89,-10'd290};
ram[57735] = {-9'd86,-10'd286};
ram[57736] = {-9'd83,-10'd283};
ram[57737] = {-9'd80,-10'd280};
ram[57738] = {-9'd77,-10'd277};
ram[57739] = {-9'd74,-10'd274};
ram[57740] = {-9'd70,-10'd271};
ram[57741] = {-9'd67,-10'd268};
ram[57742] = {-9'd64,-10'd264};
ram[57743] = {-9'd61,-10'd261};
ram[57744] = {-9'd58,-10'd258};
ram[57745] = {-9'd55,-10'd255};
ram[57746] = {-9'd52,-10'd252};
ram[57747] = {-9'd48,-10'd249};
ram[57748] = {-9'd45,-10'd246};
ram[57749] = {-9'd42,-10'd242};
ram[57750] = {-9'd39,-10'd239};
ram[57751] = {-9'd36,-10'd236};
ram[57752] = {-9'd33,-10'd233};
ram[57753] = {-9'd30,-10'd230};
ram[57754] = {-9'd26,-10'd227};
ram[57755] = {-9'd23,-10'd224};
ram[57756] = {-9'd20,-10'd220};
ram[57757] = {-9'd17,-10'd217};
ram[57758] = {-9'd14,-10'd214};
ram[57759] = {-9'd11,-10'd211};
ram[57760] = {-9'd8,-10'd208};
ram[57761] = {-9'd4,-10'd205};
ram[57762] = {-9'd1,-10'd202};
ram[57763] = {9'd2,-10'd198};
ram[57764] = {9'd5,-10'd195};
ram[57765] = {9'd8,-10'd192};
ram[57766] = {9'd11,-10'd189};
ram[57767] = {9'd14,-10'd186};
ram[57768] = {9'd18,-10'd183};
ram[57769] = {9'd21,-10'd180};
ram[57770] = {9'd24,-10'd176};
ram[57771] = {9'd27,-10'd173};
ram[57772] = {9'd30,-10'd170};
ram[57773] = {9'd33,-10'd167};
ram[57774] = {9'd36,-10'd164};
ram[57775] = {9'd40,-10'd161};
ram[57776] = {9'd43,-10'd158};
ram[57777] = {9'd46,-10'd154};
ram[57778] = {9'd49,-10'd151};
ram[57779] = {9'd52,-10'd148};
ram[57780] = {9'd55,-10'd145};
ram[57781] = {9'd58,-10'd142};
ram[57782] = {9'd62,-10'd139};
ram[57783] = {9'd65,-10'd136};
ram[57784] = {9'd68,-10'd132};
ram[57785] = {9'd71,-10'd129};
ram[57786] = {9'd74,-10'd126};
ram[57787] = {9'd77,-10'd123};
ram[57788] = {9'd80,-10'd120};
ram[57789] = {9'd84,-10'd117};
ram[57790] = {9'd87,-10'd114};
ram[57791] = {9'd90,-10'd110};
ram[57792] = {9'd93,-10'd107};
ram[57793] = {9'd96,-10'd104};
ram[57794] = {9'd99,-10'd101};
ram[57795] = {-9'd98,-10'd98};
ram[57796] = {-9'd95,-10'd95};
ram[57797] = {-9'd92,-10'd92};
ram[57798] = {-9'd88,-10'd88};
ram[57799] = {-9'd85,-10'd85};
ram[57800] = {-9'd82,-10'd82};
ram[57801] = {-9'd79,-10'd79};
ram[57802] = {-9'd76,-10'd76};
ram[57803] = {-9'd73,-10'd73};
ram[57804] = {-9'd70,-10'd70};
ram[57805] = {-9'd66,-10'd66};
ram[57806] = {-9'd63,-10'd63};
ram[57807] = {-9'd60,-10'd60};
ram[57808] = {-9'd57,-10'd57};
ram[57809] = {-9'd54,-10'd54};
ram[57810] = {-9'd51,-10'd51};
ram[57811] = {-9'd48,-10'd48};
ram[57812] = {-9'd44,-10'd44};
ram[57813] = {-9'd41,-10'd41};
ram[57814] = {-9'd38,-10'd38};
ram[57815] = {-9'd35,-10'd35};
ram[57816] = {-9'd32,-10'd32};
ram[57817] = {-9'd29,-10'd29};
ram[57818] = {-9'd26,-10'd26};
ram[57819] = {-9'd22,-10'd22};
ram[57820] = {-9'd19,-10'd19};
ram[57821] = {-9'd16,-10'd16};
ram[57822] = {-9'd13,-10'd13};
ram[57823] = {-9'd10,-10'd10};
ram[57824] = {-9'd7,-10'd7};
ram[57825] = {-9'd4,-10'd4};
ram[57826] = {9'd0,10'd0};
ram[57827] = {9'd3,10'd3};
ram[57828] = {9'd6,10'd6};
ram[57829] = {9'd9,10'd9};
ram[57830] = {9'd12,10'd12};
ram[57831] = {9'd15,10'd15};
ram[57832] = {9'd18,10'd18};
ram[57833] = {9'd21,10'd21};
ram[57834] = {9'd25,10'd25};
ram[57835] = {9'd28,10'd28};
ram[57836] = {9'd31,10'd31};
ram[57837] = {9'd34,10'd34};
ram[57838] = {9'd37,10'd37};
ram[57839] = {9'd40,10'd40};
ram[57840] = {9'd43,10'd43};
ram[57841] = {9'd47,10'd47};
ram[57842] = {9'd50,10'd50};
ram[57843] = {9'd53,10'd53};
ram[57844] = {9'd56,10'd56};
ram[57845] = {9'd59,10'd59};
ram[57846] = {9'd62,10'd62};
ram[57847] = {9'd65,10'd65};
ram[57848] = {9'd69,10'd69};
ram[57849] = {9'd72,10'd72};
ram[57850] = {9'd75,10'd75};
ram[57851] = {9'd78,10'd78};
ram[57852] = {9'd81,10'd81};
ram[57853] = {9'd84,10'd84};
ram[57854] = {9'd87,10'd87};
ram[57855] = {9'd91,10'd91};
ram[57856] = {9'd91,10'd91};
ram[57857] = {9'd94,10'd94};
ram[57858] = {9'd97,10'd97};
ram[57859] = {-9'd100,10'd100};
ram[57860] = {-9'd97,10'd103};
ram[57861] = {-9'd94,10'd106};
ram[57862] = {-9'd91,10'd109};
ram[57863] = {-9'd88,10'd113};
ram[57864] = {-9'd85,10'd116};
ram[57865] = {-9'd81,10'd119};
ram[57866] = {-9'd78,10'd122};
ram[57867] = {-9'd75,10'd125};
ram[57868] = {-9'd72,10'd128};
ram[57869] = {-9'd69,10'd131};
ram[57870] = {-9'd66,10'd135};
ram[57871] = {-9'd63,10'd138};
ram[57872] = {-9'd59,10'd141};
ram[57873] = {-9'd56,10'd144};
ram[57874] = {-9'd53,10'd147};
ram[57875] = {-9'd50,10'd150};
ram[57876] = {-9'd47,10'd153};
ram[57877] = {-9'd44,10'd157};
ram[57878] = {-9'd41,10'd160};
ram[57879] = {-9'd37,10'd163};
ram[57880] = {-9'd34,10'd166};
ram[57881] = {-9'd31,10'd169};
ram[57882] = {-9'd28,10'd172};
ram[57883] = {-9'd25,10'd175};
ram[57884] = {-9'd22,10'd179};
ram[57885] = {-9'd19,10'd182};
ram[57886] = {-9'd15,10'd185};
ram[57887] = {-9'd12,10'd188};
ram[57888] = {-9'd9,10'd191};
ram[57889] = {-9'd6,10'd194};
ram[57890] = {-9'd3,10'd197};
ram[57891] = {9'd0,10'd201};
ram[57892] = {9'd3,10'd204};
ram[57893] = {9'd7,10'd207};
ram[57894] = {9'd10,10'd210};
ram[57895] = {9'd13,10'd213};
ram[57896] = {9'd16,10'd216};
ram[57897] = {9'd19,10'd219};
ram[57898] = {9'd22,10'd223};
ram[57899] = {9'd25,10'd226};
ram[57900] = {9'd29,10'd229};
ram[57901] = {9'd32,10'd232};
ram[57902] = {9'd35,10'd235};
ram[57903] = {9'd38,10'd238};
ram[57904] = {9'd41,10'd241};
ram[57905] = {9'd44,10'd245};
ram[57906] = {9'd47,10'd248};
ram[57907] = {9'd51,10'd251};
ram[57908] = {9'd54,10'd254};
ram[57909] = {9'd57,10'd257};
ram[57910] = {9'd60,10'd260};
ram[57911] = {9'd63,10'd263};
ram[57912] = {9'd66,10'd267};
ram[57913] = {9'd69,10'd270};
ram[57914] = {9'd73,10'd273};
ram[57915] = {9'd76,10'd276};
ram[57916] = {9'd79,10'd279};
ram[57917] = {9'd82,10'd282};
ram[57918] = {9'd85,10'd285};
ram[57919] = {9'd88,10'd289};
ram[57920] = {9'd91,10'd292};
ram[57921] = {9'd95,10'd295};
ram[57922] = {9'd98,10'd298};
ram[57923] = {-9'd99,10'd301};
ram[57924] = {-9'd96,10'd304};
ram[57925] = {-9'd93,10'd307};
ram[57926] = {-9'd90,10'd311};
ram[57927] = {-9'd87,10'd314};
ram[57928] = {-9'd84,10'd317};
ram[57929] = {-9'd81,10'd320};
ram[57930] = {-9'd77,10'd323};
ram[57931] = {-9'd74,10'd326};
ram[57932] = {-9'd71,10'd329};
ram[57933] = {-9'd68,10'd333};
ram[57934] = {-9'd65,10'd336};
ram[57935] = {-9'd62,10'd339};
ram[57936] = {-9'd59,10'd342};
ram[57937] = {-9'd55,10'd345};
ram[57938] = {-9'd52,10'd348};
ram[57939] = {-9'd49,10'd351};
ram[57940] = {-9'd46,10'd354};
ram[57941] = {-9'd43,10'd358};
ram[57942] = {-9'd40,10'd361};
ram[57943] = {-9'd37,10'd364};
ram[57944] = {-9'd33,10'd367};
ram[57945] = {-9'd30,10'd370};
ram[57946] = {-9'd27,10'd373};
ram[57947] = {-9'd24,10'd376};
ram[57948] = {-9'd21,10'd380};
ram[57949] = {-9'd18,10'd383};
ram[57950] = {-9'd15,10'd386};
ram[57951] = {-9'd11,10'd389};
ram[57952] = {-9'd8,10'd392};
ram[57953] = {-9'd5,10'd395};
ram[57954] = {-9'd2,10'd398};
ram[57955] = {9'd1,-10'd399};
ram[57956] = {9'd4,-10'd396};
ram[57957] = {9'd7,-10'd393};
ram[57958] = {9'd10,-10'd390};
ram[57959] = {9'd14,-10'd387};
ram[57960] = {9'd17,-10'd384};
ram[57961] = {9'd20,-10'd381};
ram[57962] = {9'd23,-10'd377};
ram[57963] = {9'd26,-10'd374};
ram[57964] = {9'd29,-10'd371};
ram[57965] = {9'd32,-10'd368};
ram[57966] = {9'd36,-10'd365};
ram[57967] = {9'd39,-10'd362};
ram[57968] = {9'd42,-10'd359};
ram[57969] = {9'd45,-10'd355};
ram[57970] = {9'd48,-10'd352};
ram[57971] = {9'd51,-10'd349};
ram[57972] = {9'd54,-10'd346};
ram[57973] = {9'd58,-10'd343};
ram[57974] = {9'd61,-10'd340};
ram[57975] = {9'd64,-10'd337};
ram[57976] = {9'd67,-10'd334};
ram[57977] = {9'd70,-10'd330};
ram[57978] = {9'd73,-10'd327};
ram[57979] = {9'd76,-10'd324};
ram[57980] = {9'd80,-10'd321};
ram[57981] = {9'd83,-10'd318};
ram[57982] = {9'd86,-10'd315};
ram[57983] = {9'd89,-10'd312};
ram[57984] = {9'd89,-10'd312};
ram[57985] = {9'd92,-10'd308};
ram[57986] = {9'd95,-10'd305};
ram[57987] = {9'd98,-10'd302};
ram[57988] = {-9'd99,-10'd299};
ram[57989] = {-9'd96,-10'd296};
ram[57990] = {-9'd92,-10'd293};
ram[57991] = {-9'd89,-10'd290};
ram[57992] = {-9'd86,-10'd286};
ram[57993] = {-9'd83,-10'd283};
ram[57994] = {-9'd80,-10'd280};
ram[57995] = {-9'd77,-10'd277};
ram[57996] = {-9'd74,-10'd274};
ram[57997] = {-9'd70,-10'd271};
ram[57998] = {-9'd67,-10'd268};
ram[57999] = {-9'd64,-10'd264};
ram[58000] = {-9'd61,-10'd261};
ram[58001] = {-9'd58,-10'd258};
ram[58002] = {-9'd55,-10'd255};
ram[58003] = {-9'd52,-10'd252};
ram[58004] = {-9'd48,-10'd249};
ram[58005] = {-9'd45,-10'd246};
ram[58006] = {-9'd42,-10'd242};
ram[58007] = {-9'd39,-10'd239};
ram[58008] = {-9'd36,-10'd236};
ram[58009] = {-9'd33,-10'd233};
ram[58010] = {-9'd30,-10'd230};
ram[58011] = {-9'd26,-10'd227};
ram[58012] = {-9'd23,-10'd224};
ram[58013] = {-9'd20,-10'd220};
ram[58014] = {-9'd17,-10'd217};
ram[58015] = {-9'd14,-10'd214};
ram[58016] = {-9'd11,-10'd211};
ram[58017] = {-9'd8,-10'd208};
ram[58018] = {-9'd4,-10'd205};
ram[58019] = {-9'd1,-10'd202};
ram[58020] = {9'd2,-10'd198};
ram[58021] = {9'd5,-10'd195};
ram[58022] = {9'd8,-10'd192};
ram[58023] = {9'd11,-10'd189};
ram[58024] = {9'd14,-10'd186};
ram[58025] = {9'd18,-10'd183};
ram[58026] = {9'd21,-10'd180};
ram[58027] = {9'd24,-10'd176};
ram[58028] = {9'd27,-10'd173};
ram[58029] = {9'd30,-10'd170};
ram[58030] = {9'd33,-10'd167};
ram[58031] = {9'd36,-10'd164};
ram[58032] = {9'd40,-10'd161};
ram[58033] = {9'd43,-10'd158};
ram[58034] = {9'd46,-10'd154};
ram[58035] = {9'd49,-10'd151};
ram[58036] = {9'd52,-10'd148};
ram[58037] = {9'd55,-10'd145};
ram[58038] = {9'd58,-10'd142};
ram[58039] = {9'd62,-10'd139};
ram[58040] = {9'd65,-10'd136};
ram[58041] = {9'd68,-10'd132};
ram[58042] = {9'd71,-10'd129};
ram[58043] = {9'd74,-10'd126};
ram[58044] = {9'd77,-10'd123};
ram[58045] = {9'd80,-10'd120};
ram[58046] = {9'd84,-10'd117};
ram[58047] = {9'd87,-10'd114};
ram[58048] = {9'd90,-10'd110};
ram[58049] = {9'd93,-10'd107};
ram[58050] = {9'd96,-10'd104};
ram[58051] = {9'd99,-10'd101};
ram[58052] = {-9'd98,-10'd98};
ram[58053] = {-9'd95,-10'd95};
ram[58054] = {-9'd92,-10'd92};
ram[58055] = {-9'd88,-10'd88};
ram[58056] = {-9'd85,-10'd85};
ram[58057] = {-9'd82,-10'd82};
ram[58058] = {-9'd79,-10'd79};
ram[58059] = {-9'd76,-10'd76};
ram[58060] = {-9'd73,-10'd73};
ram[58061] = {-9'd70,-10'd70};
ram[58062] = {-9'd66,-10'd66};
ram[58063] = {-9'd63,-10'd63};
ram[58064] = {-9'd60,-10'd60};
ram[58065] = {-9'd57,-10'd57};
ram[58066] = {-9'd54,-10'd54};
ram[58067] = {-9'd51,-10'd51};
ram[58068] = {-9'd48,-10'd48};
ram[58069] = {-9'd44,-10'd44};
ram[58070] = {-9'd41,-10'd41};
ram[58071] = {-9'd38,-10'd38};
ram[58072] = {-9'd35,-10'd35};
ram[58073] = {-9'd32,-10'd32};
ram[58074] = {-9'd29,-10'd29};
ram[58075] = {-9'd26,-10'd26};
ram[58076] = {-9'd22,-10'd22};
ram[58077] = {-9'd19,-10'd19};
ram[58078] = {-9'd16,-10'd16};
ram[58079] = {-9'd13,-10'd13};
ram[58080] = {-9'd10,-10'd10};
ram[58081] = {-9'd7,-10'd7};
ram[58082] = {-9'd4,-10'd4};
ram[58083] = {9'd0,10'd0};
ram[58084] = {9'd3,10'd3};
ram[58085] = {9'd6,10'd6};
ram[58086] = {9'd9,10'd9};
ram[58087] = {9'd12,10'd12};
ram[58088] = {9'd15,10'd15};
ram[58089] = {9'd18,10'd18};
ram[58090] = {9'd21,10'd21};
ram[58091] = {9'd25,10'd25};
ram[58092] = {9'd28,10'd28};
ram[58093] = {9'd31,10'd31};
ram[58094] = {9'd34,10'd34};
ram[58095] = {9'd37,10'd37};
ram[58096] = {9'd40,10'd40};
ram[58097] = {9'd43,10'd43};
ram[58098] = {9'd47,10'd47};
ram[58099] = {9'd50,10'd50};
ram[58100] = {9'd53,10'd53};
ram[58101] = {9'd56,10'd56};
ram[58102] = {9'd59,10'd59};
ram[58103] = {9'd62,10'd62};
ram[58104] = {9'd65,10'd65};
ram[58105] = {9'd69,10'd69};
ram[58106] = {9'd72,10'd72};
ram[58107] = {9'd75,10'd75};
ram[58108] = {9'd78,10'd78};
ram[58109] = {9'd81,10'd81};
ram[58110] = {9'd84,10'd84};
ram[58111] = {9'd87,10'd87};
ram[58112] = {9'd87,10'd87};
ram[58113] = {9'd91,10'd91};
ram[58114] = {9'd94,10'd94};
ram[58115] = {9'd97,10'd97};
ram[58116] = {-9'd100,10'd100};
ram[58117] = {-9'd97,10'd103};
ram[58118] = {-9'd94,10'd106};
ram[58119] = {-9'd91,10'd109};
ram[58120] = {-9'd88,10'd113};
ram[58121] = {-9'd85,10'd116};
ram[58122] = {-9'd81,10'd119};
ram[58123] = {-9'd78,10'd122};
ram[58124] = {-9'd75,10'd125};
ram[58125] = {-9'd72,10'd128};
ram[58126] = {-9'd69,10'd131};
ram[58127] = {-9'd66,10'd135};
ram[58128] = {-9'd63,10'd138};
ram[58129] = {-9'd59,10'd141};
ram[58130] = {-9'd56,10'd144};
ram[58131] = {-9'd53,10'd147};
ram[58132] = {-9'd50,10'd150};
ram[58133] = {-9'd47,10'd153};
ram[58134] = {-9'd44,10'd157};
ram[58135] = {-9'd41,10'd160};
ram[58136] = {-9'd37,10'd163};
ram[58137] = {-9'd34,10'd166};
ram[58138] = {-9'd31,10'd169};
ram[58139] = {-9'd28,10'd172};
ram[58140] = {-9'd25,10'd175};
ram[58141] = {-9'd22,10'd179};
ram[58142] = {-9'd19,10'd182};
ram[58143] = {-9'd15,10'd185};
ram[58144] = {-9'd12,10'd188};
ram[58145] = {-9'd9,10'd191};
ram[58146] = {-9'd6,10'd194};
ram[58147] = {-9'd3,10'd197};
ram[58148] = {9'd0,10'd201};
ram[58149] = {9'd3,10'd204};
ram[58150] = {9'd7,10'd207};
ram[58151] = {9'd10,10'd210};
ram[58152] = {9'd13,10'd213};
ram[58153] = {9'd16,10'd216};
ram[58154] = {9'd19,10'd219};
ram[58155] = {9'd22,10'd223};
ram[58156] = {9'd25,10'd226};
ram[58157] = {9'd29,10'd229};
ram[58158] = {9'd32,10'd232};
ram[58159] = {9'd35,10'd235};
ram[58160] = {9'd38,10'd238};
ram[58161] = {9'd41,10'd241};
ram[58162] = {9'd44,10'd245};
ram[58163] = {9'd47,10'd248};
ram[58164] = {9'd51,10'd251};
ram[58165] = {9'd54,10'd254};
ram[58166] = {9'd57,10'd257};
ram[58167] = {9'd60,10'd260};
ram[58168] = {9'd63,10'd263};
ram[58169] = {9'd66,10'd267};
ram[58170] = {9'd69,10'd270};
ram[58171] = {9'd73,10'd273};
ram[58172] = {9'd76,10'd276};
ram[58173] = {9'd79,10'd279};
ram[58174] = {9'd82,10'd282};
ram[58175] = {9'd85,10'd285};
ram[58176] = {9'd88,10'd289};
ram[58177] = {9'd91,10'd292};
ram[58178] = {9'd95,10'd295};
ram[58179] = {9'd98,10'd298};
ram[58180] = {-9'd99,10'd301};
ram[58181] = {-9'd96,10'd304};
ram[58182] = {-9'd93,10'd307};
ram[58183] = {-9'd90,10'd311};
ram[58184] = {-9'd87,10'd314};
ram[58185] = {-9'd84,10'd317};
ram[58186] = {-9'd81,10'd320};
ram[58187] = {-9'd77,10'd323};
ram[58188] = {-9'd74,10'd326};
ram[58189] = {-9'd71,10'd329};
ram[58190] = {-9'd68,10'd333};
ram[58191] = {-9'd65,10'd336};
ram[58192] = {-9'd62,10'd339};
ram[58193] = {-9'd59,10'd342};
ram[58194] = {-9'd55,10'd345};
ram[58195] = {-9'd52,10'd348};
ram[58196] = {-9'd49,10'd351};
ram[58197] = {-9'd46,10'd354};
ram[58198] = {-9'd43,10'd358};
ram[58199] = {-9'd40,10'd361};
ram[58200] = {-9'd37,10'd364};
ram[58201] = {-9'd33,10'd367};
ram[58202] = {-9'd30,10'd370};
ram[58203] = {-9'd27,10'd373};
ram[58204] = {-9'd24,10'd376};
ram[58205] = {-9'd21,10'd380};
ram[58206] = {-9'd18,10'd383};
ram[58207] = {-9'd15,10'd386};
ram[58208] = {-9'd11,10'd389};
ram[58209] = {-9'd8,10'd392};
ram[58210] = {-9'd5,10'd395};
ram[58211] = {-9'd2,10'd398};
ram[58212] = {9'd1,-10'd399};
ram[58213] = {9'd4,-10'd396};
ram[58214] = {9'd7,-10'd393};
ram[58215] = {9'd10,-10'd390};
ram[58216] = {9'd14,-10'd387};
ram[58217] = {9'd17,-10'd384};
ram[58218] = {9'd20,-10'd381};
ram[58219] = {9'd23,-10'd377};
ram[58220] = {9'd26,-10'd374};
ram[58221] = {9'd29,-10'd371};
ram[58222] = {9'd32,-10'd368};
ram[58223] = {9'd36,-10'd365};
ram[58224] = {9'd39,-10'd362};
ram[58225] = {9'd42,-10'd359};
ram[58226] = {9'd45,-10'd355};
ram[58227] = {9'd48,-10'd352};
ram[58228] = {9'd51,-10'd349};
ram[58229] = {9'd54,-10'd346};
ram[58230] = {9'd58,-10'd343};
ram[58231] = {9'd61,-10'd340};
ram[58232] = {9'd64,-10'd337};
ram[58233] = {9'd67,-10'd334};
ram[58234] = {9'd70,-10'd330};
ram[58235] = {9'd73,-10'd327};
ram[58236] = {9'd76,-10'd324};
ram[58237] = {9'd80,-10'd321};
ram[58238] = {9'd83,-10'd318};
ram[58239] = {9'd86,-10'd315};
ram[58240] = {9'd86,-10'd315};
ram[58241] = {9'd89,-10'd312};
ram[58242] = {9'd92,-10'd308};
ram[58243] = {9'd95,-10'd305};
ram[58244] = {9'd98,-10'd302};
ram[58245] = {-9'd99,-10'd299};
ram[58246] = {-9'd96,-10'd296};
ram[58247] = {-9'd92,-10'd293};
ram[58248] = {-9'd89,-10'd290};
ram[58249] = {-9'd86,-10'd286};
ram[58250] = {-9'd83,-10'd283};
ram[58251] = {-9'd80,-10'd280};
ram[58252] = {-9'd77,-10'd277};
ram[58253] = {-9'd74,-10'd274};
ram[58254] = {-9'd70,-10'd271};
ram[58255] = {-9'd67,-10'd268};
ram[58256] = {-9'd64,-10'd264};
ram[58257] = {-9'd61,-10'd261};
ram[58258] = {-9'd58,-10'd258};
ram[58259] = {-9'd55,-10'd255};
ram[58260] = {-9'd52,-10'd252};
ram[58261] = {-9'd48,-10'd249};
ram[58262] = {-9'd45,-10'd246};
ram[58263] = {-9'd42,-10'd242};
ram[58264] = {-9'd39,-10'd239};
ram[58265] = {-9'd36,-10'd236};
ram[58266] = {-9'd33,-10'd233};
ram[58267] = {-9'd30,-10'd230};
ram[58268] = {-9'd26,-10'd227};
ram[58269] = {-9'd23,-10'd224};
ram[58270] = {-9'd20,-10'd220};
ram[58271] = {-9'd17,-10'd217};
ram[58272] = {-9'd14,-10'd214};
ram[58273] = {-9'd11,-10'd211};
ram[58274] = {-9'd8,-10'd208};
ram[58275] = {-9'd4,-10'd205};
ram[58276] = {-9'd1,-10'd202};
ram[58277] = {9'd2,-10'd198};
ram[58278] = {9'd5,-10'd195};
ram[58279] = {9'd8,-10'd192};
ram[58280] = {9'd11,-10'd189};
ram[58281] = {9'd14,-10'd186};
ram[58282] = {9'd18,-10'd183};
ram[58283] = {9'd21,-10'd180};
ram[58284] = {9'd24,-10'd176};
ram[58285] = {9'd27,-10'd173};
ram[58286] = {9'd30,-10'd170};
ram[58287] = {9'd33,-10'd167};
ram[58288] = {9'd36,-10'd164};
ram[58289] = {9'd40,-10'd161};
ram[58290] = {9'd43,-10'd158};
ram[58291] = {9'd46,-10'd154};
ram[58292] = {9'd49,-10'd151};
ram[58293] = {9'd52,-10'd148};
ram[58294] = {9'd55,-10'd145};
ram[58295] = {9'd58,-10'd142};
ram[58296] = {9'd62,-10'd139};
ram[58297] = {9'd65,-10'd136};
ram[58298] = {9'd68,-10'd132};
ram[58299] = {9'd71,-10'd129};
ram[58300] = {9'd74,-10'd126};
ram[58301] = {9'd77,-10'd123};
ram[58302] = {9'd80,-10'd120};
ram[58303] = {9'd84,-10'd117};
ram[58304] = {9'd87,-10'd114};
ram[58305] = {9'd90,-10'd110};
ram[58306] = {9'd93,-10'd107};
ram[58307] = {9'd96,-10'd104};
ram[58308] = {9'd99,-10'd101};
ram[58309] = {-9'd98,-10'd98};
ram[58310] = {-9'd95,-10'd95};
ram[58311] = {-9'd92,-10'd92};
ram[58312] = {-9'd88,-10'd88};
ram[58313] = {-9'd85,-10'd85};
ram[58314] = {-9'd82,-10'd82};
ram[58315] = {-9'd79,-10'd79};
ram[58316] = {-9'd76,-10'd76};
ram[58317] = {-9'd73,-10'd73};
ram[58318] = {-9'd70,-10'd70};
ram[58319] = {-9'd66,-10'd66};
ram[58320] = {-9'd63,-10'd63};
ram[58321] = {-9'd60,-10'd60};
ram[58322] = {-9'd57,-10'd57};
ram[58323] = {-9'd54,-10'd54};
ram[58324] = {-9'd51,-10'd51};
ram[58325] = {-9'd48,-10'd48};
ram[58326] = {-9'd44,-10'd44};
ram[58327] = {-9'd41,-10'd41};
ram[58328] = {-9'd38,-10'd38};
ram[58329] = {-9'd35,-10'd35};
ram[58330] = {-9'd32,-10'd32};
ram[58331] = {-9'd29,-10'd29};
ram[58332] = {-9'd26,-10'd26};
ram[58333] = {-9'd22,-10'd22};
ram[58334] = {-9'd19,-10'd19};
ram[58335] = {-9'd16,-10'd16};
ram[58336] = {-9'd13,-10'd13};
ram[58337] = {-9'd10,-10'd10};
ram[58338] = {-9'd7,-10'd7};
ram[58339] = {-9'd4,-10'd4};
ram[58340] = {9'd0,10'd0};
ram[58341] = {9'd3,10'd3};
ram[58342] = {9'd6,10'd6};
ram[58343] = {9'd9,10'd9};
ram[58344] = {9'd12,10'd12};
ram[58345] = {9'd15,10'd15};
ram[58346] = {9'd18,10'd18};
ram[58347] = {9'd21,10'd21};
ram[58348] = {9'd25,10'd25};
ram[58349] = {9'd28,10'd28};
ram[58350] = {9'd31,10'd31};
ram[58351] = {9'd34,10'd34};
ram[58352] = {9'd37,10'd37};
ram[58353] = {9'd40,10'd40};
ram[58354] = {9'd43,10'd43};
ram[58355] = {9'd47,10'd47};
ram[58356] = {9'd50,10'd50};
ram[58357] = {9'd53,10'd53};
ram[58358] = {9'd56,10'd56};
ram[58359] = {9'd59,10'd59};
ram[58360] = {9'd62,10'd62};
ram[58361] = {9'd65,10'd65};
ram[58362] = {9'd69,10'd69};
ram[58363] = {9'd72,10'd72};
ram[58364] = {9'd75,10'd75};
ram[58365] = {9'd78,10'd78};
ram[58366] = {9'd81,10'd81};
ram[58367] = {9'd84,10'd84};
ram[58368] = {9'd84,10'd84};
ram[58369] = {9'd87,10'd87};
ram[58370] = {9'd91,10'd91};
ram[58371] = {9'd94,10'd94};
ram[58372] = {9'd97,10'd97};
ram[58373] = {-9'd100,10'd100};
ram[58374] = {-9'd97,10'd103};
ram[58375] = {-9'd94,10'd106};
ram[58376] = {-9'd91,10'd109};
ram[58377] = {-9'd88,10'd113};
ram[58378] = {-9'd85,10'd116};
ram[58379] = {-9'd81,10'd119};
ram[58380] = {-9'd78,10'd122};
ram[58381] = {-9'd75,10'd125};
ram[58382] = {-9'd72,10'd128};
ram[58383] = {-9'd69,10'd131};
ram[58384] = {-9'd66,10'd135};
ram[58385] = {-9'd63,10'd138};
ram[58386] = {-9'd59,10'd141};
ram[58387] = {-9'd56,10'd144};
ram[58388] = {-9'd53,10'd147};
ram[58389] = {-9'd50,10'd150};
ram[58390] = {-9'd47,10'd153};
ram[58391] = {-9'd44,10'd157};
ram[58392] = {-9'd41,10'd160};
ram[58393] = {-9'd37,10'd163};
ram[58394] = {-9'd34,10'd166};
ram[58395] = {-9'd31,10'd169};
ram[58396] = {-9'd28,10'd172};
ram[58397] = {-9'd25,10'd175};
ram[58398] = {-9'd22,10'd179};
ram[58399] = {-9'd19,10'd182};
ram[58400] = {-9'd15,10'd185};
ram[58401] = {-9'd12,10'd188};
ram[58402] = {-9'd9,10'd191};
ram[58403] = {-9'd6,10'd194};
ram[58404] = {-9'd3,10'd197};
ram[58405] = {9'd0,10'd201};
ram[58406] = {9'd3,10'd204};
ram[58407] = {9'd7,10'd207};
ram[58408] = {9'd10,10'd210};
ram[58409] = {9'd13,10'd213};
ram[58410] = {9'd16,10'd216};
ram[58411] = {9'd19,10'd219};
ram[58412] = {9'd22,10'd223};
ram[58413] = {9'd25,10'd226};
ram[58414] = {9'd29,10'd229};
ram[58415] = {9'd32,10'd232};
ram[58416] = {9'd35,10'd235};
ram[58417] = {9'd38,10'd238};
ram[58418] = {9'd41,10'd241};
ram[58419] = {9'd44,10'd245};
ram[58420] = {9'd47,10'd248};
ram[58421] = {9'd51,10'd251};
ram[58422] = {9'd54,10'd254};
ram[58423] = {9'd57,10'd257};
ram[58424] = {9'd60,10'd260};
ram[58425] = {9'd63,10'd263};
ram[58426] = {9'd66,10'd267};
ram[58427] = {9'd69,10'd270};
ram[58428] = {9'd73,10'd273};
ram[58429] = {9'd76,10'd276};
ram[58430] = {9'd79,10'd279};
ram[58431] = {9'd82,10'd282};
ram[58432] = {9'd85,10'd285};
ram[58433] = {9'd88,10'd289};
ram[58434] = {9'd91,10'd292};
ram[58435] = {9'd95,10'd295};
ram[58436] = {9'd98,10'd298};
ram[58437] = {-9'd99,10'd301};
ram[58438] = {-9'd96,10'd304};
ram[58439] = {-9'd93,10'd307};
ram[58440] = {-9'd90,10'd311};
ram[58441] = {-9'd87,10'd314};
ram[58442] = {-9'd84,10'd317};
ram[58443] = {-9'd81,10'd320};
ram[58444] = {-9'd77,10'd323};
ram[58445] = {-9'd74,10'd326};
ram[58446] = {-9'd71,10'd329};
ram[58447] = {-9'd68,10'd333};
ram[58448] = {-9'd65,10'd336};
ram[58449] = {-9'd62,10'd339};
ram[58450] = {-9'd59,10'd342};
ram[58451] = {-9'd55,10'd345};
ram[58452] = {-9'd52,10'd348};
ram[58453] = {-9'd49,10'd351};
ram[58454] = {-9'd46,10'd354};
ram[58455] = {-9'd43,10'd358};
ram[58456] = {-9'd40,10'd361};
ram[58457] = {-9'd37,10'd364};
ram[58458] = {-9'd33,10'd367};
ram[58459] = {-9'd30,10'd370};
ram[58460] = {-9'd27,10'd373};
ram[58461] = {-9'd24,10'd376};
ram[58462] = {-9'd21,10'd380};
ram[58463] = {-9'd18,10'd383};
ram[58464] = {-9'd15,10'd386};
ram[58465] = {-9'd11,10'd389};
ram[58466] = {-9'd8,10'd392};
ram[58467] = {-9'd5,10'd395};
ram[58468] = {-9'd2,10'd398};
ram[58469] = {9'd1,-10'd399};
ram[58470] = {9'd4,-10'd396};
ram[58471] = {9'd7,-10'd393};
ram[58472] = {9'd10,-10'd390};
ram[58473] = {9'd14,-10'd387};
ram[58474] = {9'd17,-10'd384};
ram[58475] = {9'd20,-10'd381};
ram[58476] = {9'd23,-10'd377};
ram[58477] = {9'd26,-10'd374};
ram[58478] = {9'd29,-10'd371};
ram[58479] = {9'd32,-10'd368};
ram[58480] = {9'd36,-10'd365};
ram[58481] = {9'd39,-10'd362};
ram[58482] = {9'd42,-10'd359};
ram[58483] = {9'd45,-10'd355};
ram[58484] = {9'd48,-10'd352};
ram[58485] = {9'd51,-10'd349};
ram[58486] = {9'd54,-10'd346};
ram[58487] = {9'd58,-10'd343};
ram[58488] = {9'd61,-10'd340};
ram[58489] = {9'd64,-10'd337};
ram[58490] = {9'd67,-10'd334};
ram[58491] = {9'd70,-10'd330};
ram[58492] = {9'd73,-10'd327};
ram[58493] = {9'd76,-10'd324};
ram[58494] = {9'd80,-10'd321};
ram[58495] = {9'd83,-10'd318};
ram[58496] = {9'd83,-10'd318};
ram[58497] = {9'd86,-10'd315};
ram[58498] = {9'd89,-10'd312};
ram[58499] = {9'd92,-10'd308};
ram[58500] = {9'd95,-10'd305};
ram[58501] = {9'd98,-10'd302};
ram[58502] = {-9'd99,-10'd299};
ram[58503] = {-9'd96,-10'd296};
ram[58504] = {-9'd92,-10'd293};
ram[58505] = {-9'd89,-10'd290};
ram[58506] = {-9'd86,-10'd286};
ram[58507] = {-9'd83,-10'd283};
ram[58508] = {-9'd80,-10'd280};
ram[58509] = {-9'd77,-10'd277};
ram[58510] = {-9'd74,-10'd274};
ram[58511] = {-9'd70,-10'd271};
ram[58512] = {-9'd67,-10'd268};
ram[58513] = {-9'd64,-10'd264};
ram[58514] = {-9'd61,-10'd261};
ram[58515] = {-9'd58,-10'd258};
ram[58516] = {-9'd55,-10'd255};
ram[58517] = {-9'd52,-10'd252};
ram[58518] = {-9'd48,-10'd249};
ram[58519] = {-9'd45,-10'd246};
ram[58520] = {-9'd42,-10'd242};
ram[58521] = {-9'd39,-10'd239};
ram[58522] = {-9'd36,-10'd236};
ram[58523] = {-9'd33,-10'd233};
ram[58524] = {-9'd30,-10'd230};
ram[58525] = {-9'd26,-10'd227};
ram[58526] = {-9'd23,-10'd224};
ram[58527] = {-9'd20,-10'd220};
ram[58528] = {-9'd17,-10'd217};
ram[58529] = {-9'd14,-10'd214};
ram[58530] = {-9'd11,-10'd211};
ram[58531] = {-9'd8,-10'd208};
ram[58532] = {-9'd4,-10'd205};
ram[58533] = {-9'd1,-10'd202};
ram[58534] = {9'd2,-10'd198};
ram[58535] = {9'd5,-10'd195};
ram[58536] = {9'd8,-10'd192};
ram[58537] = {9'd11,-10'd189};
ram[58538] = {9'd14,-10'd186};
ram[58539] = {9'd18,-10'd183};
ram[58540] = {9'd21,-10'd180};
ram[58541] = {9'd24,-10'd176};
ram[58542] = {9'd27,-10'd173};
ram[58543] = {9'd30,-10'd170};
ram[58544] = {9'd33,-10'd167};
ram[58545] = {9'd36,-10'd164};
ram[58546] = {9'd40,-10'd161};
ram[58547] = {9'd43,-10'd158};
ram[58548] = {9'd46,-10'd154};
ram[58549] = {9'd49,-10'd151};
ram[58550] = {9'd52,-10'd148};
ram[58551] = {9'd55,-10'd145};
ram[58552] = {9'd58,-10'd142};
ram[58553] = {9'd62,-10'd139};
ram[58554] = {9'd65,-10'd136};
ram[58555] = {9'd68,-10'd132};
ram[58556] = {9'd71,-10'd129};
ram[58557] = {9'd74,-10'd126};
ram[58558] = {9'd77,-10'd123};
ram[58559] = {9'd80,-10'd120};
ram[58560] = {9'd84,-10'd117};
ram[58561] = {9'd87,-10'd114};
ram[58562] = {9'd90,-10'd110};
ram[58563] = {9'd93,-10'd107};
ram[58564] = {9'd96,-10'd104};
ram[58565] = {9'd99,-10'd101};
ram[58566] = {-9'd98,-10'd98};
ram[58567] = {-9'd95,-10'd95};
ram[58568] = {-9'd92,-10'd92};
ram[58569] = {-9'd88,-10'd88};
ram[58570] = {-9'd85,-10'd85};
ram[58571] = {-9'd82,-10'd82};
ram[58572] = {-9'd79,-10'd79};
ram[58573] = {-9'd76,-10'd76};
ram[58574] = {-9'd73,-10'd73};
ram[58575] = {-9'd70,-10'd70};
ram[58576] = {-9'd66,-10'd66};
ram[58577] = {-9'd63,-10'd63};
ram[58578] = {-9'd60,-10'd60};
ram[58579] = {-9'd57,-10'd57};
ram[58580] = {-9'd54,-10'd54};
ram[58581] = {-9'd51,-10'd51};
ram[58582] = {-9'd48,-10'd48};
ram[58583] = {-9'd44,-10'd44};
ram[58584] = {-9'd41,-10'd41};
ram[58585] = {-9'd38,-10'd38};
ram[58586] = {-9'd35,-10'd35};
ram[58587] = {-9'd32,-10'd32};
ram[58588] = {-9'd29,-10'd29};
ram[58589] = {-9'd26,-10'd26};
ram[58590] = {-9'd22,-10'd22};
ram[58591] = {-9'd19,-10'd19};
ram[58592] = {-9'd16,-10'd16};
ram[58593] = {-9'd13,-10'd13};
ram[58594] = {-9'd10,-10'd10};
ram[58595] = {-9'd7,-10'd7};
ram[58596] = {-9'd4,-10'd4};
ram[58597] = {9'd0,10'd0};
ram[58598] = {9'd3,10'd3};
ram[58599] = {9'd6,10'd6};
ram[58600] = {9'd9,10'd9};
ram[58601] = {9'd12,10'd12};
ram[58602] = {9'd15,10'd15};
ram[58603] = {9'd18,10'd18};
ram[58604] = {9'd21,10'd21};
ram[58605] = {9'd25,10'd25};
ram[58606] = {9'd28,10'd28};
ram[58607] = {9'd31,10'd31};
ram[58608] = {9'd34,10'd34};
ram[58609] = {9'd37,10'd37};
ram[58610] = {9'd40,10'd40};
ram[58611] = {9'd43,10'd43};
ram[58612] = {9'd47,10'd47};
ram[58613] = {9'd50,10'd50};
ram[58614] = {9'd53,10'd53};
ram[58615] = {9'd56,10'd56};
ram[58616] = {9'd59,10'd59};
ram[58617] = {9'd62,10'd62};
ram[58618] = {9'd65,10'd65};
ram[58619] = {9'd69,10'd69};
ram[58620] = {9'd72,10'd72};
ram[58621] = {9'd75,10'd75};
ram[58622] = {9'd78,10'd78};
ram[58623] = {9'd81,10'd81};
ram[58624] = {9'd81,10'd81};
ram[58625] = {9'd84,10'd84};
ram[58626] = {9'd87,10'd87};
ram[58627] = {9'd91,10'd91};
ram[58628] = {9'd94,10'd94};
ram[58629] = {9'd97,10'd97};
ram[58630] = {-9'd100,10'd100};
ram[58631] = {-9'd97,10'd103};
ram[58632] = {-9'd94,10'd106};
ram[58633] = {-9'd91,10'd109};
ram[58634] = {-9'd88,10'd113};
ram[58635] = {-9'd85,10'd116};
ram[58636] = {-9'd81,10'd119};
ram[58637] = {-9'd78,10'd122};
ram[58638] = {-9'd75,10'd125};
ram[58639] = {-9'd72,10'd128};
ram[58640] = {-9'd69,10'd131};
ram[58641] = {-9'd66,10'd135};
ram[58642] = {-9'd63,10'd138};
ram[58643] = {-9'd59,10'd141};
ram[58644] = {-9'd56,10'd144};
ram[58645] = {-9'd53,10'd147};
ram[58646] = {-9'd50,10'd150};
ram[58647] = {-9'd47,10'd153};
ram[58648] = {-9'd44,10'd157};
ram[58649] = {-9'd41,10'd160};
ram[58650] = {-9'd37,10'd163};
ram[58651] = {-9'd34,10'd166};
ram[58652] = {-9'd31,10'd169};
ram[58653] = {-9'd28,10'd172};
ram[58654] = {-9'd25,10'd175};
ram[58655] = {-9'd22,10'd179};
ram[58656] = {-9'd19,10'd182};
ram[58657] = {-9'd15,10'd185};
ram[58658] = {-9'd12,10'd188};
ram[58659] = {-9'd9,10'd191};
ram[58660] = {-9'd6,10'd194};
ram[58661] = {-9'd3,10'd197};
ram[58662] = {9'd0,10'd201};
ram[58663] = {9'd3,10'd204};
ram[58664] = {9'd7,10'd207};
ram[58665] = {9'd10,10'd210};
ram[58666] = {9'd13,10'd213};
ram[58667] = {9'd16,10'd216};
ram[58668] = {9'd19,10'd219};
ram[58669] = {9'd22,10'd223};
ram[58670] = {9'd25,10'd226};
ram[58671] = {9'd29,10'd229};
ram[58672] = {9'd32,10'd232};
ram[58673] = {9'd35,10'd235};
ram[58674] = {9'd38,10'd238};
ram[58675] = {9'd41,10'd241};
ram[58676] = {9'd44,10'd245};
ram[58677] = {9'd47,10'd248};
ram[58678] = {9'd51,10'd251};
ram[58679] = {9'd54,10'd254};
ram[58680] = {9'd57,10'd257};
ram[58681] = {9'd60,10'd260};
ram[58682] = {9'd63,10'd263};
ram[58683] = {9'd66,10'd267};
ram[58684] = {9'd69,10'd270};
ram[58685] = {9'd73,10'd273};
ram[58686] = {9'd76,10'd276};
ram[58687] = {9'd79,10'd279};
ram[58688] = {9'd82,10'd282};
ram[58689] = {9'd85,10'd285};
ram[58690] = {9'd88,10'd289};
ram[58691] = {9'd91,10'd292};
ram[58692] = {9'd95,10'd295};
ram[58693] = {9'd98,10'd298};
ram[58694] = {-9'd99,10'd301};
ram[58695] = {-9'd96,10'd304};
ram[58696] = {-9'd93,10'd307};
ram[58697] = {-9'd90,10'd311};
ram[58698] = {-9'd87,10'd314};
ram[58699] = {-9'd84,10'd317};
ram[58700] = {-9'd81,10'd320};
ram[58701] = {-9'd77,10'd323};
ram[58702] = {-9'd74,10'd326};
ram[58703] = {-9'd71,10'd329};
ram[58704] = {-9'd68,10'd333};
ram[58705] = {-9'd65,10'd336};
ram[58706] = {-9'd62,10'd339};
ram[58707] = {-9'd59,10'd342};
ram[58708] = {-9'd55,10'd345};
ram[58709] = {-9'd52,10'd348};
ram[58710] = {-9'd49,10'd351};
ram[58711] = {-9'd46,10'd354};
ram[58712] = {-9'd43,10'd358};
ram[58713] = {-9'd40,10'd361};
ram[58714] = {-9'd37,10'd364};
ram[58715] = {-9'd33,10'd367};
ram[58716] = {-9'd30,10'd370};
ram[58717] = {-9'd27,10'd373};
ram[58718] = {-9'd24,10'd376};
ram[58719] = {-9'd21,10'd380};
ram[58720] = {-9'd18,10'd383};
ram[58721] = {-9'd15,10'd386};
ram[58722] = {-9'd11,10'd389};
ram[58723] = {-9'd8,10'd392};
ram[58724] = {-9'd5,10'd395};
ram[58725] = {-9'd2,10'd398};
ram[58726] = {9'd1,-10'd399};
ram[58727] = {9'd4,-10'd396};
ram[58728] = {9'd7,-10'd393};
ram[58729] = {9'd10,-10'd390};
ram[58730] = {9'd14,-10'd387};
ram[58731] = {9'd17,-10'd384};
ram[58732] = {9'd20,-10'd381};
ram[58733] = {9'd23,-10'd377};
ram[58734] = {9'd26,-10'd374};
ram[58735] = {9'd29,-10'd371};
ram[58736] = {9'd32,-10'd368};
ram[58737] = {9'd36,-10'd365};
ram[58738] = {9'd39,-10'd362};
ram[58739] = {9'd42,-10'd359};
ram[58740] = {9'd45,-10'd355};
ram[58741] = {9'd48,-10'd352};
ram[58742] = {9'd51,-10'd349};
ram[58743] = {9'd54,-10'd346};
ram[58744] = {9'd58,-10'd343};
ram[58745] = {9'd61,-10'd340};
ram[58746] = {9'd64,-10'd337};
ram[58747] = {9'd67,-10'd334};
ram[58748] = {9'd70,-10'd330};
ram[58749] = {9'd73,-10'd327};
ram[58750] = {9'd76,-10'd324};
ram[58751] = {9'd80,-10'd321};
ram[58752] = {9'd80,-10'd321};
ram[58753] = {9'd83,-10'd318};
ram[58754] = {9'd86,-10'd315};
ram[58755] = {9'd89,-10'd312};
ram[58756] = {9'd92,-10'd308};
ram[58757] = {9'd95,-10'd305};
ram[58758] = {9'd98,-10'd302};
ram[58759] = {-9'd99,-10'd299};
ram[58760] = {-9'd96,-10'd296};
ram[58761] = {-9'd92,-10'd293};
ram[58762] = {-9'd89,-10'd290};
ram[58763] = {-9'd86,-10'd286};
ram[58764] = {-9'd83,-10'd283};
ram[58765] = {-9'd80,-10'd280};
ram[58766] = {-9'd77,-10'd277};
ram[58767] = {-9'd74,-10'd274};
ram[58768] = {-9'd70,-10'd271};
ram[58769] = {-9'd67,-10'd268};
ram[58770] = {-9'd64,-10'd264};
ram[58771] = {-9'd61,-10'd261};
ram[58772] = {-9'd58,-10'd258};
ram[58773] = {-9'd55,-10'd255};
ram[58774] = {-9'd52,-10'd252};
ram[58775] = {-9'd48,-10'd249};
ram[58776] = {-9'd45,-10'd246};
ram[58777] = {-9'd42,-10'd242};
ram[58778] = {-9'd39,-10'd239};
ram[58779] = {-9'd36,-10'd236};
ram[58780] = {-9'd33,-10'd233};
ram[58781] = {-9'd30,-10'd230};
ram[58782] = {-9'd26,-10'd227};
ram[58783] = {-9'd23,-10'd224};
ram[58784] = {-9'd20,-10'd220};
ram[58785] = {-9'd17,-10'd217};
ram[58786] = {-9'd14,-10'd214};
ram[58787] = {-9'd11,-10'd211};
ram[58788] = {-9'd8,-10'd208};
ram[58789] = {-9'd4,-10'd205};
ram[58790] = {-9'd1,-10'd202};
ram[58791] = {9'd2,-10'd198};
ram[58792] = {9'd5,-10'd195};
ram[58793] = {9'd8,-10'd192};
ram[58794] = {9'd11,-10'd189};
ram[58795] = {9'd14,-10'd186};
ram[58796] = {9'd18,-10'd183};
ram[58797] = {9'd21,-10'd180};
ram[58798] = {9'd24,-10'd176};
ram[58799] = {9'd27,-10'd173};
ram[58800] = {9'd30,-10'd170};
ram[58801] = {9'd33,-10'd167};
ram[58802] = {9'd36,-10'd164};
ram[58803] = {9'd40,-10'd161};
ram[58804] = {9'd43,-10'd158};
ram[58805] = {9'd46,-10'd154};
ram[58806] = {9'd49,-10'd151};
ram[58807] = {9'd52,-10'd148};
ram[58808] = {9'd55,-10'd145};
ram[58809] = {9'd58,-10'd142};
ram[58810] = {9'd62,-10'd139};
ram[58811] = {9'd65,-10'd136};
ram[58812] = {9'd68,-10'd132};
ram[58813] = {9'd71,-10'd129};
ram[58814] = {9'd74,-10'd126};
ram[58815] = {9'd77,-10'd123};
ram[58816] = {9'd80,-10'd120};
ram[58817] = {9'd84,-10'd117};
ram[58818] = {9'd87,-10'd114};
ram[58819] = {9'd90,-10'd110};
ram[58820] = {9'd93,-10'd107};
ram[58821] = {9'd96,-10'd104};
ram[58822] = {9'd99,-10'd101};
ram[58823] = {-9'd98,-10'd98};
ram[58824] = {-9'd95,-10'd95};
ram[58825] = {-9'd92,-10'd92};
ram[58826] = {-9'd88,-10'd88};
ram[58827] = {-9'd85,-10'd85};
ram[58828] = {-9'd82,-10'd82};
ram[58829] = {-9'd79,-10'd79};
ram[58830] = {-9'd76,-10'd76};
ram[58831] = {-9'd73,-10'd73};
ram[58832] = {-9'd70,-10'd70};
ram[58833] = {-9'd66,-10'd66};
ram[58834] = {-9'd63,-10'd63};
ram[58835] = {-9'd60,-10'd60};
ram[58836] = {-9'd57,-10'd57};
ram[58837] = {-9'd54,-10'd54};
ram[58838] = {-9'd51,-10'd51};
ram[58839] = {-9'd48,-10'd48};
ram[58840] = {-9'd44,-10'd44};
ram[58841] = {-9'd41,-10'd41};
ram[58842] = {-9'd38,-10'd38};
ram[58843] = {-9'd35,-10'd35};
ram[58844] = {-9'd32,-10'd32};
ram[58845] = {-9'd29,-10'd29};
ram[58846] = {-9'd26,-10'd26};
ram[58847] = {-9'd22,-10'd22};
ram[58848] = {-9'd19,-10'd19};
ram[58849] = {-9'd16,-10'd16};
ram[58850] = {-9'd13,-10'd13};
ram[58851] = {-9'd10,-10'd10};
ram[58852] = {-9'd7,-10'd7};
ram[58853] = {-9'd4,-10'd4};
ram[58854] = {9'd0,10'd0};
ram[58855] = {9'd3,10'd3};
ram[58856] = {9'd6,10'd6};
ram[58857] = {9'd9,10'd9};
ram[58858] = {9'd12,10'd12};
ram[58859] = {9'd15,10'd15};
ram[58860] = {9'd18,10'd18};
ram[58861] = {9'd21,10'd21};
ram[58862] = {9'd25,10'd25};
ram[58863] = {9'd28,10'd28};
ram[58864] = {9'd31,10'd31};
ram[58865] = {9'd34,10'd34};
ram[58866] = {9'd37,10'd37};
ram[58867] = {9'd40,10'd40};
ram[58868] = {9'd43,10'd43};
ram[58869] = {9'd47,10'd47};
ram[58870] = {9'd50,10'd50};
ram[58871] = {9'd53,10'd53};
ram[58872] = {9'd56,10'd56};
ram[58873] = {9'd59,10'd59};
ram[58874] = {9'd62,10'd62};
ram[58875] = {9'd65,10'd65};
ram[58876] = {9'd69,10'd69};
ram[58877] = {9'd72,10'd72};
ram[58878] = {9'd75,10'd75};
ram[58879] = {9'd78,10'd78};
ram[58880] = {9'd78,10'd78};
ram[58881] = {9'd81,10'd81};
ram[58882] = {9'd84,10'd84};
ram[58883] = {9'd87,10'd87};
ram[58884] = {9'd91,10'd91};
ram[58885] = {9'd94,10'd94};
ram[58886] = {9'd97,10'd97};
ram[58887] = {-9'd100,10'd100};
ram[58888] = {-9'd97,10'd103};
ram[58889] = {-9'd94,10'd106};
ram[58890] = {-9'd91,10'd109};
ram[58891] = {-9'd88,10'd113};
ram[58892] = {-9'd85,10'd116};
ram[58893] = {-9'd81,10'd119};
ram[58894] = {-9'd78,10'd122};
ram[58895] = {-9'd75,10'd125};
ram[58896] = {-9'd72,10'd128};
ram[58897] = {-9'd69,10'd131};
ram[58898] = {-9'd66,10'd135};
ram[58899] = {-9'd63,10'd138};
ram[58900] = {-9'd59,10'd141};
ram[58901] = {-9'd56,10'd144};
ram[58902] = {-9'd53,10'd147};
ram[58903] = {-9'd50,10'd150};
ram[58904] = {-9'd47,10'd153};
ram[58905] = {-9'd44,10'd157};
ram[58906] = {-9'd41,10'd160};
ram[58907] = {-9'd37,10'd163};
ram[58908] = {-9'd34,10'd166};
ram[58909] = {-9'd31,10'd169};
ram[58910] = {-9'd28,10'd172};
ram[58911] = {-9'd25,10'd175};
ram[58912] = {-9'd22,10'd179};
ram[58913] = {-9'd19,10'd182};
ram[58914] = {-9'd15,10'd185};
ram[58915] = {-9'd12,10'd188};
ram[58916] = {-9'd9,10'd191};
ram[58917] = {-9'd6,10'd194};
ram[58918] = {-9'd3,10'd197};
ram[58919] = {9'd0,10'd201};
ram[58920] = {9'd3,10'd204};
ram[58921] = {9'd7,10'd207};
ram[58922] = {9'd10,10'd210};
ram[58923] = {9'd13,10'd213};
ram[58924] = {9'd16,10'd216};
ram[58925] = {9'd19,10'd219};
ram[58926] = {9'd22,10'd223};
ram[58927] = {9'd25,10'd226};
ram[58928] = {9'd29,10'd229};
ram[58929] = {9'd32,10'd232};
ram[58930] = {9'd35,10'd235};
ram[58931] = {9'd38,10'd238};
ram[58932] = {9'd41,10'd241};
ram[58933] = {9'd44,10'd245};
ram[58934] = {9'd47,10'd248};
ram[58935] = {9'd51,10'd251};
ram[58936] = {9'd54,10'd254};
ram[58937] = {9'd57,10'd257};
ram[58938] = {9'd60,10'd260};
ram[58939] = {9'd63,10'd263};
ram[58940] = {9'd66,10'd267};
ram[58941] = {9'd69,10'd270};
ram[58942] = {9'd73,10'd273};
ram[58943] = {9'd76,10'd276};
ram[58944] = {9'd79,10'd279};
ram[58945] = {9'd82,10'd282};
ram[58946] = {9'd85,10'd285};
ram[58947] = {9'd88,10'd289};
ram[58948] = {9'd91,10'd292};
ram[58949] = {9'd95,10'd295};
ram[58950] = {9'd98,10'd298};
ram[58951] = {-9'd99,10'd301};
ram[58952] = {-9'd96,10'd304};
ram[58953] = {-9'd93,10'd307};
ram[58954] = {-9'd90,10'd311};
ram[58955] = {-9'd87,10'd314};
ram[58956] = {-9'd84,10'd317};
ram[58957] = {-9'd81,10'd320};
ram[58958] = {-9'd77,10'd323};
ram[58959] = {-9'd74,10'd326};
ram[58960] = {-9'd71,10'd329};
ram[58961] = {-9'd68,10'd333};
ram[58962] = {-9'd65,10'd336};
ram[58963] = {-9'd62,10'd339};
ram[58964] = {-9'd59,10'd342};
ram[58965] = {-9'd55,10'd345};
ram[58966] = {-9'd52,10'd348};
ram[58967] = {-9'd49,10'd351};
ram[58968] = {-9'd46,10'd354};
ram[58969] = {-9'd43,10'd358};
ram[58970] = {-9'd40,10'd361};
ram[58971] = {-9'd37,10'd364};
ram[58972] = {-9'd33,10'd367};
ram[58973] = {-9'd30,10'd370};
ram[58974] = {-9'd27,10'd373};
ram[58975] = {-9'd24,10'd376};
ram[58976] = {-9'd21,10'd380};
ram[58977] = {-9'd18,10'd383};
ram[58978] = {-9'd15,10'd386};
ram[58979] = {-9'd11,10'd389};
ram[58980] = {-9'd8,10'd392};
ram[58981] = {-9'd5,10'd395};
ram[58982] = {-9'd2,10'd398};
ram[58983] = {9'd1,-10'd399};
ram[58984] = {9'd4,-10'd396};
ram[58985] = {9'd7,-10'd393};
ram[58986] = {9'd10,-10'd390};
ram[58987] = {9'd14,-10'd387};
ram[58988] = {9'd17,-10'd384};
ram[58989] = {9'd20,-10'd381};
ram[58990] = {9'd23,-10'd377};
ram[58991] = {9'd26,-10'd374};
ram[58992] = {9'd29,-10'd371};
ram[58993] = {9'd32,-10'd368};
ram[58994] = {9'd36,-10'd365};
ram[58995] = {9'd39,-10'd362};
ram[58996] = {9'd42,-10'd359};
ram[58997] = {9'd45,-10'd355};
ram[58998] = {9'd48,-10'd352};
ram[58999] = {9'd51,-10'd349};
ram[59000] = {9'd54,-10'd346};
ram[59001] = {9'd58,-10'd343};
ram[59002] = {9'd61,-10'd340};
ram[59003] = {9'd64,-10'd337};
ram[59004] = {9'd67,-10'd334};
ram[59005] = {9'd70,-10'd330};
ram[59006] = {9'd73,-10'd327};
ram[59007] = {9'd76,-10'd324};
ram[59008] = {9'd76,-10'd324};
ram[59009] = {9'd80,-10'd321};
ram[59010] = {9'd83,-10'd318};
ram[59011] = {9'd86,-10'd315};
ram[59012] = {9'd89,-10'd312};
ram[59013] = {9'd92,-10'd308};
ram[59014] = {9'd95,-10'd305};
ram[59015] = {9'd98,-10'd302};
ram[59016] = {-9'd99,-10'd299};
ram[59017] = {-9'd96,-10'd296};
ram[59018] = {-9'd92,-10'd293};
ram[59019] = {-9'd89,-10'd290};
ram[59020] = {-9'd86,-10'd286};
ram[59021] = {-9'd83,-10'd283};
ram[59022] = {-9'd80,-10'd280};
ram[59023] = {-9'd77,-10'd277};
ram[59024] = {-9'd74,-10'd274};
ram[59025] = {-9'd70,-10'd271};
ram[59026] = {-9'd67,-10'd268};
ram[59027] = {-9'd64,-10'd264};
ram[59028] = {-9'd61,-10'd261};
ram[59029] = {-9'd58,-10'd258};
ram[59030] = {-9'd55,-10'd255};
ram[59031] = {-9'd52,-10'd252};
ram[59032] = {-9'd48,-10'd249};
ram[59033] = {-9'd45,-10'd246};
ram[59034] = {-9'd42,-10'd242};
ram[59035] = {-9'd39,-10'd239};
ram[59036] = {-9'd36,-10'd236};
ram[59037] = {-9'd33,-10'd233};
ram[59038] = {-9'd30,-10'd230};
ram[59039] = {-9'd26,-10'd227};
ram[59040] = {-9'd23,-10'd224};
ram[59041] = {-9'd20,-10'd220};
ram[59042] = {-9'd17,-10'd217};
ram[59043] = {-9'd14,-10'd214};
ram[59044] = {-9'd11,-10'd211};
ram[59045] = {-9'd8,-10'd208};
ram[59046] = {-9'd4,-10'd205};
ram[59047] = {-9'd1,-10'd202};
ram[59048] = {9'd2,-10'd198};
ram[59049] = {9'd5,-10'd195};
ram[59050] = {9'd8,-10'd192};
ram[59051] = {9'd11,-10'd189};
ram[59052] = {9'd14,-10'd186};
ram[59053] = {9'd18,-10'd183};
ram[59054] = {9'd21,-10'd180};
ram[59055] = {9'd24,-10'd176};
ram[59056] = {9'd27,-10'd173};
ram[59057] = {9'd30,-10'd170};
ram[59058] = {9'd33,-10'd167};
ram[59059] = {9'd36,-10'd164};
ram[59060] = {9'd40,-10'd161};
ram[59061] = {9'd43,-10'd158};
ram[59062] = {9'd46,-10'd154};
ram[59063] = {9'd49,-10'd151};
ram[59064] = {9'd52,-10'd148};
ram[59065] = {9'd55,-10'd145};
ram[59066] = {9'd58,-10'd142};
ram[59067] = {9'd62,-10'd139};
ram[59068] = {9'd65,-10'd136};
ram[59069] = {9'd68,-10'd132};
ram[59070] = {9'd71,-10'd129};
ram[59071] = {9'd74,-10'd126};
ram[59072] = {9'd77,-10'd123};
ram[59073] = {9'd80,-10'd120};
ram[59074] = {9'd84,-10'd117};
ram[59075] = {9'd87,-10'd114};
ram[59076] = {9'd90,-10'd110};
ram[59077] = {9'd93,-10'd107};
ram[59078] = {9'd96,-10'd104};
ram[59079] = {9'd99,-10'd101};
ram[59080] = {-9'd98,-10'd98};
ram[59081] = {-9'd95,-10'd95};
ram[59082] = {-9'd92,-10'd92};
ram[59083] = {-9'd88,-10'd88};
ram[59084] = {-9'd85,-10'd85};
ram[59085] = {-9'd82,-10'd82};
ram[59086] = {-9'd79,-10'd79};
ram[59087] = {-9'd76,-10'd76};
ram[59088] = {-9'd73,-10'd73};
ram[59089] = {-9'd70,-10'd70};
ram[59090] = {-9'd66,-10'd66};
ram[59091] = {-9'd63,-10'd63};
ram[59092] = {-9'd60,-10'd60};
ram[59093] = {-9'd57,-10'd57};
ram[59094] = {-9'd54,-10'd54};
ram[59095] = {-9'd51,-10'd51};
ram[59096] = {-9'd48,-10'd48};
ram[59097] = {-9'd44,-10'd44};
ram[59098] = {-9'd41,-10'd41};
ram[59099] = {-9'd38,-10'd38};
ram[59100] = {-9'd35,-10'd35};
ram[59101] = {-9'd32,-10'd32};
ram[59102] = {-9'd29,-10'd29};
ram[59103] = {-9'd26,-10'd26};
ram[59104] = {-9'd22,-10'd22};
ram[59105] = {-9'd19,-10'd19};
ram[59106] = {-9'd16,-10'd16};
ram[59107] = {-9'd13,-10'd13};
ram[59108] = {-9'd10,-10'd10};
ram[59109] = {-9'd7,-10'd7};
ram[59110] = {-9'd4,-10'd4};
ram[59111] = {9'd0,10'd0};
ram[59112] = {9'd3,10'd3};
ram[59113] = {9'd6,10'd6};
ram[59114] = {9'd9,10'd9};
ram[59115] = {9'd12,10'd12};
ram[59116] = {9'd15,10'd15};
ram[59117] = {9'd18,10'd18};
ram[59118] = {9'd21,10'd21};
ram[59119] = {9'd25,10'd25};
ram[59120] = {9'd28,10'd28};
ram[59121] = {9'd31,10'd31};
ram[59122] = {9'd34,10'd34};
ram[59123] = {9'd37,10'd37};
ram[59124] = {9'd40,10'd40};
ram[59125] = {9'd43,10'd43};
ram[59126] = {9'd47,10'd47};
ram[59127] = {9'd50,10'd50};
ram[59128] = {9'd53,10'd53};
ram[59129] = {9'd56,10'd56};
ram[59130] = {9'd59,10'd59};
ram[59131] = {9'd62,10'd62};
ram[59132] = {9'd65,10'd65};
ram[59133] = {9'd69,10'd69};
ram[59134] = {9'd72,10'd72};
ram[59135] = {9'd75,10'd75};
ram[59136] = {9'd75,10'd75};
ram[59137] = {9'd78,10'd78};
ram[59138] = {9'd81,10'd81};
ram[59139] = {9'd84,10'd84};
ram[59140] = {9'd87,10'd87};
ram[59141] = {9'd91,10'd91};
ram[59142] = {9'd94,10'd94};
ram[59143] = {9'd97,10'd97};
ram[59144] = {-9'd100,10'd100};
ram[59145] = {-9'd97,10'd103};
ram[59146] = {-9'd94,10'd106};
ram[59147] = {-9'd91,10'd109};
ram[59148] = {-9'd88,10'd113};
ram[59149] = {-9'd85,10'd116};
ram[59150] = {-9'd81,10'd119};
ram[59151] = {-9'd78,10'd122};
ram[59152] = {-9'd75,10'd125};
ram[59153] = {-9'd72,10'd128};
ram[59154] = {-9'd69,10'd131};
ram[59155] = {-9'd66,10'd135};
ram[59156] = {-9'd63,10'd138};
ram[59157] = {-9'd59,10'd141};
ram[59158] = {-9'd56,10'd144};
ram[59159] = {-9'd53,10'd147};
ram[59160] = {-9'd50,10'd150};
ram[59161] = {-9'd47,10'd153};
ram[59162] = {-9'd44,10'd157};
ram[59163] = {-9'd41,10'd160};
ram[59164] = {-9'd37,10'd163};
ram[59165] = {-9'd34,10'd166};
ram[59166] = {-9'd31,10'd169};
ram[59167] = {-9'd28,10'd172};
ram[59168] = {-9'd25,10'd175};
ram[59169] = {-9'd22,10'd179};
ram[59170] = {-9'd19,10'd182};
ram[59171] = {-9'd15,10'd185};
ram[59172] = {-9'd12,10'd188};
ram[59173] = {-9'd9,10'd191};
ram[59174] = {-9'd6,10'd194};
ram[59175] = {-9'd3,10'd197};
ram[59176] = {9'd0,10'd201};
ram[59177] = {9'd3,10'd204};
ram[59178] = {9'd7,10'd207};
ram[59179] = {9'd10,10'd210};
ram[59180] = {9'd13,10'd213};
ram[59181] = {9'd16,10'd216};
ram[59182] = {9'd19,10'd219};
ram[59183] = {9'd22,10'd223};
ram[59184] = {9'd25,10'd226};
ram[59185] = {9'd29,10'd229};
ram[59186] = {9'd32,10'd232};
ram[59187] = {9'd35,10'd235};
ram[59188] = {9'd38,10'd238};
ram[59189] = {9'd41,10'd241};
ram[59190] = {9'd44,10'd245};
ram[59191] = {9'd47,10'd248};
ram[59192] = {9'd51,10'd251};
ram[59193] = {9'd54,10'd254};
ram[59194] = {9'd57,10'd257};
ram[59195] = {9'd60,10'd260};
ram[59196] = {9'd63,10'd263};
ram[59197] = {9'd66,10'd267};
ram[59198] = {9'd69,10'd270};
ram[59199] = {9'd73,10'd273};
ram[59200] = {9'd76,10'd276};
ram[59201] = {9'd79,10'd279};
ram[59202] = {9'd82,10'd282};
ram[59203] = {9'd85,10'd285};
ram[59204] = {9'd88,10'd289};
ram[59205] = {9'd91,10'd292};
ram[59206] = {9'd95,10'd295};
ram[59207] = {9'd98,10'd298};
ram[59208] = {-9'd99,10'd301};
ram[59209] = {-9'd96,10'd304};
ram[59210] = {-9'd93,10'd307};
ram[59211] = {-9'd90,10'd311};
ram[59212] = {-9'd87,10'd314};
ram[59213] = {-9'd84,10'd317};
ram[59214] = {-9'd81,10'd320};
ram[59215] = {-9'd77,10'd323};
ram[59216] = {-9'd74,10'd326};
ram[59217] = {-9'd71,10'd329};
ram[59218] = {-9'd68,10'd333};
ram[59219] = {-9'd65,10'd336};
ram[59220] = {-9'd62,10'd339};
ram[59221] = {-9'd59,10'd342};
ram[59222] = {-9'd55,10'd345};
ram[59223] = {-9'd52,10'd348};
ram[59224] = {-9'd49,10'd351};
ram[59225] = {-9'd46,10'd354};
ram[59226] = {-9'd43,10'd358};
ram[59227] = {-9'd40,10'd361};
ram[59228] = {-9'd37,10'd364};
ram[59229] = {-9'd33,10'd367};
ram[59230] = {-9'd30,10'd370};
ram[59231] = {-9'd27,10'd373};
ram[59232] = {-9'd24,10'd376};
ram[59233] = {-9'd21,10'd380};
ram[59234] = {-9'd18,10'd383};
ram[59235] = {-9'd15,10'd386};
ram[59236] = {-9'd11,10'd389};
ram[59237] = {-9'd8,10'd392};
ram[59238] = {-9'd5,10'd395};
ram[59239] = {-9'd2,10'd398};
ram[59240] = {9'd1,-10'd399};
ram[59241] = {9'd4,-10'd396};
ram[59242] = {9'd7,-10'd393};
ram[59243] = {9'd10,-10'd390};
ram[59244] = {9'd14,-10'd387};
ram[59245] = {9'd17,-10'd384};
ram[59246] = {9'd20,-10'd381};
ram[59247] = {9'd23,-10'd377};
ram[59248] = {9'd26,-10'd374};
ram[59249] = {9'd29,-10'd371};
ram[59250] = {9'd32,-10'd368};
ram[59251] = {9'd36,-10'd365};
ram[59252] = {9'd39,-10'd362};
ram[59253] = {9'd42,-10'd359};
ram[59254] = {9'd45,-10'd355};
ram[59255] = {9'd48,-10'd352};
ram[59256] = {9'd51,-10'd349};
ram[59257] = {9'd54,-10'd346};
ram[59258] = {9'd58,-10'd343};
ram[59259] = {9'd61,-10'd340};
ram[59260] = {9'd64,-10'd337};
ram[59261] = {9'd67,-10'd334};
ram[59262] = {9'd70,-10'd330};
ram[59263] = {9'd73,-10'd327};
ram[59264] = {9'd73,-10'd327};
ram[59265] = {9'd76,-10'd324};
ram[59266] = {9'd80,-10'd321};
ram[59267] = {9'd83,-10'd318};
ram[59268] = {9'd86,-10'd315};
ram[59269] = {9'd89,-10'd312};
ram[59270] = {9'd92,-10'd308};
ram[59271] = {9'd95,-10'd305};
ram[59272] = {9'd98,-10'd302};
ram[59273] = {-9'd99,-10'd299};
ram[59274] = {-9'd96,-10'd296};
ram[59275] = {-9'd92,-10'd293};
ram[59276] = {-9'd89,-10'd290};
ram[59277] = {-9'd86,-10'd286};
ram[59278] = {-9'd83,-10'd283};
ram[59279] = {-9'd80,-10'd280};
ram[59280] = {-9'd77,-10'd277};
ram[59281] = {-9'd74,-10'd274};
ram[59282] = {-9'd70,-10'd271};
ram[59283] = {-9'd67,-10'd268};
ram[59284] = {-9'd64,-10'd264};
ram[59285] = {-9'd61,-10'd261};
ram[59286] = {-9'd58,-10'd258};
ram[59287] = {-9'd55,-10'd255};
ram[59288] = {-9'd52,-10'd252};
ram[59289] = {-9'd48,-10'd249};
ram[59290] = {-9'd45,-10'd246};
ram[59291] = {-9'd42,-10'd242};
ram[59292] = {-9'd39,-10'd239};
ram[59293] = {-9'd36,-10'd236};
ram[59294] = {-9'd33,-10'd233};
ram[59295] = {-9'd30,-10'd230};
ram[59296] = {-9'd26,-10'd227};
ram[59297] = {-9'd23,-10'd224};
ram[59298] = {-9'd20,-10'd220};
ram[59299] = {-9'd17,-10'd217};
ram[59300] = {-9'd14,-10'd214};
ram[59301] = {-9'd11,-10'd211};
ram[59302] = {-9'd8,-10'd208};
ram[59303] = {-9'd4,-10'd205};
ram[59304] = {-9'd1,-10'd202};
ram[59305] = {9'd2,-10'd198};
ram[59306] = {9'd5,-10'd195};
ram[59307] = {9'd8,-10'd192};
ram[59308] = {9'd11,-10'd189};
ram[59309] = {9'd14,-10'd186};
ram[59310] = {9'd18,-10'd183};
ram[59311] = {9'd21,-10'd180};
ram[59312] = {9'd24,-10'd176};
ram[59313] = {9'd27,-10'd173};
ram[59314] = {9'd30,-10'd170};
ram[59315] = {9'd33,-10'd167};
ram[59316] = {9'd36,-10'd164};
ram[59317] = {9'd40,-10'd161};
ram[59318] = {9'd43,-10'd158};
ram[59319] = {9'd46,-10'd154};
ram[59320] = {9'd49,-10'd151};
ram[59321] = {9'd52,-10'd148};
ram[59322] = {9'd55,-10'd145};
ram[59323] = {9'd58,-10'd142};
ram[59324] = {9'd62,-10'd139};
ram[59325] = {9'd65,-10'd136};
ram[59326] = {9'd68,-10'd132};
ram[59327] = {9'd71,-10'd129};
ram[59328] = {9'd74,-10'd126};
ram[59329] = {9'd77,-10'd123};
ram[59330] = {9'd80,-10'd120};
ram[59331] = {9'd84,-10'd117};
ram[59332] = {9'd87,-10'd114};
ram[59333] = {9'd90,-10'd110};
ram[59334] = {9'd93,-10'd107};
ram[59335] = {9'd96,-10'd104};
ram[59336] = {9'd99,-10'd101};
ram[59337] = {-9'd98,-10'd98};
ram[59338] = {-9'd95,-10'd95};
ram[59339] = {-9'd92,-10'd92};
ram[59340] = {-9'd88,-10'd88};
ram[59341] = {-9'd85,-10'd85};
ram[59342] = {-9'd82,-10'd82};
ram[59343] = {-9'd79,-10'd79};
ram[59344] = {-9'd76,-10'd76};
ram[59345] = {-9'd73,-10'd73};
ram[59346] = {-9'd70,-10'd70};
ram[59347] = {-9'd66,-10'd66};
ram[59348] = {-9'd63,-10'd63};
ram[59349] = {-9'd60,-10'd60};
ram[59350] = {-9'd57,-10'd57};
ram[59351] = {-9'd54,-10'd54};
ram[59352] = {-9'd51,-10'd51};
ram[59353] = {-9'd48,-10'd48};
ram[59354] = {-9'd44,-10'd44};
ram[59355] = {-9'd41,-10'd41};
ram[59356] = {-9'd38,-10'd38};
ram[59357] = {-9'd35,-10'd35};
ram[59358] = {-9'd32,-10'd32};
ram[59359] = {-9'd29,-10'd29};
ram[59360] = {-9'd26,-10'd26};
ram[59361] = {-9'd22,-10'd22};
ram[59362] = {-9'd19,-10'd19};
ram[59363] = {-9'd16,-10'd16};
ram[59364] = {-9'd13,-10'd13};
ram[59365] = {-9'd10,-10'd10};
ram[59366] = {-9'd7,-10'd7};
ram[59367] = {-9'd4,-10'd4};
ram[59368] = {9'd0,10'd0};
ram[59369] = {9'd3,10'd3};
ram[59370] = {9'd6,10'd6};
ram[59371] = {9'd9,10'd9};
ram[59372] = {9'd12,10'd12};
ram[59373] = {9'd15,10'd15};
ram[59374] = {9'd18,10'd18};
ram[59375] = {9'd21,10'd21};
ram[59376] = {9'd25,10'd25};
ram[59377] = {9'd28,10'd28};
ram[59378] = {9'd31,10'd31};
ram[59379] = {9'd34,10'd34};
ram[59380] = {9'd37,10'd37};
ram[59381] = {9'd40,10'd40};
ram[59382] = {9'd43,10'd43};
ram[59383] = {9'd47,10'd47};
ram[59384] = {9'd50,10'd50};
ram[59385] = {9'd53,10'd53};
ram[59386] = {9'd56,10'd56};
ram[59387] = {9'd59,10'd59};
ram[59388] = {9'd62,10'd62};
ram[59389] = {9'd65,10'd65};
ram[59390] = {9'd69,10'd69};
ram[59391] = {9'd72,10'd72};
ram[59392] = {9'd72,10'd72};
ram[59393] = {9'd75,10'd75};
ram[59394] = {9'd78,10'd78};
ram[59395] = {9'd81,10'd81};
ram[59396] = {9'd84,10'd84};
ram[59397] = {9'd87,10'd87};
ram[59398] = {9'd91,10'd91};
ram[59399] = {9'd94,10'd94};
ram[59400] = {9'd97,10'd97};
ram[59401] = {-9'd100,10'd100};
ram[59402] = {-9'd97,10'd103};
ram[59403] = {-9'd94,10'd106};
ram[59404] = {-9'd91,10'd109};
ram[59405] = {-9'd88,10'd113};
ram[59406] = {-9'd85,10'd116};
ram[59407] = {-9'd81,10'd119};
ram[59408] = {-9'd78,10'd122};
ram[59409] = {-9'd75,10'd125};
ram[59410] = {-9'd72,10'd128};
ram[59411] = {-9'd69,10'd131};
ram[59412] = {-9'd66,10'd135};
ram[59413] = {-9'd63,10'd138};
ram[59414] = {-9'd59,10'd141};
ram[59415] = {-9'd56,10'd144};
ram[59416] = {-9'd53,10'd147};
ram[59417] = {-9'd50,10'd150};
ram[59418] = {-9'd47,10'd153};
ram[59419] = {-9'd44,10'd157};
ram[59420] = {-9'd41,10'd160};
ram[59421] = {-9'd37,10'd163};
ram[59422] = {-9'd34,10'd166};
ram[59423] = {-9'd31,10'd169};
ram[59424] = {-9'd28,10'd172};
ram[59425] = {-9'd25,10'd175};
ram[59426] = {-9'd22,10'd179};
ram[59427] = {-9'd19,10'd182};
ram[59428] = {-9'd15,10'd185};
ram[59429] = {-9'd12,10'd188};
ram[59430] = {-9'd9,10'd191};
ram[59431] = {-9'd6,10'd194};
ram[59432] = {-9'd3,10'd197};
ram[59433] = {9'd0,10'd201};
ram[59434] = {9'd3,10'd204};
ram[59435] = {9'd7,10'd207};
ram[59436] = {9'd10,10'd210};
ram[59437] = {9'd13,10'd213};
ram[59438] = {9'd16,10'd216};
ram[59439] = {9'd19,10'd219};
ram[59440] = {9'd22,10'd223};
ram[59441] = {9'd25,10'd226};
ram[59442] = {9'd29,10'd229};
ram[59443] = {9'd32,10'd232};
ram[59444] = {9'd35,10'd235};
ram[59445] = {9'd38,10'd238};
ram[59446] = {9'd41,10'd241};
ram[59447] = {9'd44,10'd245};
ram[59448] = {9'd47,10'd248};
ram[59449] = {9'd51,10'd251};
ram[59450] = {9'd54,10'd254};
ram[59451] = {9'd57,10'd257};
ram[59452] = {9'd60,10'd260};
ram[59453] = {9'd63,10'd263};
ram[59454] = {9'd66,10'd267};
ram[59455] = {9'd69,10'd270};
ram[59456] = {9'd73,10'd273};
ram[59457] = {9'd76,10'd276};
ram[59458] = {9'd79,10'd279};
ram[59459] = {9'd82,10'd282};
ram[59460] = {9'd85,10'd285};
ram[59461] = {9'd88,10'd289};
ram[59462] = {9'd91,10'd292};
ram[59463] = {9'd95,10'd295};
ram[59464] = {9'd98,10'd298};
ram[59465] = {-9'd99,10'd301};
ram[59466] = {-9'd96,10'd304};
ram[59467] = {-9'd93,10'd307};
ram[59468] = {-9'd90,10'd311};
ram[59469] = {-9'd87,10'd314};
ram[59470] = {-9'd84,10'd317};
ram[59471] = {-9'd81,10'd320};
ram[59472] = {-9'd77,10'd323};
ram[59473] = {-9'd74,10'd326};
ram[59474] = {-9'd71,10'd329};
ram[59475] = {-9'd68,10'd333};
ram[59476] = {-9'd65,10'd336};
ram[59477] = {-9'd62,10'd339};
ram[59478] = {-9'd59,10'd342};
ram[59479] = {-9'd55,10'd345};
ram[59480] = {-9'd52,10'd348};
ram[59481] = {-9'd49,10'd351};
ram[59482] = {-9'd46,10'd354};
ram[59483] = {-9'd43,10'd358};
ram[59484] = {-9'd40,10'd361};
ram[59485] = {-9'd37,10'd364};
ram[59486] = {-9'd33,10'd367};
ram[59487] = {-9'd30,10'd370};
ram[59488] = {-9'd27,10'd373};
ram[59489] = {-9'd24,10'd376};
ram[59490] = {-9'd21,10'd380};
ram[59491] = {-9'd18,10'd383};
ram[59492] = {-9'd15,10'd386};
ram[59493] = {-9'd11,10'd389};
ram[59494] = {-9'd8,10'd392};
ram[59495] = {-9'd5,10'd395};
ram[59496] = {-9'd2,10'd398};
ram[59497] = {9'd1,-10'd399};
ram[59498] = {9'd4,-10'd396};
ram[59499] = {9'd7,-10'd393};
ram[59500] = {9'd10,-10'd390};
ram[59501] = {9'd14,-10'd387};
ram[59502] = {9'd17,-10'd384};
ram[59503] = {9'd20,-10'd381};
ram[59504] = {9'd23,-10'd377};
ram[59505] = {9'd26,-10'd374};
ram[59506] = {9'd29,-10'd371};
ram[59507] = {9'd32,-10'd368};
ram[59508] = {9'd36,-10'd365};
ram[59509] = {9'd39,-10'd362};
ram[59510] = {9'd42,-10'd359};
ram[59511] = {9'd45,-10'd355};
ram[59512] = {9'd48,-10'd352};
ram[59513] = {9'd51,-10'd349};
ram[59514] = {9'd54,-10'd346};
ram[59515] = {9'd58,-10'd343};
ram[59516] = {9'd61,-10'd340};
ram[59517] = {9'd64,-10'd337};
ram[59518] = {9'd67,-10'd334};
ram[59519] = {9'd70,-10'd330};
ram[59520] = {9'd70,-10'd330};
ram[59521] = {9'd73,-10'd327};
ram[59522] = {9'd76,-10'd324};
ram[59523] = {9'd80,-10'd321};
ram[59524] = {9'd83,-10'd318};
ram[59525] = {9'd86,-10'd315};
ram[59526] = {9'd89,-10'd312};
ram[59527] = {9'd92,-10'd308};
ram[59528] = {9'd95,-10'd305};
ram[59529] = {9'd98,-10'd302};
ram[59530] = {-9'd99,-10'd299};
ram[59531] = {-9'd96,-10'd296};
ram[59532] = {-9'd92,-10'd293};
ram[59533] = {-9'd89,-10'd290};
ram[59534] = {-9'd86,-10'd286};
ram[59535] = {-9'd83,-10'd283};
ram[59536] = {-9'd80,-10'd280};
ram[59537] = {-9'd77,-10'd277};
ram[59538] = {-9'd74,-10'd274};
ram[59539] = {-9'd70,-10'd271};
ram[59540] = {-9'd67,-10'd268};
ram[59541] = {-9'd64,-10'd264};
ram[59542] = {-9'd61,-10'd261};
ram[59543] = {-9'd58,-10'd258};
ram[59544] = {-9'd55,-10'd255};
ram[59545] = {-9'd52,-10'd252};
ram[59546] = {-9'd48,-10'd249};
ram[59547] = {-9'd45,-10'd246};
ram[59548] = {-9'd42,-10'd242};
ram[59549] = {-9'd39,-10'd239};
ram[59550] = {-9'd36,-10'd236};
ram[59551] = {-9'd33,-10'd233};
ram[59552] = {-9'd30,-10'd230};
ram[59553] = {-9'd26,-10'd227};
ram[59554] = {-9'd23,-10'd224};
ram[59555] = {-9'd20,-10'd220};
ram[59556] = {-9'd17,-10'd217};
ram[59557] = {-9'd14,-10'd214};
ram[59558] = {-9'd11,-10'd211};
ram[59559] = {-9'd8,-10'd208};
ram[59560] = {-9'd4,-10'd205};
ram[59561] = {-9'd1,-10'd202};
ram[59562] = {9'd2,-10'd198};
ram[59563] = {9'd5,-10'd195};
ram[59564] = {9'd8,-10'd192};
ram[59565] = {9'd11,-10'd189};
ram[59566] = {9'd14,-10'd186};
ram[59567] = {9'd18,-10'd183};
ram[59568] = {9'd21,-10'd180};
ram[59569] = {9'd24,-10'd176};
ram[59570] = {9'd27,-10'd173};
ram[59571] = {9'd30,-10'd170};
ram[59572] = {9'd33,-10'd167};
ram[59573] = {9'd36,-10'd164};
ram[59574] = {9'd40,-10'd161};
ram[59575] = {9'd43,-10'd158};
ram[59576] = {9'd46,-10'd154};
ram[59577] = {9'd49,-10'd151};
ram[59578] = {9'd52,-10'd148};
ram[59579] = {9'd55,-10'd145};
ram[59580] = {9'd58,-10'd142};
ram[59581] = {9'd62,-10'd139};
ram[59582] = {9'd65,-10'd136};
ram[59583] = {9'd68,-10'd132};
ram[59584] = {9'd71,-10'd129};
ram[59585] = {9'd74,-10'd126};
ram[59586] = {9'd77,-10'd123};
ram[59587] = {9'd80,-10'd120};
ram[59588] = {9'd84,-10'd117};
ram[59589] = {9'd87,-10'd114};
ram[59590] = {9'd90,-10'd110};
ram[59591] = {9'd93,-10'd107};
ram[59592] = {9'd96,-10'd104};
ram[59593] = {9'd99,-10'd101};
ram[59594] = {-9'd98,-10'd98};
ram[59595] = {-9'd95,-10'd95};
ram[59596] = {-9'd92,-10'd92};
ram[59597] = {-9'd88,-10'd88};
ram[59598] = {-9'd85,-10'd85};
ram[59599] = {-9'd82,-10'd82};
ram[59600] = {-9'd79,-10'd79};
ram[59601] = {-9'd76,-10'd76};
ram[59602] = {-9'd73,-10'd73};
ram[59603] = {-9'd70,-10'd70};
ram[59604] = {-9'd66,-10'd66};
ram[59605] = {-9'd63,-10'd63};
ram[59606] = {-9'd60,-10'd60};
ram[59607] = {-9'd57,-10'd57};
ram[59608] = {-9'd54,-10'd54};
ram[59609] = {-9'd51,-10'd51};
ram[59610] = {-9'd48,-10'd48};
ram[59611] = {-9'd44,-10'd44};
ram[59612] = {-9'd41,-10'd41};
ram[59613] = {-9'd38,-10'd38};
ram[59614] = {-9'd35,-10'd35};
ram[59615] = {-9'd32,-10'd32};
ram[59616] = {-9'd29,-10'd29};
ram[59617] = {-9'd26,-10'd26};
ram[59618] = {-9'd22,-10'd22};
ram[59619] = {-9'd19,-10'd19};
ram[59620] = {-9'd16,-10'd16};
ram[59621] = {-9'd13,-10'd13};
ram[59622] = {-9'd10,-10'd10};
ram[59623] = {-9'd7,-10'd7};
ram[59624] = {-9'd4,-10'd4};
ram[59625] = {9'd0,10'd0};
ram[59626] = {9'd3,10'd3};
ram[59627] = {9'd6,10'd6};
ram[59628] = {9'd9,10'd9};
ram[59629] = {9'd12,10'd12};
ram[59630] = {9'd15,10'd15};
ram[59631] = {9'd18,10'd18};
ram[59632] = {9'd21,10'd21};
ram[59633] = {9'd25,10'd25};
ram[59634] = {9'd28,10'd28};
ram[59635] = {9'd31,10'd31};
ram[59636] = {9'd34,10'd34};
ram[59637] = {9'd37,10'd37};
ram[59638] = {9'd40,10'd40};
ram[59639] = {9'd43,10'd43};
ram[59640] = {9'd47,10'd47};
ram[59641] = {9'd50,10'd50};
ram[59642] = {9'd53,10'd53};
ram[59643] = {9'd56,10'd56};
ram[59644] = {9'd59,10'd59};
ram[59645] = {9'd62,10'd62};
ram[59646] = {9'd65,10'd65};
ram[59647] = {9'd69,10'd69};
ram[59648] = {9'd69,10'd69};
ram[59649] = {9'd72,10'd72};
ram[59650] = {9'd75,10'd75};
ram[59651] = {9'd78,10'd78};
ram[59652] = {9'd81,10'd81};
ram[59653] = {9'd84,10'd84};
ram[59654] = {9'd87,10'd87};
ram[59655] = {9'd91,10'd91};
ram[59656] = {9'd94,10'd94};
ram[59657] = {9'd97,10'd97};
ram[59658] = {-9'd100,10'd100};
ram[59659] = {-9'd97,10'd103};
ram[59660] = {-9'd94,10'd106};
ram[59661] = {-9'd91,10'd109};
ram[59662] = {-9'd88,10'd113};
ram[59663] = {-9'd85,10'd116};
ram[59664] = {-9'd81,10'd119};
ram[59665] = {-9'd78,10'd122};
ram[59666] = {-9'd75,10'd125};
ram[59667] = {-9'd72,10'd128};
ram[59668] = {-9'd69,10'd131};
ram[59669] = {-9'd66,10'd135};
ram[59670] = {-9'd63,10'd138};
ram[59671] = {-9'd59,10'd141};
ram[59672] = {-9'd56,10'd144};
ram[59673] = {-9'd53,10'd147};
ram[59674] = {-9'd50,10'd150};
ram[59675] = {-9'd47,10'd153};
ram[59676] = {-9'd44,10'd157};
ram[59677] = {-9'd41,10'd160};
ram[59678] = {-9'd37,10'd163};
ram[59679] = {-9'd34,10'd166};
ram[59680] = {-9'd31,10'd169};
ram[59681] = {-9'd28,10'd172};
ram[59682] = {-9'd25,10'd175};
ram[59683] = {-9'd22,10'd179};
ram[59684] = {-9'd19,10'd182};
ram[59685] = {-9'd15,10'd185};
ram[59686] = {-9'd12,10'd188};
ram[59687] = {-9'd9,10'd191};
ram[59688] = {-9'd6,10'd194};
ram[59689] = {-9'd3,10'd197};
ram[59690] = {9'd0,10'd201};
ram[59691] = {9'd3,10'd204};
ram[59692] = {9'd7,10'd207};
ram[59693] = {9'd10,10'd210};
ram[59694] = {9'd13,10'd213};
ram[59695] = {9'd16,10'd216};
ram[59696] = {9'd19,10'd219};
ram[59697] = {9'd22,10'd223};
ram[59698] = {9'd25,10'd226};
ram[59699] = {9'd29,10'd229};
ram[59700] = {9'd32,10'd232};
ram[59701] = {9'd35,10'd235};
ram[59702] = {9'd38,10'd238};
ram[59703] = {9'd41,10'd241};
ram[59704] = {9'd44,10'd245};
ram[59705] = {9'd47,10'd248};
ram[59706] = {9'd51,10'd251};
ram[59707] = {9'd54,10'd254};
ram[59708] = {9'd57,10'd257};
ram[59709] = {9'd60,10'd260};
ram[59710] = {9'd63,10'd263};
ram[59711] = {9'd66,10'd267};
ram[59712] = {9'd69,10'd270};
ram[59713] = {9'd73,10'd273};
ram[59714] = {9'd76,10'd276};
ram[59715] = {9'd79,10'd279};
ram[59716] = {9'd82,10'd282};
ram[59717] = {9'd85,10'd285};
ram[59718] = {9'd88,10'd289};
ram[59719] = {9'd91,10'd292};
ram[59720] = {9'd95,10'd295};
ram[59721] = {9'd98,10'd298};
ram[59722] = {-9'd99,10'd301};
ram[59723] = {-9'd96,10'd304};
ram[59724] = {-9'd93,10'd307};
ram[59725] = {-9'd90,10'd311};
ram[59726] = {-9'd87,10'd314};
ram[59727] = {-9'd84,10'd317};
ram[59728] = {-9'd81,10'd320};
ram[59729] = {-9'd77,10'd323};
ram[59730] = {-9'd74,10'd326};
ram[59731] = {-9'd71,10'd329};
ram[59732] = {-9'd68,10'd333};
ram[59733] = {-9'd65,10'd336};
ram[59734] = {-9'd62,10'd339};
ram[59735] = {-9'd59,10'd342};
ram[59736] = {-9'd55,10'd345};
ram[59737] = {-9'd52,10'd348};
ram[59738] = {-9'd49,10'd351};
ram[59739] = {-9'd46,10'd354};
ram[59740] = {-9'd43,10'd358};
ram[59741] = {-9'd40,10'd361};
ram[59742] = {-9'd37,10'd364};
ram[59743] = {-9'd33,10'd367};
ram[59744] = {-9'd30,10'd370};
ram[59745] = {-9'd27,10'd373};
ram[59746] = {-9'd24,10'd376};
ram[59747] = {-9'd21,10'd380};
ram[59748] = {-9'd18,10'd383};
ram[59749] = {-9'd15,10'd386};
ram[59750] = {-9'd11,10'd389};
ram[59751] = {-9'd8,10'd392};
ram[59752] = {-9'd5,10'd395};
ram[59753] = {-9'd2,10'd398};
ram[59754] = {9'd1,-10'd399};
ram[59755] = {9'd4,-10'd396};
ram[59756] = {9'd7,-10'd393};
ram[59757] = {9'd10,-10'd390};
ram[59758] = {9'd14,-10'd387};
ram[59759] = {9'd17,-10'd384};
ram[59760] = {9'd20,-10'd381};
ram[59761] = {9'd23,-10'd377};
ram[59762] = {9'd26,-10'd374};
ram[59763] = {9'd29,-10'd371};
ram[59764] = {9'd32,-10'd368};
ram[59765] = {9'd36,-10'd365};
ram[59766] = {9'd39,-10'd362};
ram[59767] = {9'd42,-10'd359};
ram[59768] = {9'd45,-10'd355};
ram[59769] = {9'd48,-10'd352};
ram[59770] = {9'd51,-10'd349};
ram[59771] = {9'd54,-10'd346};
ram[59772] = {9'd58,-10'd343};
ram[59773] = {9'd61,-10'd340};
ram[59774] = {9'd64,-10'd337};
ram[59775] = {9'd67,-10'd334};
ram[59776] = {9'd67,-10'd334};
ram[59777] = {9'd70,-10'd330};
ram[59778] = {9'd73,-10'd327};
ram[59779] = {9'd76,-10'd324};
ram[59780] = {9'd80,-10'd321};
ram[59781] = {9'd83,-10'd318};
ram[59782] = {9'd86,-10'd315};
ram[59783] = {9'd89,-10'd312};
ram[59784] = {9'd92,-10'd308};
ram[59785] = {9'd95,-10'd305};
ram[59786] = {9'd98,-10'd302};
ram[59787] = {-9'd99,-10'd299};
ram[59788] = {-9'd96,-10'd296};
ram[59789] = {-9'd92,-10'd293};
ram[59790] = {-9'd89,-10'd290};
ram[59791] = {-9'd86,-10'd286};
ram[59792] = {-9'd83,-10'd283};
ram[59793] = {-9'd80,-10'd280};
ram[59794] = {-9'd77,-10'd277};
ram[59795] = {-9'd74,-10'd274};
ram[59796] = {-9'd70,-10'd271};
ram[59797] = {-9'd67,-10'd268};
ram[59798] = {-9'd64,-10'd264};
ram[59799] = {-9'd61,-10'd261};
ram[59800] = {-9'd58,-10'd258};
ram[59801] = {-9'd55,-10'd255};
ram[59802] = {-9'd52,-10'd252};
ram[59803] = {-9'd48,-10'd249};
ram[59804] = {-9'd45,-10'd246};
ram[59805] = {-9'd42,-10'd242};
ram[59806] = {-9'd39,-10'd239};
ram[59807] = {-9'd36,-10'd236};
ram[59808] = {-9'd33,-10'd233};
ram[59809] = {-9'd30,-10'd230};
ram[59810] = {-9'd26,-10'd227};
ram[59811] = {-9'd23,-10'd224};
ram[59812] = {-9'd20,-10'd220};
ram[59813] = {-9'd17,-10'd217};
ram[59814] = {-9'd14,-10'd214};
ram[59815] = {-9'd11,-10'd211};
ram[59816] = {-9'd8,-10'd208};
ram[59817] = {-9'd4,-10'd205};
ram[59818] = {-9'd1,-10'd202};
ram[59819] = {9'd2,-10'd198};
ram[59820] = {9'd5,-10'd195};
ram[59821] = {9'd8,-10'd192};
ram[59822] = {9'd11,-10'd189};
ram[59823] = {9'd14,-10'd186};
ram[59824] = {9'd18,-10'd183};
ram[59825] = {9'd21,-10'd180};
ram[59826] = {9'd24,-10'd176};
ram[59827] = {9'd27,-10'd173};
ram[59828] = {9'd30,-10'd170};
ram[59829] = {9'd33,-10'd167};
ram[59830] = {9'd36,-10'd164};
ram[59831] = {9'd40,-10'd161};
ram[59832] = {9'd43,-10'd158};
ram[59833] = {9'd46,-10'd154};
ram[59834] = {9'd49,-10'd151};
ram[59835] = {9'd52,-10'd148};
ram[59836] = {9'd55,-10'd145};
ram[59837] = {9'd58,-10'd142};
ram[59838] = {9'd62,-10'd139};
ram[59839] = {9'd65,-10'd136};
ram[59840] = {9'd68,-10'd132};
ram[59841] = {9'd71,-10'd129};
ram[59842] = {9'd74,-10'd126};
ram[59843] = {9'd77,-10'd123};
ram[59844] = {9'd80,-10'd120};
ram[59845] = {9'd84,-10'd117};
ram[59846] = {9'd87,-10'd114};
ram[59847] = {9'd90,-10'd110};
ram[59848] = {9'd93,-10'd107};
ram[59849] = {9'd96,-10'd104};
ram[59850] = {9'd99,-10'd101};
ram[59851] = {-9'd98,-10'd98};
ram[59852] = {-9'd95,-10'd95};
ram[59853] = {-9'd92,-10'd92};
ram[59854] = {-9'd88,-10'd88};
ram[59855] = {-9'd85,-10'd85};
ram[59856] = {-9'd82,-10'd82};
ram[59857] = {-9'd79,-10'd79};
ram[59858] = {-9'd76,-10'd76};
ram[59859] = {-9'd73,-10'd73};
ram[59860] = {-9'd70,-10'd70};
ram[59861] = {-9'd66,-10'd66};
ram[59862] = {-9'd63,-10'd63};
ram[59863] = {-9'd60,-10'd60};
ram[59864] = {-9'd57,-10'd57};
ram[59865] = {-9'd54,-10'd54};
ram[59866] = {-9'd51,-10'd51};
ram[59867] = {-9'd48,-10'd48};
ram[59868] = {-9'd44,-10'd44};
ram[59869] = {-9'd41,-10'd41};
ram[59870] = {-9'd38,-10'd38};
ram[59871] = {-9'd35,-10'd35};
ram[59872] = {-9'd32,-10'd32};
ram[59873] = {-9'd29,-10'd29};
ram[59874] = {-9'd26,-10'd26};
ram[59875] = {-9'd22,-10'd22};
ram[59876] = {-9'd19,-10'd19};
ram[59877] = {-9'd16,-10'd16};
ram[59878] = {-9'd13,-10'd13};
ram[59879] = {-9'd10,-10'd10};
ram[59880] = {-9'd7,-10'd7};
ram[59881] = {-9'd4,-10'd4};
ram[59882] = {9'd0,10'd0};
ram[59883] = {9'd3,10'd3};
ram[59884] = {9'd6,10'd6};
ram[59885] = {9'd9,10'd9};
ram[59886] = {9'd12,10'd12};
ram[59887] = {9'd15,10'd15};
ram[59888] = {9'd18,10'd18};
ram[59889] = {9'd21,10'd21};
ram[59890] = {9'd25,10'd25};
ram[59891] = {9'd28,10'd28};
ram[59892] = {9'd31,10'd31};
ram[59893] = {9'd34,10'd34};
ram[59894] = {9'd37,10'd37};
ram[59895] = {9'd40,10'd40};
ram[59896] = {9'd43,10'd43};
ram[59897] = {9'd47,10'd47};
ram[59898] = {9'd50,10'd50};
ram[59899] = {9'd53,10'd53};
ram[59900] = {9'd56,10'd56};
ram[59901] = {9'd59,10'd59};
ram[59902] = {9'd62,10'd62};
ram[59903] = {9'd65,10'd65};
ram[59904] = {9'd65,10'd65};
ram[59905] = {9'd69,10'd69};
ram[59906] = {9'd72,10'd72};
ram[59907] = {9'd75,10'd75};
ram[59908] = {9'd78,10'd78};
ram[59909] = {9'd81,10'd81};
ram[59910] = {9'd84,10'd84};
ram[59911] = {9'd87,10'd87};
ram[59912] = {9'd91,10'd91};
ram[59913] = {9'd94,10'd94};
ram[59914] = {9'd97,10'd97};
ram[59915] = {-9'd100,10'd100};
ram[59916] = {-9'd97,10'd103};
ram[59917] = {-9'd94,10'd106};
ram[59918] = {-9'd91,10'd109};
ram[59919] = {-9'd88,10'd113};
ram[59920] = {-9'd85,10'd116};
ram[59921] = {-9'd81,10'd119};
ram[59922] = {-9'd78,10'd122};
ram[59923] = {-9'd75,10'd125};
ram[59924] = {-9'd72,10'd128};
ram[59925] = {-9'd69,10'd131};
ram[59926] = {-9'd66,10'd135};
ram[59927] = {-9'd63,10'd138};
ram[59928] = {-9'd59,10'd141};
ram[59929] = {-9'd56,10'd144};
ram[59930] = {-9'd53,10'd147};
ram[59931] = {-9'd50,10'd150};
ram[59932] = {-9'd47,10'd153};
ram[59933] = {-9'd44,10'd157};
ram[59934] = {-9'd41,10'd160};
ram[59935] = {-9'd37,10'd163};
ram[59936] = {-9'd34,10'd166};
ram[59937] = {-9'd31,10'd169};
ram[59938] = {-9'd28,10'd172};
ram[59939] = {-9'd25,10'd175};
ram[59940] = {-9'd22,10'd179};
ram[59941] = {-9'd19,10'd182};
ram[59942] = {-9'd15,10'd185};
ram[59943] = {-9'd12,10'd188};
ram[59944] = {-9'd9,10'd191};
ram[59945] = {-9'd6,10'd194};
ram[59946] = {-9'd3,10'd197};
ram[59947] = {9'd0,10'd201};
ram[59948] = {9'd3,10'd204};
ram[59949] = {9'd7,10'd207};
ram[59950] = {9'd10,10'd210};
ram[59951] = {9'd13,10'd213};
ram[59952] = {9'd16,10'd216};
ram[59953] = {9'd19,10'd219};
ram[59954] = {9'd22,10'd223};
ram[59955] = {9'd25,10'd226};
ram[59956] = {9'd29,10'd229};
ram[59957] = {9'd32,10'd232};
ram[59958] = {9'd35,10'd235};
ram[59959] = {9'd38,10'd238};
ram[59960] = {9'd41,10'd241};
ram[59961] = {9'd44,10'd245};
ram[59962] = {9'd47,10'd248};
ram[59963] = {9'd51,10'd251};
ram[59964] = {9'd54,10'd254};
ram[59965] = {9'd57,10'd257};
ram[59966] = {9'd60,10'd260};
ram[59967] = {9'd63,10'd263};
ram[59968] = {9'd66,10'd267};
ram[59969] = {9'd69,10'd270};
ram[59970] = {9'd73,10'd273};
ram[59971] = {9'd76,10'd276};
ram[59972] = {9'd79,10'd279};
ram[59973] = {9'd82,10'd282};
ram[59974] = {9'd85,10'd285};
ram[59975] = {9'd88,10'd289};
ram[59976] = {9'd91,10'd292};
ram[59977] = {9'd95,10'd295};
ram[59978] = {9'd98,10'd298};
ram[59979] = {-9'd99,10'd301};
ram[59980] = {-9'd96,10'd304};
ram[59981] = {-9'd93,10'd307};
ram[59982] = {-9'd90,10'd311};
ram[59983] = {-9'd87,10'd314};
ram[59984] = {-9'd84,10'd317};
ram[59985] = {-9'd81,10'd320};
ram[59986] = {-9'd77,10'd323};
ram[59987] = {-9'd74,10'd326};
ram[59988] = {-9'd71,10'd329};
ram[59989] = {-9'd68,10'd333};
ram[59990] = {-9'd65,10'd336};
ram[59991] = {-9'd62,10'd339};
ram[59992] = {-9'd59,10'd342};
ram[59993] = {-9'd55,10'd345};
ram[59994] = {-9'd52,10'd348};
ram[59995] = {-9'd49,10'd351};
ram[59996] = {-9'd46,10'd354};
ram[59997] = {-9'd43,10'd358};
ram[59998] = {-9'd40,10'd361};
ram[59999] = {-9'd37,10'd364};
ram[60000] = {-9'd33,10'd367};
ram[60001] = {-9'd30,10'd370};
ram[60002] = {-9'd27,10'd373};
ram[60003] = {-9'd24,10'd376};
ram[60004] = {-9'd21,10'd380};
ram[60005] = {-9'd18,10'd383};
ram[60006] = {-9'd15,10'd386};
ram[60007] = {-9'd11,10'd389};
ram[60008] = {-9'd8,10'd392};
ram[60009] = {-9'd5,10'd395};
ram[60010] = {-9'd2,10'd398};
ram[60011] = {9'd1,-10'd399};
ram[60012] = {9'd4,-10'd396};
ram[60013] = {9'd7,-10'd393};
ram[60014] = {9'd10,-10'd390};
ram[60015] = {9'd14,-10'd387};
ram[60016] = {9'd17,-10'd384};
ram[60017] = {9'd20,-10'd381};
ram[60018] = {9'd23,-10'd377};
ram[60019] = {9'd26,-10'd374};
ram[60020] = {9'd29,-10'd371};
ram[60021] = {9'd32,-10'd368};
ram[60022] = {9'd36,-10'd365};
ram[60023] = {9'd39,-10'd362};
ram[60024] = {9'd42,-10'd359};
ram[60025] = {9'd45,-10'd355};
ram[60026] = {9'd48,-10'd352};
ram[60027] = {9'd51,-10'd349};
ram[60028] = {9'd54,-10'd346};
ram[60029] = {9'd58,-10'd343};
ram[60030] = {9'd61,-10'd340};
ram[60031] = {9'd64,-10'd337};
ram[60032] = {9'd64,-10'd337};
ram[60033] = {9'd67,-10'd334};
ram[60034] = {9'd70,-10'd330};
ram[60035] = {9'd73,-10'd327};
ram[60036] = {9'd76,-10'd324};
ram[60037] = {9'd80,-10'd321};
ram[60038] = {9'd83,-10'd318};
ram[60039] = {9'd86,-10'd315};
ram[60040] = {9'd89,-10'd312};
ram[60041] = {9'd92,-10'd308};
ram[60042] = {9'd95,-10'd305};
ram[60043] = {9'd98,-10'd302};
ram[60044] = {-9'd99,-10'd299};
ram[60045] = {-9'd96,-10'd296};
ram[60046] = {-9'd92,-10'd293};
ram[60047] = {-9'd89,-10'd290};
ram[60048] = {-9'd86,-10'd286};
ram[60049] = {-9'd83,-10'd283};
ram[60050] = {-9'd80,-10'd280};
ram[60051] = {-9'd77,-10'd277};
ram[60052] = {-9'd74,-10'd274};
ram[60053] = {-9'd70,-10'd271};
ram[60054] = {-9'd67,-10'd268};
ram[60055] = {-9'd64,-10'd264};
ram[60056] = {-9'd61,-10'd261};
ram[60057] = {-9'd58,-10'd258};
ram[60058] = {-9'd55,-10'd255};
ram[60059] = {-9'd52,-10'd252};
ram[60060] = {-9'd48,-10'd249};
ram[60061] = {-9'd45,-10'd246};
ram[60062] = {-9'd42,-10'd242};
ram[60063] = {-9'd39,-10'd239};
ram[60064] = {-9'd36,-10'd236};
ram[60065] = {-9'd33,-10'd233};
ram[60066] = {-9'd30,-10'd230};
ram[60067] = {-9'd26,-10'd227};
ram[60068] = {-9'd23,-10'd224};
ram[60069] = {-9'd20,-10'd220};
ram[60070] = {-9'd17,-10'd217};
ram[60071] = {-9'd14,-10'd214};
ram[60072] = {-9'd11,-10'd211};
ram[60073] = {-9'd8,-10'd208};
ram[60074] = {-9'd4,-10'd205};
ram[60075] = {-9'd1,-10'd202};
ram[60076] = {9'd2,-10'd198};
ram[60077] = {9'd5,-10'd195};
ram[60078] = {9'd8,-10'd192};
ram[60079] = {9'd11,-10'd189};
ram[60080] = {9'd14,-10'd186};
ram[60081] = {9'd18,-10'd183};
ram[60082] = {9'd21,-10'd180};
ram[60083] = {9'd24,-10'd176};
ram[60084] = {9'd27,-10'd173};
ram[60085] = {9'd30,-10'd170};
ram[60086] = {9'd33,-10'd167};
ram[60087] = {9'd36,-10'd164};
ram[60088] = {9'd40,-10'd161};
ram[60089] = {9'd43,-10'd158};
ram[60090] = {9'd46,-10'd154};
ram[60091] = {9'd49,-10'd151};
ram[60092] = {9'd52,-10'd148};
ram[60093] = {9'd55,-10'd145};
ram[60094] = {9'd58,-10'd142};
ram[60095] = {9'd62,-10'd139};
ram[60096] = {9'd65,-10'd136};
ram[60097] = {9'd68,-10'd132};
ram[60098] = {9'd71,-10'd129};
ram[60099] = {9'd74,-10'd126};
ram[60100] = {9'd77,-10'd123};
ram[60101] = {9'd80,-10'd120};
ram[60102] = {9'd84,-10'd117};
ram[60103] = {9'd87,-10'd114};
ram[60104] = {9'd90,-10'd110};
ram[60105] = {9'd93,-10'd107};
ram[60106] = {9'd96,-10'd104};
ram[60107] = {9'd99,-10'd101};
ram[60108] = {-9'd98,-10'd98};
ram[60109] = {-9'd95,-10'd95};
ram[60110] = {-9'd92,-10'd92};
ram[60111] = {-9'd88,-10'd88};
ram[60112] = {-9'd85,-10'd85};
ram[60113] = {-9'd82,-10'd82};
ram[60114] = {-9'd79,-10'd79};
ram[60115] = {-9'd76,-10'd76};
ram[60116] = {-9'd73,-10'd73};
ram[60117] = {-9'd70,-10'd70};
ram[60118] = {-9'd66,-10'd66};
ram[60119] = {-9'd63,-10'd63};
ram[60120] = {-9'd60,-10'd60};
ram[60121] = {-9'd57,-10'd57};
ram[60122] = {-9'd54,-10'd54};
ram[60123] = {-9'd51,-10'd51};
ram[60124] = {-9'd48,-10'd48};
ram[60125] = {-9'd44,-10'd44};
ram[60126] = {-9'd41,-10'd41};
ram[60127] = {-9'd38,-10'd38};
ram[60128] = {-9'd35,-10'd35};
ram[60129] = {-9'd32,-10'd32};
ram[60130] = {-9'd29,-10'd29};
ram[60131] = {-9'd26,-10'd26};
ram[60132] = {-9'd22,-10'd22};
ram[60133] = {-9'd19,-10'd19};
ram[60134] = {-9'd16,-10'd16};
ram[60135] = {-9'd13,-10'd13};
ram[60136] = {-9'd10,-10'd10};
ram[60137] = {-9'd7,-10'd7};
ram[60138] = {-9'd4,-10'd4};
ram[60139] = {9'd0,10'd0};
ram[60140] = {9'd3,10'd3};
ram[60141] = {9'd6,10'd6};
ram[60142] = {9'd9,10'd9};
ram[60143] = {9'd12,10'd12};
ram[60144] = {9'd15,10'd15};
ram[60145] = {9'd18,10'd18};
ram[60146] = {9'd21,10'd21};
ram[60147] = {9'd25,10'd25};
ram[60148] = {9'd28,10'd28};
ram[60149] = {9'd31,10'd31};
ram[60150] = {9'd34,10'd34};
ram[60151] = {9'd37,10'd37};
ram[60152] = {9'd40,10'd40};
ram[60153] = {9'd43,10'd43};
ram[60154] = {9'd47,10'd47};
ram[60155] = {9'd50,10'd50};
ram[60156] = {9'd53,10'd53};
ram[60157] = {9'd56,10'd56};
ram[60158] = {9'd59,10'd59};
ram[60159] = {9'd62,10'd62};
ram[60160] = {9'd62,10'd62};
ram[60161] = {9'd65,10'd65};
ram[60162] = {9'd69,10'd69};
ram[60163] = {9'd72,10'd72};
ram[60164] = {9'd75,10'd75};
ram[60165] = {9'd78,10'd78};
ram[60166] = {9'd81,10'd81};
ram[60167] = {9'd84,10'd84};
ram[60168] = {9'd87,10'd87};
ram[60169] = {9'd91,10'd91};
ram[60170] = {9'd94,10'd94};
ram[60171] = {9'd97,10'd97};
ram[60172] = {-9'd100,10'd100};
ram[60173] = {-9'd97,10'd103};
ram[60174] = {-9'd94,10'd106};
ram[60175] = {-9'd91,10'd109};
ram[60176] = {-9'd88,10'd113};
ram[60177] = {-9'd85,10'd116};
ram[60178] = {-9'd81,10'd119};
ram[60179] = {-9'd78,10'd122};
ram[60180] = {-9'd75,10'd125};
ram[60181] = {-9'd72,10'd128};
ram[60182] = {-9'd69,10'd131};
ram[60183] = {-9'd66,10'd135};
ram[60184] = {-9'd63,10'd138};
ram[60185] = {-9'd59,10'd141};
ram[60186] = {-9'd56,10'd144};
ram[60187] = {-9'd53,10'd147};
ram[60188] = {-9'd50,10'd150};
ram[60189] = {-9'd47,10'd153};
ram[60190] = {-9'd44,10'd157};
ram[60191] = {-9'd41,10'd160};
ram[60192] = {-9'd37,10'd163};
ram[60193] = {-9'd34,10'd166};
ram[60194] = {-9'd31,10'd169};
ram[60195] = {-9'd28,10'd172};
ram[60196] = {-9'd25,10'd175};
ram[60197] = {-9'd22,10'd179};
ram[60198] = {-9'd19,10'd182};
ram[60199] = {-9'd15,10'd185};
ram[60200] = {-9'd12,10'd188};
ram[60201] = {-9'd9,10'd191};
ram[60202] = {-9'd6,10'd194};
ram[60203] = {-9'd3,10'd197};
ram[60204] = {9'd0,10'd201};
ram[60205] = {9'd3,10'd204};
ram[60206] = {9'd7,10'd207};
ram[60207] = {9'd10,10'd210};
ram[60208] = {9'd13,10'd213};
ram[60209] = {9'd16,10'd216};
ram[60210] = {9'd19,10'd219};
ram[60211] = {9'd22,10'd223};
ram[60212] = {9'd25,10'd226};
ram[60213] = {9'd29,10'd229};
ram[60214] = {9'd32,10'd232};
ram[60215] = {9'd35,10'd235};
ram[60216] = {9'd38,10'd238};
ram[60217] = {9'd41,10'd241};
ram[60218] = {9'd44,10'd245};
ram[60219] = {9'd47,10'd248};
ram[60220] = {9'd51,10'd251};
ram[60221] = {9'd54,10'd254};
ram[60222] = {9'd57,10'd257};
ram[60223] = {9'd60,10'd260};
ram[60224] = {9'd63,10'd263};
ram[60225] = {9'd66,10'd267};
ram[60226] = {9'd69,10'd270};
ram[60227] = {9'd73,10'd273};
ram[60228] = {9'd76,10'd276};
ram[60229] = {9'd79,10'd279};
ram[60230] = {9'd82,10'd282};
ram[60231] = {9'd85,10'd285};
ram[60232] = {9'd88,10'd289};
ram[60233] = {9'd91,10'd292};
ram[60234] = {9'd95,10'd295};
ram[60235] = {9'd98,10'd298};
ram[60236] = {-9'd99,10'd301};
ram[60237] = {-9'd96,10'd304};
ram[60238] = {-9'd93,10'd307};
ram[60239] = {-9'd90,10'd311};
ram[60240] = {-9'd87,10'd314};
ram[60241] = {-9'd84,10'd317};
ram[60242] = {-9'd81,10'd320};
ram[60243] = {-9'd77,10'd323};
ram[60244] = {-9'd74,10'd326};
ram[60245] = {-9'd71,10'd329};
ram[60246] = {-9'd68,10'd333};
ram[60247] = {-9'd65,10'd336};
ram[60248] = {-9'd62,10'd339};
ram[60249] = {-9'd59,10'd342};
ram[60250] = {-9'd55,10'd345};
ram[60251] = {-9'd52,10'd348};
ram[60252] = {-9'd49,10'd351};
ram[60253] = {-9'd46,10'd354};
ram[60254] = {-9'd43,10'd358};
ram[60255] = {-9'd40,10'd361};
ram[60256] = {-9'd37,10'd364};
ram[60257] = {-9'd33,10'd367};
ram[60258] = {-9'd30,10'd370};
ram[60259] = {-9'd27,10'd373};
ram[60260] = {-9'd24,10'd376};
ram[60261] = {-9'd21,10'd380};
ram[60262] = {-9'd18,10'd383};
ram[60263] = {-9'd15,10'd386};
ram[60264] = {-9'd11,10'd389};
ram[60265] = {-9'd8,10'd392};
ram[60266] = {-9'd5,10'd395};
ram[60267] = {-9'd2,10'd398};
ram[60268] = {9'd1,-10'd399};
ram[60269] = {9'd4,-10'd396};
ram[60270] = {9'd7,-10'd393};
ram[60271] = {9'd10,-10'd390};
ram[60272] = {9'd14,-10'd387};
ram[60273] = {9'd17,-10'd384};
ram[60274] = {9'd20,-10'd381};
ram[60275] = {9'd23,-10'd377};
ram[60276] = {9'd26,-10'd374};
ram[60277] = {9'd29,-10'd371};
ram[60278] = {9'd32,-10'd368};
ram[60279] = {9'd36,-10'd365};
ram[60280] = {9'd39,-10'd362};
ram[60281] = {9'd42,-10'd359};
ram[60282] = {9'd45,-10'd355};
ram[60283] = {9'd48,-10'd352};
ram[60284] = {9'd51,-10'd349};
ram[60285] = {9'd54,-10'd346};
ram[60286] = {9'd58,-10'd343};
ram[60287] = {9'd61,-10'd340};
ram[60288] = {9'd61,-10'd340};
ram[60289] = {9'd64,-10'd337};
ram[60290] = {9'd67,-10'd334};
ram[60291] = {9'd70,-10'd330};
ram[60292] = {9'd73,-10'd327};
ram[60293] = {9'd76,-10'd324};
ram[60294] = {9'd80,-10'd321};
ram[60295] = {9'd83,-10'd318};
ram[60296] = {9'd86,-10'd315};
ram[60297] = {9'd89,-10'd312};
ram[60298] = {9'd92,-10'd308};
ram[60299] = {9'd95,-10'd305};
ram[60300] = {9'd98,-10'd302};
ram[60301] = {-9'd99,-10'd299};
ram[60302] = {-9'd96,-10'd296};
ram[60303] = {-9'd92,-10'd293};
ram[60304] = {-9'd89,-10'd290};
ram[60305] = {-9'd86,-10'd286};
ram[60306] = {-9'd83,-10'd283};
ram[60307] = {-9'd80,-10'd280};
ram[60308] = {-9'd77,-10'd277};
ram[60309] = {-9'd74,-10'd274};
ram[60310] = {-9'd70,-10'd271};
ram[60311] = {-9'd67,-10'd268};
ram[60312] = {-9'd64,-10'd264};
ram[60313] = {-9'd61,-10'd261};
ram[60314] = {-9'd58,-10'd258};
ram[60315] = {-9'd55,-10'd255};
ram[60316] = {-9'd52,-10'd252};
ram[60317] = {-9'd48,-10'd249};
ram[60318] = {-9'd45,-10'd246};
ram[60319] = {-9'd42,-10'd242};
ram[60320] = {-9'd39,-10'd239};
ram[60321] = {-9'd36,-10'd236};
ram[60322] = {-9'd33,-10'd233};
ram[60323] = {-9'd30,-10'd230};
ram[60324] = {-9'd26,-10'd227};
ram[60325] = {-9'd23,-10'd224};
ram[60326] = {-9'd20,-10'd220};
ram[60327] = {-9'd17,-10'd217};
ram[60328] = {-9'd14,-10'd214};
ram[60329] = {-9'd11,-10'd211};
ram[60330] = {-9'd8,-10'd208};
ram[60331] = {-9'd4,-10'd205};
ram[60332] = {-9'd1,-10'd202};
ram[60333] = {9'd2,-10'd198};
ram[60334] = {9'd5,-10'd195};
ram[60335] = {9'd8,-10'd192};
ram[60336] = {9'd11,-10'd189};
ram[60337] = {9'd14,-10'd186};
ram[60338] = {9'd18,-10'd183};
ram[60339] = {9'd21,-10'd180};
ram[60340] = {9'd24,-10'd176};
ram[60341] = {9'd27,-10'd173};
ram[60342] = {9'd30,-10'd170};
ram[60343] = {9'd33,-10'd167};
ram[60344] = {9'd36,-10'd164};
ram[60345] = {9'd40,-10'd161};
ram[60346] = {9'd43,-10'd158};
ram[60347] = {9'd46,-10'd154};
ram[60348] = {9'd49,-10'd151};
ram[60349] = {9'd52,-10'd148};
ram[60350] = {9'd55,-10'd145};
ram[60351] = {9'd58,-10'd142};
ram[60352] = {9'd62,-10'd139};
ram[60353] = {9'd65,-10'd136};
ram[60354] = {9'd68,-10'd132};
ram[60355] = {9'd71,-10'd129};
ram[60356] = {9'd74,-10'd126};
ram[60357] = {9'd77,-10'd123};
ram[60358] = {9'd80,-10'd120};
ram[60359] = {9'd84,-10'd117};
ram[60360] = {9'd87,-10'd114};
ram[60361] = {9'd90,-10'd110};
ram[60362] = {9'd93,-10'd107};
ram[60363] = {9'd96,-10'd104};
ram[60364] = {9'd99,-10'd101};
ram[60365] = {-9'd98,-10'd98};
ram[60366] = {-9'd95,-10'd95};
ram[60367] = {-9'd92,-10'd92};
ram[60368] = {-9'd88,-10'd88};
ram[60369] = {-9'd85,-10'd85};
ram[60370] = {-9'd82,-10'd82};
ram[60371] = {-9'd79,-10'd79};
ram[60372] = {-9'd76,-10'd76};
ram[60373] = {-9'd73,-10'd73};
ram[60374] = {-9'd70,-10'd70};
ram[60375] = {-9'd66,-10'd66};
ram[60376] = {-9'd63,-10'd63};
ram[60377] = {-9'd60,-10'd60};
ram[60378] = {-9'd57,-10'd57};
ram[60379] = {-9'd54,-10'd54};
ram[60380] = {-9'd51,-10'd51};
ram[60381] = {-9'd48,-10'd48};
ram[60382] = {-9'd44,-10'd44};
ram[60383] = {-9'd41,-10'd41};
ram[60384] = {-9'd38,-10'd38};
ram[60385] = {-9'd35,-10'd35};
ram[60386] = {-9'd32,-10'd32};
ram[60387] = {-9'd29,-10'd29};
ram[60388] = {-9'd26,-10'd26};
ram[60389] = {-9'd22,-10'd22};
ram[60390] = {-9'd19,-10'd19};
ram[60391] = {-9'd16,-10'd16};
ram[60392] = {-9'd13,-10'd13};
ram[60393] = {-9'd10,-10'd10};
ram[60394] = {-9'd7,-10'd7};
ram[60395] = {-9'd4,-10'd4};
ram[60396] = {9'd0,10'd0};
ram[60397] = {9'd3,10'd3};
ram[60398] = {9'd6,10'd6};
ram[60399] = {9'd9,10'd9};
ram[60400] = {9'd12,10'd12};
ram[60401] = {9'd15,10'd15};
ram[60402] = {9'd18,10'd18};
ram[60403] = {9'd21,10'd21};
ram[60404] = {9'd25,10'd25};
ram[60405] = {9'd28,10'd28};
ram[60406] = {9'd31,10'd31};
ram[60407] = {9'd34,10'd34};
ram[60408] = {9'd37,10'd37};
ram[60409] = {9'd40,10'd40};
ram[60410] = {9'd43,10'd43};
ram[60411] = {9'd47,10'd47};
ram[60412] = {9'd50,10'd50};
ram[60413] = {9'd53,10'd53};
ram[60414] = {9'd56,10'd56};
ram[60415] = {9'd59,10'd59};
ram[60416] = {9'd59,10'd59};
ram[60417] = {9'd62,10'd62};
ram[60418] = {9'd65,10'd65};
ram[60419] = {9'd69,10'd69};
ram[60420] = {9'd72,10'd72};
ram[60421] = {9'd75,10'd75};
ram[60422] = {9'd78,10'd78};
ram[60423] = {9'd81,10'd81};
ram[60424] = {9'd84,10'd84};
ram[60425] = {9'd87,10'd87};
ram[60426] = {9'd91,10'd91};
ram[60427] = {9'd94,10'd94};
ram[60428] = {9'd97,10'd97};
ram[60429] = {-9'd100,10'd100};
ram[60430] = {-9'd97,10'd103};
ram[60431] = {-9'd94,10'd106};
ram[60432] = {-9'd91,10'd109};
ram[60433] = {-9'd88,10'd113};
ram[60434] = {-9'd85,10'd116};
ram[60435] = {-9'd81,10'd119};
ram[60436] = {-9'd78,10'd122};
ram[60437] = {-9'd75,10'd125};
ram[60438] = {-9'd72,10'd128};
ram[60439] = {-9'd69,10'd131};
ram[60440] = {-9'd66,10'd135};
ram[60441] = {-9'd63,10'd138};
ram[60442] = {-9'd59,10'd141};
ram[60443] = {-9'd56,10'd144};
ram[60444] = {-9'd53,10'd147};
ram[60445] = {-9'd50,10'd150};
ram[60446] = {-9'd47,10'd153};
ram[60447] = {-9'd44,10'd157};
ram[60448] = {-9'd41,10'd160};
ram[60449] = {-9'd37,10'd163};
ram[60450] = {-9'd34,10'd166};
ram[60451] = {-9'd31,10'd169};
ram[60452] = {-9'd28,10'd172};
ram[60453] = {-9'd25,10'd175};
ram[60454] = {-9'd22,10'd179};
ram[60455] = {-9'd19,10'd182};
ram[60456] = {-9'd15,10'd185};
ram[60457] = {-9'd12,10'd188};
ram[60458] = {-9'd9,10'd191};
ram[60459] = {-9'd6,10'd194};
ram[60460] = {-9'd3,10'd197};
ram[60461] = {9'd0,10'd201};
ram[60462] = {9'd3,10'd204};
ram[60463] = {9'd7,10'd207};
ram[60464] = {9'd10,10'd210};
ram[60465] = {9'd13,10'd213};
ram[60466] = {9'd16,10'd216};
ram[60467] = {9'd19,10'd219};
ram[60468] = {9'd22,10'd223};
ram[60469] = {9'd25,10'd226};
ram[60470] = {9'd29,10'd229};
ram[60471] = {9'd32,10'd232};
ram[60472] = {9'd35,10'd235};
ram[60473] = {9'd38,10'd238};
ram[60474] = {9'd41,10'd241};
ram[60475] = {9'd44,10'd245};
ram[60476] = {9'd47,10'd248};
ram[60477] = {9'd51,10'd251};
ram[60478] = {9'd54,10'd254};
ram[60479] = {9'd57,10'd257};
ram[60480] = {9'd60,10'd260};
ram[60481] = {9'd63,10'd263};
ram[60482] = {9'd66,10'd267};
ram[60483] = {9'd69,10'd270};
ram[60484] = {9'd73,10'd273};
ram[60485] = {9'd76,10'd276};
ram[60486] = {9'd79,10'd279};
ram[60487] = {9'd82,10'd282};
ram[60488] = {9'd85,10'd285};
ram[60489] = {9'd88,10'd289};
ram[60490] = {9'd91,10'd292};
ram[60491] = {9'd95,10'd295};
ram[60492] = {9'd98,10'd298};
ram[60493] = {-9'd99,10'd301};
ram[60494] = {-9'd96,10'd304};
ram[60495] = {-9'd93,10'd307};
ram[60496] = {-9'd90,10'd311};
ram[60497] = {-9'd87,10'd314};
ram[60498] = {-9'd84,10'd317};
ram[60499] = {-9'd81,10'd320};
ram[60500] = {-9'd77,10'd323};
ram[60501] = {-9'd74,10'd326};
ram[60502] = {-9'd71,10'd329};
ram[60503] = {-9'd68,10'd333};
ram[60504] = {-9'd65,10'd336};
ram[60505] = {-9'd62,10'd339};
ram[60506] = {-9'd59,10'd342};
ram[60507] = {-9'd55,10'd345};
ram[60508] = {-9'd52,10'd348};
ram[60509] = {-9'd49,10'd351};
ram[60510] = {-9'd46,10'd354};
ram[60511] = {-9'd43,10'd358};
ram[60512] = {-9'd40,10'd361};
ram[60513] = {-9'd37,10'd364};
ram[60514] = {-9'd33,10'd367};
ram[60515] = {-9'd30,10'd370};
ram[60516] = {-9'd27,10'd373};
ram[60517] = {-9'd24,10'd376};
ram[60518] = {-9'd21,10'd380};
ram[60519] = {-9'd18,10'd383};
ram[60520] = {-9'd15,10'd386};
ram[60521] = {-9'd11,10'd389};
ram[60522] = {-9'd8,10'd392};
ram[60523] = {-9'd5,10'd395};
ram[60524] = {-9'd2,10'd398};
ram[60525] = {9'd1,-10'd399};
ram[60526] = {9'd4,-10'd396};
ram[60527] = {9'd7,-10'd393};
ram[60528] = {9'd10,-10'd390};
ram[60529] = {9'd14,-10'd387};
ram[60530] = {9'd17,-10'd384};
ram[60531] = {9'd20,-10'd381};
ram[60532] = {9'd23,-10'd377};
ram[60533] = {9'd26,-10'd374};
ram[60534] = {9'd29,-10'd371};
ram[60535] = {9'd32,-10'd368};
ram[60536] = {9'd36,-10'd365};
ram[60537] = {9'd39,-10'd362};
ram[60538] = {9'd42,-10'd359};
ram[60539] = {9'd45,-10'd355};
ram[60540] = {9'd48,-10'd352};
ram[60541] = {9'd51,-10'd349};
ram[60542] = {9'd54,-10'd346};
ram[60543] = {9'd58,-10'd343};
ram[60544] = {9'd58,-10'd343};
ram[60545] = {9'd61,-10'd340};
ram[60546] = {9'd64,-10'd337};
ram[60547] = {9'd67,-10'd334};
ram[60548] = {9'd70,-10'd330};
ram[60549] = {9'd73,-10'd327};
ram[60550] = {9'd76,-10'd324};
ram[60551] = {9'd80,-10'd321};
ram[60552] = {9'd83,-10'd318};
ram[60553] = {9'd86,-10'd315};
ram[60554] = {9'd89,-10'd312};
ram[60555] = {9'd92,-10'd308};
ram[60556] = {9'd95,-10'd305};
ram[60557] = {9'd98,-10'd302};
ram[60558] = {-9'd99,-10'd299};
ram[60559] = {-9'd96,-10'd296};
ram[60560] = {-9'd92,-10'd293};
ram[60561] = {-9'd89,-10'd290};
ram[60562] = {-9'd86,-10'd286};
ram[60563] = {-9'd83,-10'd283};
ram[60564] = {-9'd80,-10'd280};
ram[60565] = {-9'd77,-10'd277};
ram[60566] = {-9'd74,-10'd274};
ram[60567] = {-9'd70,-10'd271};
ram[60568] = {-9'd67,-10'd268};
ram[60569] = {-9'd64,-10'd264};
ram[60570] = {-9'd61,-10'd261};
ram[60571] = {-9'd58,-10'd258};
ram[60572] = {-9'd55,-10'd255};
ram[60573] = {-9'd52,-10'd252};
ram[60574] = {-9'd48,-10'd249};
ram[60575] = {-9'd45,-10'd246};
ram[60576] = {-9'd42,-10'd242};
ram[60577] = {-9'd39,-10'd239};
ram[60578] = {-9'd36,-10'd236};
ram[60579] = {-9'd33,-10'd233};
ram[60580] = {-9'd30,-10'd230};
ram[60581] = {-9'd26,-10'd227};
ram[60582] = {-9'd23,-10'd224};
ram[60583] = {-9'd20,-10'd220};
ram[60584] = {-9'd17,-10'd217};
ram[60585] = {-9'd14,-10'd214};
ram[60586] = {-9'd11,-10'd211};
ram[60587] = {-9'd8,-10'd208};
ram[60588] = {-9'd4,-10'd205};
ram[60589] = {-9'd1,-10'd202};
ram[60590] = {9'd2,-10'd198};
ram[60591] = {9'd5,-10'd195};
ram[60592] = {9'd8,-10'd192};
ram[60593] = {9'd11,-10'd189};
ram[60594] = {9'd14,-10'd186};
ram[60595] = {9'd18,-10'd183};
ram[60596] = {9'd21,-10'd180};
ram[60597] = {9'd24,-10'd176};
ram[60598] = {9'd27,-10'd173};
ram[60599] = {9'd30,-10'd170};
ram[60600] = {9'd33,-10'd167};
ram[60601] = {9'd36,-10'd164};
ram[60602] = {9'd40,-10'd161};
ram[60603] = {9'd43,-10'd158};
ram[60604] = {9'd46,-10'd154};
ram[60605] = {9'd49,-10'd151};
ram[60606] = {9'd52,-10'd148};
ram[60607] = {9'd55,-10'd145};
ram[60608] = {9'd58,-10'd142};
ram[60609] = {9'd62,-10'd139};
ram[60610] = {9'd65,-10'd136};
ram[60611] = {9'd68,-10'd132};
ram[60612] = {9'd71,-10'd129};
ram[60613] = {9'd74,-10'd126};
ram[60614] = {9'd77,-10'd123};
ram[60615] = {9'd80,-10'd120};
ram[60616] = {9'd84,-10'd117};
ram[60617] = {9'd87,-10'd114};
ram[60618] = {9'd90,-10'd110};
ram[60619] = {9'd93,-10'd107};
ram[60620] = {9'd96,-10'd104};
ram[60621] = {9'd99,-10'd101};
ram[60622] = {-9'd98,-10'd98};
ram[60623] = {-9'd95,-10'd95};
ram[60624] = {-9'd92,-10'd92};
ram[60625] = {-9'd88,-10'd88};
ram[60626] = {-9'd85,-10'd85};
ram[60627] = {-9'd82,-10'd82};
ram[60628] = {-9'd79,-10'd79};
ram[60629] = {-9'd76,-10'd76};
ram[60630] = {-9'd73,-10'd73};
ram[60631] = {-9'd70,-10'd70};
ram[60632] = {-9'd66,-10'd66};
ram[60633] = {-9'd63,-10'd63};
ram[60634] = {-9'd60,-10'd60};
ram[60635] = {-9'd57,-10'd57};
ram[60636] = {-9'd54,-10'd54};
ram[60637] = {-9'd51,-10'd51};
ram[60638] = {-9'd48,-10'd48};
ram[60639] = {-9'd44,-10'd44};
ram[60640] = {-9'd41,-10'd41};
ram[60641] = {-9'd38,-10'd38};
ram[60642] = {-9'd35,-10'd35};
ram[60643] = {-9'd32,-10'd32};
ram[60644] = {-9'd29,-10'd29};
ram[60645] = {-9'd26,-10'd26};
ram[60646] = {-9'd22,-10'd22};
ram[60647] = {-9'd19,-10'd19};
ram[60648] = {-9'd16,-10'd16};
ram[60649] = {-9'd13,-10'd13};
ram[60650] = {-9'd10,-10'd10};
ram[60651] = {-9'd7,-10'd7};
ram[60652] = {-9'd4,-10'd4};
ram[60653] = {9'd0,10'd0};
ram[60654] = {9'd3,10'd3};
ram[60655] = {9'd6,10'd6};
ram[60656] = {9'd9,10'd9};
ram[60657] = {9'd12,10'd12};
ram[60658] = {9'd15,10'd15};
ram[60659] = {9'd18,10'd18};
ram[60660] = {9'd21,10'd21};
ram[60661] = {9'd25,10'd25};
ram[60662] = {9'd28,10'd28};
ram[60663] = {9'd31,10'd31};
ram[60664] = {9'd34,10'd34};
ram[60665] = {9'd37,10'd37};
ram[60666] = {9'd40,10'd40};
ram[60667] = {9'd43,10'd43};
ram[60668] = {9'd47,10'd47};
ram[60669] = {9'd50,10'd50};
ram[60670] = {9'd53,10'd53};
ram[60671] = {9'd56,10'd56};
ram[60672] = {9'd56,10'd56};
ram[60673] = {9'd59,10'd59};
ram[60674] = {9'd62,10'd62};
ram[60675] = {9'd65,10'd65};
ram[60676] = {9'd69,10'd69};
ram[60677] = {9'd72,10'd72};
ram[60678] = {9'd75,10'd75};
ram[60679] = {9'd78,10'd78};
ram[60680] = {9'd81,10'd81};
ram[60681] = {9'd84,10'd84};
ram[60682] = {9'd87,10'd87};
ram[60683] = {9'd91,10'd91};
ram[60684] = {9'd94,10'd94};
ram[60685] = {9'd97,10'd97};
ram[60686] = {-9'd100,10'd100};
ram[60687] = {-9'd97,10'd103};
ram[60688] = {-9'd94,10'd106};
ram[60689] = {-9'd91,10'd109};
ram[60690] = {-9'd88,10'd113};
ram[60691] = {-9'd85,10'd116};
ram[60692] = {-9'd81,10'd119};
ram[60693] = {-9'd78,10'd122};
ram[60694] = {-9'd75,10'd125};
ram[60695] = {-9'd72,10'd128};
ram[60696] = {-9'd69,10'd131};
ram[60697] = {-9'd66,10'd135};
ram[60698] = {-9'd63,10'd138};
ram[60699] = {-9'd59,10'd141};
ram[60700] = {-9'd56,10'd144};
ram[60701] = {-9'd53,10'd147};
ram[60702] = {-9'd50,10'd150};
ram[60703] = {-9'd47,10'd153};
ram[60704] = {-9'd44,10'd157};
ram[60705] = {-9'd41,10'd160};
ram[60706] = {-9'd37,10'd163};
ram[60707] = {-9'd34,10'd166};
ram[60708] = {-9'd31,10'd169};
ram[60709] = {-9'd28,10'd172};
ram[60710] = {-9'd25,10'd175};
ram[60711] = {-9'd22,10'd179};
ram[60712] = {-9'd19,10'd182};
ram[60713] = {-9'd15,10'd185};
ram[60714] = {-9'd12,10'd188};
ram[60715] = {-9'd9,10'd191};
ram[60716] = {-9'd6,10'd194};
ram[60717] = {-9'd3,10'd197};
ram[60718] = {9'd0,10'd201};
ram[60719] = {9'd3,10'd204};
ram[60720] = {9'd7,10'd207};
ram[60721] = {9'd10,10'd210};
ram[60722] = {9'd13,10'd213};
ram[60723] = {9'd16,10'd216};
ram[60724] = {9'd19,10'd219};
ram[60725] = {9'd22,10'd223};
ram[60726] = {9'd25,10'd226};
ram[60727] = {9'd29,10'd229};
ram[60728] = {9'd32,10'd232};
ram[60729] = {9'd35,10'd235};
ram[60730] = {9'd38,10'd238};
ram[60731] = {9'd41,10'd241};
ram[60732] = {9'd44,10'd245};
ram[60733] = {9'd47,10'd248};
ram[60734] = {9'd51,10'd251};
ram[60735] = {9'd54,10'd254};
ram[60736] = {9'd57,10'd257};
ram[60737] = {9'd60,10'd260};
ram[60738] = {9'd63,10'd263};
ram[60739] = {9'd66,10'd267};
ram[60740] = {9'd69,10'd270};
ram[60741] = {9'd73,10'd273};
ram[60742] = {9'd76,10'd276};
ram[60743] = {9'd79,10'd279};
ram[60744] = {9'd82,10'd282};
ram[60745] = {9'd85,10'd285};
ram[60746] = {9'd88,10'd289};
ram[60747] = {9'd91,10'd292};
ram[60748] = {9'd95,10'd295};
ram[60749] = {9'd98,10'd298};
ram[60750] = {-9'd99,10'd301};
ram[60751] = {-9'd96,10'd304};
ram[60752] = {-9'd93,10'd307};
ram[60753] = {-9'd90,10'd311};
ram[60754] = {-9'd87,10'd314};
ram[60755] = {-9'd84,10'd317};
ram[60756] = {-9'd81,10'd320};
ram[60757] = {-9'd77,10'd323};
ram[60758] = {-9'd74,10'd326};
ram[60759] = {-9'd71,10'd329};
ram[60760] = {-9'd68,10'd333};
ram[60761] = {-9'd65,10'd336};
ram[60762] = {-9'd62,10'd339};
ram[60763] = {-9'd59,10'd342};
ram[60764] = {-9'd55,10'd345};
ram[60765] = {-9'd52,10'd348};
ram[60766] = {-9'd49,10'd351};
ram[60767] = {-9'd46,10'd354};
ram[60768] = {-9'd43,10'd358};
ram[60769] = {-9'd40,10'd361};
ram[60770] = {-9'd37,10'd364};
ram[60771] = {-9'd33,10'd367};
ram[60772] = {-9'd30,10'd370};
ram[60773] = {-9'd27,10'd373};
ram[60774] = {-9'd24,10'd376};
ram[60775] = {-9'd21,10'd380};
ram[60776] = {-9'd18,10'd383};
ram[60777] = {-9'd15,10'd386};
ram[60778] = {-9'd11,10'd389};
ram[60779] = {-9'd8,10'd392};
ram[60780] = {-9'd5,10'd395};
ram[60781] = {-9'd2,10'd398};
ram[60782] = {9'd1,-10'd399};
ram[60783] = {9'd4,-10'd396};
ram[60784] = {9'd7,-10'd393};
ram[60785] = {9'd10,-10'd390};
ram[60786] = {9'd14,-10'd387};
ram[60787] = {9'd17,-10'd384};
ram[60788] = {9'd20,-10'd381};
ram[60789] = {9'd23,-10'd377};
ram[60790] = {9'd26,-10'd374};
ram[60791] = {9'd29,-10'd371};
ram[60792] = {9'd32,-10'd368};
ram[60793] = {9'd36,-10'd365};
ram[60794] = {9'd39,-10'd362};
ram[60795] = {9'd42,-10'd359};
ram[60796] = {9'd45,-10'd355};
ram[60797] = {9'd48,-10'd352};
ram[60798] = {9'd51,-10'd349};
ram[60799] = {9'd54,-10'd346};
ram[60800] = {9'd54,-10'd346};
ram[60801] = {9'd58,-10'd343};
ram[60802] = {9'd61,-10'd340};
ram[60803] = {9'd64,-10'd337};
ram[60804] = {9'd67,-10'd334};
ram[60805] = {9'd70,-10'd330};
ram[60806] = {9'd73,-10'd327};
ram[60807] = {9'd76,-10'd324};
ram[60808] = {9'd80,-10'd321};
ram[60809] = {9'd83,-10'd318};
ram[60810] = {9'd86,-10'd315};
ram[60811] = {9'd89,-10'd312};
ram[60812] = {9'd92,-10'd308};
ram[60813] = {9'd95,-10'd305};
ram[60814] = {9'd98,-10'd302};
ram[60815] = {-9'd99,-10'd299};
ram[60816] = {-9'd96,-10'd296};
ram[60817] = {-9'd92,-10'd293};
ram[60818] = {-9'd89,-10'd290};
ram[60819] = {-9'd86,-10'd286};
ram[60820] = {-9'd83,-10'd283};
ram[60821] = {-9'd80,-10'd280};
ram[60822] = {-9'd77,-10'd277};
ram[60823] = {-9'd74,-10'd274};
ram[60824] = {-9'd70,-10'd271};
ram[60825] = {-9'd67,-10'd268};
ram[60826] = {-9'd64,-10'd264};
ram[60827] = {-9'd61,-10'd261};
ram[60828] = {-9'd58,-10'd258};
ram[60829] = {-9'd55,-10'd255};
ram[60830] = {-9'd52,-10'd252};
ram[60831] = {-9'd48,-10'd249};
ram[60832] = {-9'd45,-10'd246};
ram[60833] = {-9'd42,-10'd242};
ram[60834] = {-9'd39,-10'd239};
ram[60835] = {-9'd36,-10'd236};
ram[60836] = {-9'd33,-10'd233};
ram[60837] = {-9'd30,-10'd230};
ram[60838] = {-9'd26,-10'd227};
ram[60839] = {-9'd23,-10'd224};
ram[60840] = {-9'd20,-10'd220};
ram[60841] = {-9'd17,-10'd217};
ram[60842] = {-9'd14,-10'd214};
ram[60843] = {-9'd11,-10'd211};
ram[60844] = {-9'd8,-10'd208};
ram[60845] = {-9'd4,-10'd205};
ram[60846] = {-9'd1,-10'd202};
ram[60847] = {9'd2,-10'd198};
ram[60848] = {9'd5,-10'd195};
ram[60849] = {9'd8,-10'd192};
ram[60850] = {9'd11,-10'd189};
ram[60851] = {9'd14,-10'd186};
ram[60852] = {9'd18,-10'd183};
ram[60853] = {9'd21,-10'd180};
ram[60854] = {9'd24,-10'd176};
ram[60855] = {9'd27,-10'd173};
ram[60856] = {9'd30,-10'd170};
ram[60857] = {9'd33,-10'd167};
ram[60858] = {9'd36,-10'd164};
ram[60859] = {9'd40,-10'd161};
ram[60860] = {9'd43,-10'd158};
ram[60861] = {9'd46,-10'd154};
ram[60862] = {9'd49,-10'd151};
ram[60863] = {9'd52,-10'd148};
ram[60864] = {9'd55,-10'd145};
ram[60865] = {9'd58,-10'd142};
ram[60866] = {9'd62,-10'd139};
ram[60867] = {9'd65,-10'd136};
ram[60868] = {9'd68,-10'd132};
ram[60869] = {9'd71,-10'd129};
ram[60870] = {9'd74,-10'd126};
ram[60871] = {9'd77,-10'd123};
ram[60872] = {9'd80,-10'd120};
ram[60873] = {9'd84,-10'd117};
ram[60874] = {9'd87,-10'd114};
ram[60875] = {9'd90,-10'd110};
ram[60876] = {9'd93,-10'd107};
ram[60877] = {9'd96,-10'd104};
ram[60878] = {9'd99,-10'd101};
ram[60879] = {-9'd98,-10'd98};
ram[60880] = {-9'd95,-10'd95};
ram[60881] = {-9'd92,-10'd92};
ram[60882] = {-9'd88,-10'd88};
ram[60883] = {-9'd85,-10'd85};
ram[60884] = {-9'd82,-10'd82};
ram[60885] = {-9'd79,-10'd79};
ram[60886] = {-9'd76,-10'd76};
ram[60887] = {-9'd73,-10'd73};
ram[60888] = {-9'd70,-10'd70};
ram[60889] = {-9'd66,-10'd66};
ram[60890] = {-9'd63,-10'd63};
ram[60891] = {-9'd60,-10'd60};
ram[60892] = {-9'd57,-10'd57};
ram[60893] = {-9'd54,-10'd54};
ram[60894] = {-9'd51,-10'd51};
ram[60895] = {-9'd48,-10'd48};
ram[60896] = {-9'd44,-10'd44};
ram[60897] = {-9'd41,-10'd41};
ram[60898] = {-9'd38,-10'd38};
ram[60899] = {-9'd35,-10'd35};
ram[60900] = {-9'd32,-10'd32};
ram[60901] = {-9'd29,-10'd29};
ram[60902] = {-9'd26,-10'd26};
ram[60903] = {-9'd22,-10'd22};
ram[60904] = {-9'd19,-10'd19};
ram[60905] = {-9'd16,-10'd16};
ram[60906] = {-9'd13,-10'd13};
ram[60907] = {-9'd10,-10'd10};
ram[60908] = {-9'd7,-10'd7};
ram[60909] = {-9'd4,-10'd4};
ram[60910] = {9'd0,10'd0};
ram[60911] = {9'd3,10'd3};
ram[60912] = {9'd6,10'd6};
ram[60913] = {9'd9,10'd9};
ram[60914] = {9'd12,10'd12};
ram[60915] = {9'd15,10'd15};
ram[60916] = {9'd18,10'd18};
ram[60917] = {9'd21,10'd21};
ram[60918] = {9'd25,10'd25};
ram[60919] = {9'd28,10'd28};
ram[60920] = {9'd31,10'd31};
ram[60921] = {9'd34,10'd34};
ram[60922] = {9'd37,10'd37};
ram[60923] = {9'd40,10'd40};
ram[60924] = {9'd43,10'd43};
ram[60925] = {9'd47,10'd47};
ram[60926] = {9'd50,10'd50};
ram[60927] = {9'd53,10'd53};
ram[60928] = {9'd53,10'd53};
ram[60929] = {9'd56,10'd56};
ram[60930] = {9'd59,10'd59};
ram[60931] = {9'd62,10'd62};
ram[60932] = {9'd65,10'd65};
ram[60933] = {9'd69,10'd69};
ram[60934] = {9'd72,10'd72};
ram[60935] = {9'd75,10'd75};
ram[60936] = {9'd78,10'd78};
ram[60937] = {9'd81,10'd81};
ram[60938] = {9'd84,10'd84};
ram[60939] = {9'd87,10'd87};
ram[60940] = {9'd91,10'd91};
ram[60941] = {9'd94,10'd94};
ram[60942] = {9'd97,10'd97};
ram[60943] = {-9'd100,10'd100};
ram[60944] = {-9'd97,10'd103};
ram[60945] = {-9'd94,10'd106};
ram[60946] = {-9'd91,10'd109};
ram[60947] = {-9'd88,10'd113};
ram[60948] = {-9'd85,10'd116};
ram[60949] = {-9'd81,10'd119};
ram[60950] = {-9'd78,10'd122};
ram[60951] = {-9'd75,10'd125};
ram[60952] = {-9'd72,10'd128};
ram[60953] = {-9'd69,10'd131};
ram[60954] = {-9'd66,10'd135};
ram[60955] = {-9'd63,10'd138};
ram[60956] = {-9'd59,10'd141};
ram[60957] = {-9'd56,10'd144};
ram[60958] = {-9'd53,10'd147};
ram[60959] = {-9'd50,10'd150};
ram[60960] = {-9'd47,10'd153};
ram[60961] = {-9'd44,10'd157};
ram[60962] = {-9'd41,10'd160};
ram[60963] = {-9'd37,10'd163};
ram[60964] = {-9'd34,10'd166};
ram[60965] = {-9'd31,10'd169};
ram[60966] = {-9'd28,10'd172};
ram[60967] = {-9'd25,10'd175};
ram[60968] = {-9'd22,10'd179};
ram[60969] = {-9'd19,10'd182};
ram[60970] = {-9'd15,10'd185};
ram[60971] = {-9'd12,10'd188};
ram[60972] = {-9'd9,10'd191};
ram[60973] = {-9'd6,10'd194};
ram[60974] = {-9'd3,10'd197};
ram[60975] = {9'd0,10'd201};
ram[60976] = {9'd3,10'd204};
ram[60977] = {9'd7,10'd207};
ram[60978] = {9'd10,10'd210};
ram[60979] = {9'd13,10'd213};
ram[60980] = {9'd16,10'd216};
ram[60981] = {9'd19,10'd219};
ram[60982] = {9'd22,10'd223};
ram[60983] = {9'd25,10'd226};
ram[60984] = {9'd29,10'd229};
ram[60985] = {9'd32,10'd232};
ram[60986] = {9'd35,10'd235};
ram[60987] = {9'd38,10'd238};
ram[60988] = {9'd41,10'd241};
ram[60989] = {9'd44,10'd245};
ram[60990] = {9'd47,10'd248};
ram[60991] = {9'd51,10'd251};
ram[60992] = {9'd54,10'd254};
ram[60993] = {9'd57,10'd257};
ram[60994] = {9'd60,10'd260};
ram[60995] = {9'd63,10'd263};
ram[60996] = {9'd66,10'd267};
ram[60997] = {9'd69,10'd270};
ram[60998] = {9'd73,10'd273};
ram[60999] = {9'd76,10'd276};
ram[61000] = {9'd79,10'd279};
ram[61001] = {9'd82,10'd282};
ram[61002] = {9'd85,10'd285};
ram[61003] = {9'd88,10'd289};
ram[61004] = {9'd91,10'd292};
ram[61005] = {9'd95,10'd295};
ram[61006] = {9'd98,10'd298};
ram[61007] = {-9'd99,10'd301};
ram[61008] = {-9'd96,10'd304};
ram[61009] = {-9'd93,10'd307};
ram[61010] = {-9'd90,10'd311};
ram[61011] = {-9'd87,10'd314};
ram[61012] = {-9'd84,10'd317};
ram[61013] = {-9'd81,10'd320};
ram[61014] = {-9'd77,10'd323};
ram[61015] = {-9'd74,10'd326};
ram[61016] = {-9'd71,10'd329};
ram[61017] = {-9'd68,10'd333};
ram[61018] = {-9'd65,10'd336};
ram[61019] = {-9'd62,10'd339};
ram[61020] = {-9'd59,10'd342};
ram[61021] = {-9'd55,10'd345};
ram[61022] = {-9'd52,10'd348};
ram[61023] = {-9'd49,10'd351};
ram[61024] = {-9'd46,10'd354};
ram[61025] = {-9'd43,10'd358};
ram[61026] = {-9'd40,10'd361};
ram[61027] = {-9'd37,10'd364};
ram[61028] = {-9'd33,10'd367};
ram[61029] = {-9'd30,10'd370};
ram[61030] = {-9'd27,10'd373};
ram[61031] = {-9'd24,10'd376};
ram[61032] = {-9'd21,10'd380};
ram[61033] = {-9'd18,10'd383};
ram[61034] = {-9'd15,10'd386};
ram[61035] = {-9'd11,10'd389};
ram[61036] = {-9'd8,10'd392};
ram[61037] = {-9'd5,10'd395};
ram[61038] = {-9'd2,10'd398};
ram[61039] = {9'd1,-10'd399};
ram[61040] = {9'd4,-10'd396};
ram[61041] = {9'd7,-10'd393};
ram[61042] = {9'd10,-10'd390};
ram[61043] = {9'd14,-10'd387};
ram[61044] = {9'd17,-10'd384};
ram[61045] = {9'd20,-10'd381};
ram[61046] = {9'd23,-10'd377};
ram[61047] = {9'd26,-10'd374};
ram[61048] = {9'd29,-10'd371};
ram[61049] = {9'd32,-10'd368};
ram[61050] = {9'd36,-10'd365};
ram[61051] = {9'd39,-10'd362};
ram[61052] = {9'd42,-10'd359};
ram[61053] = {9'd45,-10'd355};
ram[61054] = {9'd48,-10'd352};
ram[61055] = {9'd51,-10'd349};
ram[61056] = {9'd51,-10'd349};
ram[61057] = {9'd54,-10'd346};
ram[61058] = {9'd58,-10'd343};
ram[61059] = {9'd61,-10'd340};
ram[61060] = {9'd64,-10'd337};
ram[61061] = {9'd67,-10'd334};
ram[61062] = {9'd70,-10'd330};
ram[61063] = {9'd73,-10'd327};
ram[61064] = {9'd76,-10'd324};
ram[61065] = {9'd80,-10'd321};
ram[61066] = {9'd83,-10'd318};
ram[61067] = {9'd86,-10'd315};
ram[61068] = {9'd89,-10'd312};
ram[61069] = {9'd92,-10'd308};
ram[61070] = {9'd95,-10'd305};
ram[61071] = {9'd98,-10'd302};
ram[61072] = {-9'd99,-10'd299};
ram[61073] = {-9'd96,-10'd296};
ram[61074] = {-9'd92,-10'd293};
ram[61075] = {-9'd89,-10'd290};
ram[61076] = {-9'd86,-10'd286};
ram[61077] = {-9'd83,-10'd283};
ram[61078] = {-9'd80,-10'd280};
ram[61079] = {-9'd77,-10'd277};
ram[61080] = {-9'd74,-10'd274};
ram[61081] = {-9'd70,-10'd271};
ram[61082] = {-9'd67,-10'd268};
ram[61083] = {-9'd64,-10'd264};
ram[61084] = {-9'd61,-10'd261};
ram[61085] = {-9'd58,-10'd258};
ram[61086] = {-9'd55,-10'd255};
ram[61087] = {-9'd52,-10'd252};
ram[61088] = {-9'd48,-10'd249};
ram[61089] = {-9'd45,-10'd246};
ram[61090] = {-9'd42,-10'd242};
ram[61091] = {-9'd39,-10'd239};
ram[61092] = {-9'd36,-10'd236};
ram[61093] = {-9'd33,-10'd233};
ram[61094] = {-9'd30,-10'd230};
ram[61095] = {-9'd26,-10'd227};
ram[61096] = {-9'd23,-10'd224};
ram[61097] = {-9'd20,-10'd220};
ram[61098] = {-9'd17,-10'd217};
ram[61099] = {-9'd14,-10'd214};
ram[61100] = {-9'd11,-10'd211};
ram[61101] = {-9'd8,-10'd208};
ram[61102] = {-9'd4,-10'd205};
ram[61103] = {-9'd1,-10'd202};
ram[61104] = {9'd2,-10'd198};
ram[61105] = {9'd5,-10'd195};
ram[61106] = {9'd8,-10'd192};
ram[61107] = {9'd11,-10'd189};
ram[61108] = {9'd14,-10'd186};
ram[61109] = {9'd18,-10'd183};
ram[61110] = {9'd21,-10'd180};
ram[61111] = {9'd24,-10'd176};
ram[61112] = {9'd27,-10'd173};
ram[61113] = {9'd30,-10'd170};
ram[61114] = {9'd33,-10'd167};
ram[61115] = {9'd36,-10'd164};
ram[61116] = {9'd40,-10'd161};
ram[61117] = {9'd43,-10'd158};
ram[61118] = {9'd46,-10'd154};
ram[61119] = {9'd49,-10'd151};
ram[61120] = {9'd52,-10'd148};
ram[61121] = {9'd55,-10'd145};
ram[61122] = {9'd58,-10'd142};
ram[61123] = {9'd62,-10'd139};
ram[61124] = {9'd65,-10'd136};
ram[61125] = {9'd68,-10'd132};
ram[61126] = {9'd71,-10'd129};
ram[61127] = {9'd74,-10'd126};
ram[61128] = {9'd77,-10'd123};
ram[61129] = {9'd80,-10'd120};
ram[61130] = {9'd84,-10'd117};
ram[61131] = {9'd87,-10'd114};
ram[61132] = {9'd90,-10'd110};
ram[61133] = {9'd93,-10'd107};
ram[61134] = {9'd96,-10'd104};
ram[61135] = {9'd99,-10'd101};
ram[61136] = {-9'd98,-10'd98};
ram[61137] = {-9'd95,-10'd95};
ram[61138] = {-9'd92,-10'd92};
ram[61139] = {-9'd88,-10'd88};
ram[61140] = {-9'd85,-10'd85};
ram[61141] = {-9'd82,-10'd82};
ram[61142] = {-9'd79,-10'd79};
ram[61143] = {-9'd76,-10'd76};
ram[61144] = {-9'd73,-10'd73};
ram[61145] = {-9'd70,-10'd70};
ram[61146] = {-9'd66,-10'd66};
ram[61147] = {-9'd63,-10'd63};
ram[61148] = {-9'd60,-10'd60};
ram[61149] = {-9'd57,-10'd57};
ram[61150] = {-9'd54,-10'd54};
ram[61151] = {-9'd51,-10'd51};
ram[61152] = {-9'd48,-10'd48};
ram[61153] = {-9'd44,-10'd44};
ram[61154] = {-9'd41,-10'd41};
ram[61155] = {-9'd38,-10'd38};
ram[61156] = {-9'd35,-10'd35};
ram[61157] = {-9'd32,-10'd32};
ram[61158] = {-9'd29,-10'd29};
ram[61159] = {-9'd26,-10'd26};
ram[61160] = {-9'd22,-10'd22};
ram[61161] = {-9'd19,-10'd19};
ram[61162] = {-9'd16,-10'd16};
ram[61163] = {-9'd13,-10'd13};
ram[61164] = {-9'd10,-10'd10};
ram[61165] = {-9'd7,-10'd7};
ram[61166] = {-9'd4,-10'd4};
ram[61167] = {9'd0,10'd0};
ram[61168] = {9'd3,10'd3};
ram[61169] = {9'd6,10'd6};
ram[61170] = {9'd9,10'd9};
ram[61171] = {9'd12,10'd12};
ram[61172] = {9'd15,10'd15};
ram[61173] = {9'd18,10'd18};
ram[61174] = {9'd21,10'd21};
ram[61175] = {9'd25,10'd25};
ram[61176] = {9'd28,10'd28};
ram[61177] = {9'd31,10'd31};
ram[61178] = {9'd34,10'd34};
ram[61179] = {9'd37,10'd37};
ram[61180] = {9'd40,10'd40};
ram[61181] = {9'd43,10'd43};
ram[61182] = {9'd47,10'd47};
ram[61183] = {9'd50,10'd50};
ram[61184] = {9'd50,10'd50};
ram[61185] = {9'd53,10'd53};
ram[61186] = {9'd56,10'd56};
ram[61187] = {9'd59,10'd59};
ram[61188] = {9'd62,10'd62};
ram[61189] = {9'd65,10'd65};
ram[61190] = {9'd69,10'd69};
ram[61191] = {9'd72,10'd72};
ram[61192] = {9'd75,10'd75};
ram[61193] = {9'd78,10'd78};
ram[61194] = {9'd81,10'd81};
ram[61195] = {9'd84,10'd84};
ram[61196] = {9'd87,10'd87};
ram[61197] = {9'd91,10'd91};
ram[61198] = {9'd94,10'd94};
ram[61199] = {9'd97,10'd97};
ram[61200] = {-9'd100,10'd100};
ram[61201] = {-9'd97,10'd103};
ram[61202] = {-9'd94,10'd106};
ram[61203] = {-9'd91,10'd109};
ram[61204] = {-9'd88,10'd113};
ram[61205] = {-9'd85,10'd116};
ram[61206] = {-9'd81,10'd119};
ram[61207] = {-9'd78,10'd122};
ram[61208] = {-9'd75,10'd125};
ram[61209] = {-9'd72,10'd128};
ram[61210] = {-9'd69,10'd131};
ram[61211] = {-9'd66,10'd135};
ram[61212] = {-9'd63,10'd138};
ram[61213] = {-9'd59,10'd141};
ram[61214] = {-9'd56,10'd144};
ram[61215] = {-9'd53,10'd147};
ram[61216] = {-9'd50,10'd150};
ram[61217] = {-9'd47,10'd153};
ram[61218] = {-9'd44,10'd157};
ram[61219] = {-9'd41,10'd160};
ram[61220] = {-9'd37,10'd163};
ram[61221] = {-9'd34,10'd166};
ram[61222] = {-9'd31,10'd169};
ram[61223] = {-9'd28,10'd172};
ram[61224] = {-9'd25,10'd175};
ram[61225] = {-9'd22,10'd179};
ram[61226] = {-9'd19,10'd182};
ram[61227] = {-9'd15,10'd185};
ram[61228] = {-9'd12,10'd188};
ram[61229] = {-9'd9,10'd191};
ram[61230] = {-9'd6,10'd194};
ram[61231] = {-9'd3,10'd197};
ram[61232] = {9'd0,10'd201};
ram[61233] = {9'd3,10'd204};
ram[61234] = {9'd7,10'd207};
ram[61235] = {9'd10,10'd210};
ram[61236] = {9'd13,10'd213};
ram[61237] = {9'd16,10'd216};
ram[61238] = {9'd19,10'd219};
ram[61239] = {9'd22,10'd223};
ram[61240] = {9'd25,10'd226};
ram[61241] = {9'd29,10'd229};
ram[61242] = {9'd32,10'd232};
ram[61243] = {9'd35,10'd235};
ram[61244] = {9'd38,10'd238};
ram[61245] = {9'd41,10'd241};
ram[61246] = {9'd44,10'd245};
ram[61247] = {9'd47,10'd248};
ram[61248] = {9'd51,10'd251};
ram[61249] = {9'd54,10'd254};
ram[61250] = {9'd57,10'd257};
ram[61251] = {9'd60,10'd260};
ram[61252] = {9'd63,10'd263};
ram[61253] = {9'd66,10'd267};
ram[61254] = {9'd69,10'd270};
ram[61255] = {9'd73,10'd273};
ram[61256] = {9'd76,10'd276};
ram[61257] = {9'd79,10'd279};
ram[61258] = {9'd82,10'd282};
ram[61259] = {9'd85,10'd285};
ram[61260] = {9'd88,10'd289};
ram[61261] = {9'd91,10'd292};
ram[61262] = {9'd95,10'd295};
ram[61263] = {9'd98,10'd298};
ram[61264] = {-9'd99,10'd301};
ram[61265] = {-9'd96,10'd304};
ram[61266] = {-9'd93,10'd307};
ram[61267] = {-9'd90,10'd311};
ram[61268] = {-9'd87,10'd314};
ram[61269] = {-9'd84,10'd317};
ram[61270] = {-9'd81,10'd320};
ram[61271] = {-9'd77,10'd323};
ram[61272] = {-9'd74,10'd326};
ram[61273] = {-9'd71,10'd329};
ram[61274] = {-9'd68,10'd333};
ram[61275] = {-9'd65,10'd336};
ram[61276] = {-9'd62,10'd339};
ram[61277] = {-9'd59,10'd342};
ram[61278] = {-9'd55,10'd345};
ram[61279] = {-9'd52,10'd348};
ram[61280] = {-9'd49,10'd351};
ram[61281] = {-9'd46,10'd354};
ram[61282] = {-9'd43,10'd358};
ram[61283] = {-9'd40,10'd361};
ram[61284] = {-9'd37,10'd364};
ram[61285] = {-9'd33,10'd367};
ram[61286] = {-9'd30,10'd370};
ram[61287] = {-9'd27,10'd373};
ram[61288] = {-9'd24,10'd376};
ram[61289] = {-9'd21,10'd380};
ram[61290] = {-9'd18,10'd383};
ram[61291] = {-9'd15,10'd386};
ram[61292] = {-9'd11,10'd389};
ram[61293] = {-9'd8,10'd392};
ram[61294] = {-9'd5,10'd395};
ram[61295] = {-9'd2,10'd398};
ram[61296] = {9'd1,-10'd399};
ram[61297] = {9'd4,-10'd396};
ram[61298] = {9'd7,-10'd393};
ram[61299] = {9'd10,-10'd390};
ram[61300] = {9'd14,-10'd387};
ram[61301] = {9'd17,-10'd384};
ram[61302] = {9'd20,-10'd381};
ram[61303] = {9'd23,-10'd377};
ram[61304] = {9'd26,-10'd374};
ram[61305] = {9'd29,-10'd371};
ram[61306] = {9'd32,-10'd368};
ram[61307] = {9'd36,-10'd365};
ram[61308] = {9'd39,-10'd362};
ram[61309] = {9'd42,-10'd359};
ram[61310] = {9'd45,-10'd355};
ram[61311] = {9'd48,-10'd352};
ram[61312] = {9'd48,-10'd352};
ram[61313] = {9'd51,-10'd349};
ram[61314] = {9'd54,-10'd346};
ram[61315] = {9'd58,-10'd343};
ram[61316] = {9'd61,-10'd340};
ram[61317] = {9'd64,-10'd337};
ram[61318] = {9'd67,-10'd334};
ram[61319] = {9'd70,-10'd330};
ram[61320] = {9'd73,-10'd327};
ram[61321] = {9'd76,-10'd324};
ram[61322] = {9'd80,-10'd321};
ram[61323] = {9'd83,-10'd318};
ram[61324] = {9'd86,-10'd315};
ram[61325] = {9'd89,-10'd312};
ram[61326] = {9'd92,-10'd308};
ram[61327] = {9'd95,-10'd305};
ram[61328] = {9'd98,-10'd302};
ram[61329] = {-9'd99,-10'd299};
ram[61330] = {-9'd96,-10'd296};
ram[61331] = {-9'd92,-10'd293};
ram[61332] = {-9'd89,-10'd290};
ram[61333] = {-9'd86,-10'd286};
ram[61334] = {-9'd83,-10'd283};
ram[61335] = {-9'd80,-10'd280};
ram[61336] = {-9'd77,-10'd277};
ram[61337] = {-9'd74,-10'd274};
ram[61338] = {-9'd70,-10'd271};
ram[61339] = {-9'd67,-10'd268};
ram[61340] = {-9'd64,-10'd264};
ram[61341] = {-9'd61,-10'd261};
ram[61342] = {-9'd58,-10'd258};
ram[61343] = {-9'd55,-10'd255};
ram[61344] = {-9'd52,-10'd252};
ram[61345] = {-9'd48,-10'd249};
ram[61346] = {-9'd45,-10'd246};
ram[61347] = {-9'd42,-10'd242};
ram[61348] = {-9'd39,-10'd239};
ram[61349] = {-9'd36,-10'd236};
ram[61350] = {-9'd33,-10'd233};
ram[61351] = {-9'd30,-10'd230};
ram[61352] = {-9'd26,-10'd227};
ram[61353] = {-9'd23,-10'd224};
ram[61354] = {-9'd20,-10'd220};
ram[61355] = {-9'd17,-10'd217};
ram[61356] = {-9'd14,-10'd214};
ram[61357] = {-9'd11,-10'd211};
ram[61358] = {-9'd8,-10'd208};
ram[61359] = {-9'd4,-10'd205};
ram[61360] = {-9'd1,-10'd202};
ram[61361] = {9'd2,-10'd198};
ram[61362] = {9'd5,-10'd195};
ram[61363] = {9'd8,-10'd192};
ram[61364] = {9'd11,-10'd189};
ram[61365] = {9'd14,-10'd186};
ram[61366] = {9'd18,-10'd183};
ram[61367] = {9'd21,-10'd180};
ram[61368] = {9'd24,-10'd176};
ram[61369] = {9'd27,-10'd173};
ram[61370] = {9'd30,-10'd170};
ram[61371] = {9'd33,-10'd167};
ram[61372] = {9'd36,-10'd164};
ram[61373] = {9'd40,-10'd161};
ram[61374] = {9'd43,-10'd158};
ram[61375] = {9'd46,-10'd154};
ram[61376] = {9'd49,-10'd151};
ram[61377] = {9'd52,-10'd148};
ram[61378] = {9'd55,-10'd145};
ram[61379] = {9'd58,-10'd142};
ram[61380] = {9'd62,-10'd139};
ram[61381] = {9'd65,-10'd136};
ram[61382] = {9'd68,-10'd132};
ram[61383] = {9'd71,-10'd129};
ram[61384] = {9'd74,-10'd126};
ram[61385] = {9'd77,-10'd123};
ram[61386] = {9'd80,-10'd120};
ram[61387] = {9'd84,-10'd117};
ram[61388] = {9'd87,-10'd114};
ram[61389] = {9'd90,-10'd110};
ram[61390] = {9'd93,-10'd107};
ram[61391] = {9'd96,-10'd104};
ram[61392] = {9'd99,-10'd101};
ram[61393] = {-9'd98,-10'd98};
ram[61394] = {-9'd95,-10'd95};
ram[61395] = {-9'd92,-10'd92};
ram[61396] = {-9'd88,-10'd88};
ram[61397] = {-9'd85,-10'd85};
ram[61398] = {-9'd82,-10'd82};
ram[61399] = {-9'd79,-10'd79};
ram[61400] = {-9'd76,-10'd76};
ram[61401] = {-9'd73,-10'd73};
ram[61402] = {-9'd70,-10'd70};
ram[61403] = {-9'd66,-10'd66};
ram[61404] = {-9'd63,-10'd63};
ram[61405] = {-9'd60,-10'd60};
ram[61406] = {-9'd57,-10'd57};
ram[61407] = {-9'd54,-10'd54};
ram[61408] = {-9'd51,-10'd51};
ram[61409] = {-9'd48,-10'd48};
ram[61410] = {-9'd44,-10'd44};
ram[61411] = {-9'd41,-10'd41};
ram[61412] = {-9'd38,-10'd38};
ram[61413] = {-9'd35,-10'd35};
ram[61414] = {-9'd32,-10'd32};
ram[61415] = {-9'd29,-10'd29};
ram[61416] = {-9'd26,-10'd26};
ram[61417] = {-9'd22,-10'd22};
ram[61418] = {-9'd19,-10'd19};
ram[61419] = {-9'd16,-10'd16};
ram[61420] = {-9'd13,-10'd13};
ram[61421] = {-9'd10,-10'd10};
ram[61422] = {-9'd7,-10'd7};
ram[61423] = {-9'd4,-10'd4};
ram[61424] = {9'd0,10'd0};
ram[61425] = {9'd3,10'd3};
ram[61426] = {9'd6,10'd6};
ram[61427] = {9'd9,10'd9};
ram[61428] = {9'd12,10'd12};
ram[61429] = {9'd15,10'd15};
ram[61430] = {9'd18,10'd18};
ram[61431] = {9'd21,10'd21};
ram[61432] = {9'd25,10'd25};
ram[61433] = {9'd28,10'd28};
ram[61434] = {9'd31,10'd31};
ram[61435] = {9'd34,10'd34};
ram[61436] = {9'd37,10'd37};
ram[61437] = {9'd40,10'd40};
ram[61438] = {9'd43,10'd43};
ram[61439] = {9'd47,10'd47};
ram[61440] = {9'd47,10'd47};
ram[61441] = {9'd50,10'd50};
ram[61442] = {9'd53,10'd53};
ram[61443] = {9'd56,10'd56};
ram[61444] = {9'd59,10'd59};
ram[61445] = {9'd62,10'd62};
ram[61446] = {9'd65,10'd65};
ram[61447] = {9'd69,10'd69};
ram[61448] = {9'd72,10'd72};
ram[61449] = {9'd75,10'd75};
ram[61450] = {9'd78,10'd78};
ram[61451] = {9'd81,10'd81};
ram[61452] = {9'd84,10'd84};
ram[61453] = {9'd87,10'd87};
ram[61454] = {9'd91,10'd91};
ram[61455] = {9'd94,10'd94};
ram[61456] = {9'd97,10'd97};
ram[61457] = {-9'd100,10'd100};
ram[61458] = {-9'd97,10'd103};
ram[61459] = {-9'd94,10'd106};
ram[61460] = {-9'd91,10'd109};
ram[61461] = {-9'd88,10'd113};
ram[61462] = {-9'd85,10'd116};
ram[61463] = {-9'd81,10'd119};
ram[61464] = {-9'd78,10'd122};
ram[61465] = {-9'd75,10'd125};
ram[61466] = {-9'd72,10'd128};
ram[61467] = {-9'd69,10'd131};
ram[61468] = {-9'd66,10'd135};
ram[61469] = {-9'd63,10'd138};
ram[61470] = {-9'd59,10'd141};
ram[61471] = {-9'd56,10'd144};
ram[61472] = {-9'd53,10'd147};
ram[61473] = {-9'd50,10'd150};
ram[61474] = {-9'd47,10'd153};
ram[61475] = {-9'd44,10'd157};
ram[61476] = {-9'd41,10'd160};
ram[61477] = {-9'd37,10'd163};
ram[61478] = {-9'd34,10'd166};
ram[61479] = {-9'd31,10'd169};
ram[61480] = {-9'd28,10'd172};
ram[61481] = {-9'd25,10'd175};
ram[61482] = {-9'd22,10'd179};
ram[61483] = {-9'd19,10'd182};
ram[61484] = {-9'd15,10'd185};
ram[61485] = {-9'd12,10'd188};
ram[61486] = {-9'd9,10'd191};
ram[61487] = {-9'd6,10'd194};
ram[61488] = {-9'd3,10'd197};
ram[61489] = {9'd0,10'd201};
ram[61490] = {9'd3,10'd204};
ram[61491] = {9'd7,10'd207};
ram[61492] = {9'd10,10'd210};
ram[61493] = {9'd13,10'd213};
ram[61494] = {9'd16,10'd216};
ram[61495] = {9'd19,10'd219};
ram[61496] = {9'd22,10'd223};
ram[61497] = {9'd25,10'd226};
ram[61498] = {9'd29,10'd229};
ram[61499] = {9'd32,10'd232};
ram[61500] = {9'd35,10'd235};
ram[61501] = {9'd38,10'd238};
ram[61502] = {9'd41,10'd241};
ram[61503] = {9'd44,10'd245};
ram[61504] = {9'd47,10'd248};
ram[61505] = {9'd51,10'd251};
ram[61506] = {9'd54,10'd254};
ram[61507] = {9'd57,10'd257};
ram[61508] = {9'd60,10'd260};
ram[61509] = {9'd63,10'd263};
ram[61510] = {9'd66,10'd267};
ram[61511] = {9'd69,10'd270};
ram[61512] = {9'd73,10'd273};
ram[61513] = {9'd76,10'd276};
ram[61514] = {9'd79,10'd279};
ram[61515] = {9'd82,10'd282};
ram[61516] = {9'd85,10'd285};
ram[61517] = {9'd88,10'd289};
ram[61518] = {9'd91,10'd292};
ram[61519] = {9'd95,10'd295};
ram[61520] = {9'd98,10'd298};
ram[61521] = {-9'd99,10'd301};
ram[61522] = {-9'd96,10'd304};
ram[61523] = {-9'd93,10'd307};
ram[61524] = {-9'd90,10'd311};
ram[61525] = {-9'd87,10'd314};
ram[61526] = {-9'd84,10'd317};
ram[61527] = {-9'd81,10'd320};
ram[61528] = {-9'd77,10'd323};
ram[61529] = {-9'd74,10'd326};
ram[61530] = {-9'd71,10'd329};
ram[61531] = {-9'd68,10'd333};
ram[61532] = {-9'd65,10'd336};
ram[61533] = {-9'd62,10'd339};
ram[61534] = {-9'd59,10'd342};
ram[61535] = {-9'd55,10'd345};
ram[61536] = {-9'd52,10'd348};
ram[61537] = {-9'd49,10'd351};
ram[61538] = {-9'd46,10'd354};
ram[61539] = {-9'd43,10'd358};
ram[61540] = {-9'd40,10'd361};
ram[61541] = {-9'd37,10'd364};
ram[61542] = {-9'd33,10'd367};
ram[61543] = {-9'd30,10'd370};
ram[61544] = {-9'd27,10'd373};
ram[61545] = {-9'd24,10'd376};
ram[61546] = {-9'd21,10'd380};
ram[61547] = {-9'd18,10'd383};
ram[61548] = {-9'd15,10'd386};
ram[61549] = {-9'd11,10'd389};
ram[61550] = {-9'd8,10'd392};
ram[61551] = {-9'd5,10'd395};
ram[61552] = {-9'd2,10'd398};
ram[61553] = {9'd1,-10'd399};
ram[61554] = {9'd4,-10'd396};
ram[61555] = {9'd7,-10'd393};
ram[61556] = {9'd10,-10'd390};
ram[61557] = {9'd14,-10'd387};
ram[61558] = {9'd17,-10'd384};
ram[61559] = {9'd20,-10'd381};
ram[61560] = {9'd23,-10'd377};
ram[61561] = {9'd26,-10'd374};
ram[61562] = {9'd29,-10'd371};
ram[61563] = {9'd32,-10'd368};
ram[61564] = {9'd36,-10'd365};
ram[61565] = {9'd39,-10'd362};
ram[61566] = {9'd42,-10'd359};
ram[61567] = {9'd45,-10'd355};
ram[61568] = {9'd45,-10'd355};
ram[61569] = {9'd48,-10'd352};
ram[61570] = {9'd51,-10'd349};
ram[61571] = {9'd54,-10'd346};
ram[61572] = {9'd58,-10'd343};
ram[61573] = {9'd61,-10'd340};
ram[61574] = {9'd64,-10'd337};
ram[61575] = {9'd67,-10'd334};
ram[61576] = {9'd70,-10'd330};
ram[61577] = {9'd73,-10'd327};
ram[61578] = {9'd76,-10'd324};
ram[61579] = {9'd80,-10'd321};
ram[61580] = {9'd83,-10'd318};
ram[61581] = {9'd86,-10'd315};
ram[61582] = {9'd89,-10'd312};
ram[61583] = {9'd92,-10'd308};
ram[61584] = {9'd95,-10'd305};
ram[61585] = {9'd98,-10'd302};
ram[61586] = {-9'd99,-10'd299};
ram[61587] = {-9'd96,-10'd296};
ram[61588] = {-9'd92,-10'd293};
ram[61589] = {-9'd89,-10'd290};
ram[61590] = {-9'd86,-10'd286};
ram[61591] = {-9'd83,-10'd283};
ram[61592] = {-9'd80,-10'd280};
ram[61593] = {-9'd77,-10'd277};
ram[61594] = {-9'd74,-10'd274};
ram[61595] = {-9'd70,-10'd271};
ram[61596] = {-9'd67,-10'd268};
ram[61597] = {-9'd64,-10'd264};
ram[61598] = {-9'd61,-10'd261};
ram[61599] = {-9'd58,-10'd258};
ram[61600] = {-9'd55,-10'd255};
ram[61601] = {-9'd52,-10'd252};
ram[61602] = {-9'd48,-10'd249};
ram[61603] = {-9'd45,-10'd246};
ram[61604] = {-9'd42,-10'd242};
ram[61605] = {-9'd39,-10'd239};
ram[61606] = {-9'd36,-10'd236};
ram[61607] = {-9'd33,-10'd233};
ram[61608] = {-9'd30,-10'd230};
ram[61609] = {-9'd26,-10'd227};
ram[61610] = {-9'd23,-10'd224};
ram[61611] = {-9'd20,-10'd220};
ram[61612] = {-9'd17,-10'd217};
ram[61613] = {-9'd14,-10'd214};
ram[61614] = {-9'd11,-10'd211};
ram[61615] = {-9'd8,-10'd208};
ram[61616] = {-9'd4,-10'd205};
ram[61617] = {-9'd1,-10'd202};
ram[61618] = {9'd2,-10'd198};
ram[61619] = {9'd5,-10'd195};
ram[61620] = {9'd8,-10'd192};
ram[61621] = {9'd11,-10'd189};
ram[61622] = {9'd14,-10'd186};
ram[61623] = {9'd18,-10'd183};
ram[61624] = {9'd21,-10'd180};
ram[61625] = {9'd24,-10'd176};
ram[61626] = {9'd27,-10'd173};
ram[61627] = {9'd30,-10'd170};
ram[61628] = {9'd33,-10'd167};
ram[61629] = {9'd36,-10'd164};
ram[61630] = {9'd40,-10'd161};
ram[61631] = {9'd43,-10'd158};
ram[61632] = {9'd46,-10'd154};
ram[61633] = {9'd49,-10'd151};
ram[61634] = {9'd52,-10'd148};
ram[61635] = {9'd55,-10'd145};
ram[61636] = {9'd58,-10'd142};
ram[61637] = {9'd62,-10'd139};
ram[61638] = {9'd65,-10'd136};
ram[61639] = {9'd68,-10'd132};
ram[61640] = {9'd71,-10'd129};
ram[61641] = {9'd74,-10'd126};
ram[61642] = {9'd77,-10'd123};
ram[61643] = {9'd80,-10'd120};
ram[61644] = {9'd84,-10'd117};
ram[61645] = {9'd87,-10'd114};
ram[61646] = {9'd90,-10'd110};
ram[61647] = {9'd93,-10'd107};
ram[61648] = {9'd96,-10'd104};
ram[61649] = {9'd99,-10'd101};
ram[61650] = {-9'd98,-10'd98};
ram[61651] = {-9'd95,-10'd95};
ram[61652] = {-9'd92,-10'd92};
ram[61653] = {-9'd88,-10'd88};
ram[61654] = {-9'd85,-10'd85};
ram[61655] = {-9'd82,-10'd82};
ram[61656] = {-9'd79,-10'd79};
ram[61657] = {-9'd76,-10'd76};
ram[61658] = {-9'd73,-10'd73};
ram[61659] = {-9'd70,-10'd70};
ram[61660] = {-9'd66,-10'd66};
ram[61661] = {-9'd63,-10'd63};
ram[61662] = {-9'd60,-10'd60};
ram[61663] = {-9'd57,-10'd57};
ram[61664] = {-9'd54,-10'd54};
ram[61665] = {-9'd51,-10'd51};
ram[61666] = {-9'd48,-10'd48};
ram[61667] = {-9'd44,-10'd44};
ram[61668] = {-9'd41,-10'd41};
ram[61669] = {-9'd38,-10'd38};
ram[61670] = {-9'd35,-10'd35};
ram[61671] = {-9'd32,-10'd32};
ram[61672] = {-9'd29,-10'd29};
ram[61673] = {-9'd26,-10'd26};
ram[61674] = {-9'd22,-10'd22};
ram[61675] = {-9'd19,-10'd19};
ram[61676] = {-9'd16,-10'd16};
ram[61677] = {-9'd13,-10'd13};
ram[61678] = {-9'd10,-10'd10};
ram[61679] = {-9'd7,-10'd7};
ram[61680] = {-9'd4,-10'd4};
ram[61681] = {9'd0,10'd0};
ram[61682] = {9'd3,10'd3};
ram[61683] = {9'd6,10'd6};
ram[61684] = {9'd9,10'd9};
ram[61685] = {9'd12,10'd12};
ram[61686] = {9'd15,10'd15};
ram[61687] = {9'd18,10'd18};
ram[61688] = {9'd21,10'd21};
ram[61689] = {9'd25,10'd25};
ram[61690] = {9'd28,10'd28};
ram[61691] = {9'd31,10'd31};
ram[61692] = {9'd34,10'd34};
ram[61693] = {9'd37,10'd37};
ram[61694] = {9'd40,10'd40};
ram[61695] = {9'd43,10'd43};
ram[61696] = {9'd43,10'd43};
ram[61697] = {9'd47,10'd47};
ram[61698] = {9'd50,10'd50};
ram[61699] = {9'd53,10'd53};
ram[61700] = {9'd56,10'd56};
ram[61701] = {9'd59,10'd59};
ram[61702] = {9'd62,10'd62};
ram[61703] = {9'd65,10'd65};
ram[61704] = {9'd69,10'd69};
ram[61705] = {9'd72,10'd72};
ram[61706] = {9'd75,10'd75};
ram[61707] = {9'd78,10'd78};
ram[61708] = {9'd81,10'd81};
ram[61709] = {9'd84,10'd84};
ram[61710] = {9'd87,10'd87};
ram[61711] = {9'd91,10'd91};
ram[61712] = {9'd94,10'd94};
ram[61713] = {9'd97,10'd97};
ram[61714] = {-9'd100,10'd100};
ram[61715] = {-9'd97,10'd103};
ram[61716] = {-9'd94,10'd106};
ram[61717] = {-9'd91,10'd109};
ram[61718] = {-9'd88,10'd113};
ram[61719] = {-9'd85,10'd116};
ram[61720] = {-9'd81,10'd119};
ram[61721] = {-9'd78,10'd122};
ram[61722] = {-9'd75,10'd125};
ram[61723] = {-9'd72,10'd128};
ram[61724] = {-9'd69,10'd131};
ram[61725] = {-9'd66,10'd135};
ram[61726] = {-9'd63,10'd138};
ram[61727] = {-9'd59,10'd141};
ram[61728] = {-9'd56,10'd144};
ram[61729] = {-9'd53,10'd147};
ram[61730] = {-9'd50,10'd150};
ram[61731] = {-9'd47,10'd153};
ram[61732] = {-9'd44,10'd157};
ram[61733] = {-9'd41,10'd160};
ram[61734] = {-9'd37,10'd163};
ram[61735] = {-9'd34,10'd166};
ram[61736] = {-9'd31,10'd169};
ram[61737] = {-9'd28,10'd172};
ram[61738] = {-9'd25,10'd175};
ram[61739] = {-9'd22,10'd179};
ram[61740] = {-9'd19,10'd182};
ram[61741] = {-9'd15,10'd185};
ram[61742] = {-9'd12,10'd188};
ram[61743] = {-9'd9,10'd191};
ram[61744] = {-9'd6,10'd194};
ram[61745] = {-9'd3,10'd197};
ram[61746] = {9'd0,10'd201};
ram[61747] = {9'd3,10'd204};
ram[61748] = {9'd7,10'd207};
ram[61749] = {9'd10,10'd210};
ram[61750] = {9'd13,10'd213};
ram[61751] = {9'd16,10'd216};
ram[61752] = {9'd19,10'd219};
ram[61753] = {9'd22,10'd223};
ram[61754] = {9'd25,10'd226};
ram[61755] = {9'd29,10'd229};
ram[61756] = {9'd32,10'd232};
ram[61757] = {9'd35,10'd235};
ram[61758] = {9'd38,10'd238};
ram[61759] = {9'd41,10'd241};
ram[61760] = {9'd44,10'd245};
ram[61761] = {9'd47,10'd248};
ram[61762] = {9'd51,10'd251};
ram[61763] = {9'd54,10'd254};
ram[61764] = {9'd57,10'd257};
ram[61765] = {9'd60,10'd260};
ram[61766] = {9'd63,10'd263};
ram[61767] = {9'd66,10'd267};
ram[61768] = {9'd69,10'd270};
ram[61769] = {9'd73,10'd273};
ram[61770] = {9'd76,10'd276};
ram[61771] = {9'd79,10'd279};
ram[61772] = {9'd82,10'd282};
ram[61773] = {9'd85,10'd285};
ram[61774] = {9'd88,10'd289};
ram[61775] = {9'd91,10'd292};
ram[61776] = {9'd95,10'd295};
ram[61777] = {9'd98,10'd298};
ram[61778] = {-9'd99,10'd301};
ram[61779] = {-9'd96,10'd304};
ram[61780] = {-9'd93,10'd307};
ram[61781] = {-9'd90,10'd311};
ram[61782] = {-9'd87,10'd314};
ram[61783] = {-9'd84,10'd317};
ram[61784] = {-9'd81,10'd320};
ram[61785] = {-9'd77,10'd323};
ram[61786] = {-9'd74,10'd326};
ram[61787] = {-9'd71,10'd329};
ram[61788] = {-9'd68,10'd333};
ram[61789] = {-9'd65,10'd336};
ram[61790] = {-9'd62,10'd339};
ram[61791] = {-9'd59,10'd342};
ram[61792] = {-9'd55,10'd345};
ram[61793] = {-9'd52,10'd348};
ram[61794] = {-9'd49,10'd351};
ram[61795] = {-9'd46,10'd354};
ram[61796] = {-9'd43,10'd358};
ram[61797] = {-9'd40,10'd361};
ram[61798] = {-9'd37,10'd364};
ram[61799] = {-9'd33,10'd367};
ram[61800] = {-9'd30,10'd370};
ram[61801] = {-9'd27,10'd373};
ram[61802] = {-9'd24,10'd376};
ram[61803] = {-9'd21,10'd380};
ram[61804] = {-9'd18,10'd383};
ram[61805] = {-9'd15,10'd386};
ram[61806] = {-9'd11,10'd389};
ram[61807] = {-9'd8,10'd392};
ram[61808] = {-9'd5,10'd395};
ram[61809] = {-9'd2,10'd398};
ram[61810] = {9'd1,-10'd399};
ram[61811] = {9'd4,-10'd396};
ram[61812] = {9'd7,-10'd393};
ram[61813] = {9'd10,-10'd390};
ram[61814] = {9'd14,-10'd387};
ram[61815] = {9'd17,-10'd384};
ram[61816] = {9'd20,-10'd381};
ram[61817] = {9'd23,-10'd377};
ram[61818] = {9'd26,-10'd374};
ram[61819] = {9'd29,-10'd371};
ram[61820] = {9'd32,-10'd368};
ram[61821] = {9'd36,-10'd365};
ram[61822] = {9'd39,-10'd362};
ram[61823] = {9'd42,-10'd359};
ram[61824] = {9'd42,-10'd359};
ram[61825] = {9'd45,-10'd355};
ram[61826] = {9'd48,-10'd352};
ram[61827] = {9'd51,-10'd349};
ram[61828] = {9'd54,-10'd346};
ram[61829] = {9'd58,-10'd343};
ram[61830] = {9'd61,-10'd340};
ram[61831] = {9'd64,-10'd337};
ram[61832] = {9'd67,-10'd334};
ram[61833] = {9'd70,-10'd330};
ram[61834] = {9'd73,-10'd327};
ram[61835] = {9'd76,-10'd324};
ram[61836] = {9'd80,-10'd321};
ram[61837] = {9'd83,-10'd318};
ram[61838] = {9'd86,-10'd315};
ram[61839] = {9'd89,-10'd312};
ram[61840] = {9'd92,-10'd308};
ram[61841] = {9'd95,-10'd305};
ram[61842] = {9'd98,-10'd302};
ram[61843] = {-9'd99,-10'd299};
ram[61844] = {-9'd96,-10'd296};
ram[61845] = {-9'd92,-10'd293};
ram[61846] = {-9'd89,-10'd290};
ram[61847] = {-9'd86,-10'd286};
ram[61848] = {-9'd83,-10'd283};
ram[61849] = {-9'd80,-10'd280};
ram[61850] = {-9'd77,-10'd277};
ram[61851] = {-9'd74,-10'd274};
ram[61852] = {-9'd70,-10'd271};
ram[61853] = {-9'd67,-10'd268};
ram[61854] = {-9'd64,-10'd264};
ram[61855] = {-9'd61,-10'd261};
ram[61856] = {-9'd58,-10'd258};
ram[61857] = {-9'd55,-10'd255};
ram[61858] = {-9'd52,-10'd252};
ram[61859] = {-9'd48,-10'd249};
ram[61860] = {-9'd45,-10'd246};
ram[61861] = {-9'd42,-10'd242};
ram[61862] = {-9'd39,-10'd239};
ram[61863] = {-9'd36,-10'd236};
ram[61864] = {-9'd33,-10'd233};
ram[61865] = {-9'd30,-10'd230};
ram[61866] = {-9'd26,-10'd227};
ram[61867] = {-9'd23,-10'd224};
ram[61868] = {-9'd20,-10'd220};
ram[61869] = {-9'd17,-10'd217};
ram[61870] = {-9'd14,-10'd214};
ram[61871] = {-9'd11,-10'd211};
ram[61872] = {-9'd8,-10'd208};
ram[61873] = {-9'd4,-10'd205};
ram[61874] = {-9'd1,-10'd202};
ram[61875] = {9'd2,-10'd198};
ram[61876] = {9'd5,-10'd195};
ram[61877] = {9'd8,-10'd192};
ram[61878] = {9'd11,-10'd189};
ram[61879] = {9'd14,-10'd186};
ram[61880] = {9'd18,-10'd183};
ram[61881] = {9'd21,-10'd180};
ram[61882] = {9'd24,-10'd176};
ram[61883] = {9'd27,-10'd173};
ram[61884] = {9'd30,-10'd170};
ram[61885] = {9'd33,-10'd167};
ram[61886] = {9'd36,-10'd164};
ram[61887] = {9'd40,-10'd161};
ram[61888] = {9'd43,-10'd158};
ram[61889] = {9'd46,-10'd154};
ram[61890] = {9'd49,-10'd151};
ram[61891] = {9'd52,-10'd148};
ram[61892] = {9'd55,-10'd145};
ram[61893] = {9'd58,-10'd142};
ram[61894] = {9'd62,-10'd139};
ram[61895] = {9'd65,-10'd136};
ram[61896] = {9'd68,-10'd132};
ram[61897] = {9'd71,-10'd129};
ram[61898] = {9'd74,-10'd126};
ram[61899] = {9'd77,-10'd123};
ram[61900] = {9'd80,-10'd120};
ram[61901] = {9'd84,-10'd117};
ram[61902] = {9'd87,-10'd114};
ram[61903] = {9'd90,-10'd110};
ram[61904] = {9'd93,-10'd107};
ram[61905] = {9'd96,-10'd104};
ram[61906] = {9'd99,-10'd101};
ram[61907] = {-9'd98,-10'd98};
ram[61908] = {-9'd95,-10'd95};
ram[61909] = {-9'd92,-10'd92};
ram[61910] = {-9'd88,-10'd88};
ram[61911] = {-9'd85,-10'd85};
ram[61912] = {-9'd82,-10'd82};
ram[61913] = {-9'd79,-10'd79};
ram[61914] = {-9'd76,-10'd76};
ram[61915] = {-9'd73,-10'd73};
ram[61916] = {-9'd70,-10'd70};
ram[61917] = {-9'd66,-10'd66};
ram[61918] = {-9'd63,-10'd63};
ram[61919] = {-9'd60,-10'd60};
ram[61920] = {-9'd57,-10'd57};
ram[61921] = {-9'd54,-10'd54};
ram[61922] = {-9'd51,-10'd51};
ram[61923] = {-9'd48,-10'd48};
ram[61924] = {-9'd44,-10'd44};
ram[61925] = {-9'd41,-10'd41};
ram[61926] = {-9'd38,-10'd38};
ram[61927] = {-9'd35,-10'd35};
ram[61928] = {-9'd32,-10'd32};
ram[61929] = {-9'd29,-10'd29};
ram[61930] = {-9'd26,-10'd26};
ram[61931] = {-9'd22,-10'd22};
ram[61932] = {-9'd19,-10'd19};
ram[61933] = {-9'd16,-10'd16};
ram[61934] = {-9'd13,-10'd13};
ram[61935] = {-9'd10,-10'd10};
ram[61936] = {-9'd7,-10'd7};
ram[61937] = {-9'd4,-10'd4};
ram[61938] = {9'd0,10'd0};
ram[61939] = {9'd3,10'd3};
ram[61940] = {9'd6,10'd6};
ram[61941] = {9'd9,10'd9};
ram[61942] = {9'd12,10'd12};
ram[61943] = {9'd15,10'd15};
ram[61944] = {9'd18,10'd18};
ram[61945] = {9'd21,10'd21};
ram[61946] = {9'd25,10'd25};
ram[61947] = {9'd28,10'd28};
ram[61948] = {9'd31,10'd31};
ram[61949] = {9'd34,10'd34};
ram[61950] = {9'd37,10'd37};
ram[61951] = {9'd40,10'd40};
ram[61952] = {9'd40,10'd40};
ram[61953] = {9'd43,10'd43};
ram[61954] = {9'd47,10'd47};
ram[61955] = {9'd50,10'd50};
ram[61956] = {9'd53,10'd53};
ram[61957] = {9'd56,10'd56};
ram[61958] = {9'd59,10'd59};
ram[61959] = {9'd62,10'd62};
ram[61960] = {9'd65,10'd65};
ram[61961] = {9'd69,10'd69};
ram[61962] = {9'd72,10'd72};
ram[61963] = {9'd75,10'd75};
ram[61964] = {9'd78,10'd78};
ram[61965] = {9'd81,10'd81};
ram[61966] = {9'd84,10'd84};
ram[61967] = {9'd87,10'd87};
ram[61968] = {9'd91,10'd91};
ram[61969] = {9'd94,10'd94};
ram[61970] = {9'd97,10'd97};
ram[61971] = {-9'd100,10'd100};
ram[61972] = {-9'd97,10'd103};
ram[61973] = {-9'd94,10'd106};
ram[61974] = {-9'd91,10'd109};
ram[61975] = {-9'd88,10'd113};
ram[61976] = {-9'd85,10'd116};
ram[61977] = {-9'd81,10'd119};
ram[61978] = {-9'd78,10'd122};
ram[61979] = {-9'd75,10'd125};
ram[61980] = {-9'd72,10'd128};
ram[61981] = {-9'd69,10'd131};
ram[61982] = {-9'd66,10'd135};
ram[61983] = {-9'd63,10'd138};
ram[61984] = {-9'd59,10'd141};
ram[61985] = {-9'd56,10'd144};
ram[61986] = {-9'd53,10'd147};
ram[61987] = {-9'd50,10'd150};
ram[61988] = {-9'd47,10'd153};
ram[61989] = {-9'd44,10'd157};
ram[61990] = {-9'd41,10'd160};
ram[61991] = {-9'd37,10'd163};
ram[61992] = {-9'd34,10'd166};
ram[61993] = {-9'd31,10'd169};
ram[61994] = {-9'd28,10'd172};
ram[61995] = {-9'd25,10'd175};
ram[61996] = {-9'd22,10'd179};
ram[61997] = {-9'd19,10'd182};
ram[61998] = {-9'd15,10'd185};
ram[61999] = {-9'd12,10'd188};
ram[62000] = {-9'd9,10'd191};
ram[62001] = {-9'd6,10'd194};
ram[62002] = {-9'd3,10'd197};
ram[62003] = {9'd0,10'd201};
ram[62004] = {9'd3,10'd204};
ram[62005] = {9'd7,10'd207};
ram[62006] = {9'd10,10'd210};
ram[62007] = {9'd13,10'd213};
ram[62008] = {9'd16,10'd216};
ram[62009] = {9'd19,10'd219};
ram[62010] = {9'd22,10'd223};
ram[62011] = {9'd25,10'd226};
ram[62012] = {9'd29,10'd229};
ram[62013] = {9'd32,10'd232};
ram[62014] = {9'd35,10'd235};
ram[62015] = {9'd38,10'd238};
ram[62016] = {9'd41,10'd241};
ram[62017] = {9'd44,10'd245};
ram[62018] = {9'd47,10'd248};
ram[62019] = {9'd51,10'd251};
ram[62020] = {9'd54,10'd254};
ram[62021] = {9'd57,10'd257};
ram[62022] = {9'd60,10'd260};
ram[62023] = {9'd63,10'd263};
ram[62024] = {9'd66,10'd267};
ram[62025] = {9'd69,10'd270};
ram[62026] = {9'd73,10'd273};
ram[62027] = {9'd76,10'd276};
ram[62028] = {9'd79,10'd279};
ram[62029] = {9'd82,10'd282};
ram[62030] = {9'd85,10'd285};
ram[62031] = {9'd88,10'd289};
ram[62032] = {9'd91,10'd292};
ram[62033] = {9'd95,10'd295};
ram[62034] = {9'd98,10'd298};
ram[62035] = {-9'd99,10'd301};
ram[62036] = {-9'd96,10'd304};
ram[62037] = {-9'd93,10'd307};
ram[62038] = {-9'd90,10'd311};
ram[62039] = {-9'd87,10'd314};
ram[62040] = {-9'd84,10'd317};
ram[62041] = {-9'd81,10'd320};
ram[62042] = {-9'd77,10'd323};
ram[62043] = {-9'd74,10'd326};
ram[62044] = {-9'd71,10'd329};
ram[62045] = {-9'd68,10'd333};
ram[62046] = {-9'd65,10'd336};
ram[62047] = {-9'd62,10'd339};
ram[62048] = {-9'd59,10'd342};
ram[62049] = {-9'd55,10'd345};
ram[62050] = {-9'd52,10'd348};
ram[62051] = {-9'd49,10'd351};
ram[62052] = {-9'd46,10'd354};
ram[62053] = {-9'd43,10'd358};
ram[62054] = {-9'd40,10'd361};
ram[62055] = {-9'd37,10'd364};
ram[62056] = {-9'd33,10'd367};
ram[62057] = {-9'd30,10'd370};
ram[62058] = {-9'd27,10'd373};
ram[62059] = {-9'd24,10'd376};
ram[62060] = {-9'd21,10'd380};
ram[62061] = {-9'd18,10'd383};
ram[62062] = {-9'd15,10'd386};
ram[62063] = {-9'd11,10'd389};
ram[62064] = {-9'd8,10'd392};
ram[62065] = {-9'd5,10'd395};
ram[62066] = {-9'd2,10'd398};
ram[62067] = {9'd1,-10'd399};
ram[62068] = {9'd4,-10'd396};
ram[62069] = {9'd7,-10'd393};
ram[62070] = {9'd10,-10'd390};
ram[62071] = {9'd14,-10'd387};
ram[62072] = {9'd17,-10'd384};
ram[62073] = {9'd20,-10'd381};
ram[62074] = {9'd23,-10'd377};
ram[62075] = {9'd26,-10'd374};
ram[62076] = {9'd29,-10'd371};
ram[62077] = {9'd32,-10'd368};
ram[62078] = {9'd36,-10'd365};
ram[62079] = {9'd39,-10'd362};
ram[62080] = {9'd39,-10'd362};
ram[62081] = {9'd42,-10'd359};
ram[62082] = {9'd45,-10'd355};
ram[62083] = {9'd48,-10'd352};
ram[62084] = {9'd51,-10'd349};
ram[62085] = {9'd54,-10'd346};
ram[62086] = {9'd58,-10'd343};
ram[62087] = {9'd61,-10'd340};
ram[62088] = {9'd64,-10'd337};
ram[62089] = {9'd67,-10'd334};
ram[62090] = {9'd70,-10'd330};
ram[62091] = {9'd73,-10'd327};
ram[62092] = {9'd76,-10'd324};
ram[62093] = {9'd80,-10'd321};
ram[62094] = {9'd83,-10'd318};
ram[62095] = {9'd86,-10'd315};
ram[62096] = {9'd89,-10'd312};
ram[62097] = {9'd92,-10'd308};
ram[62098] = {9'd95,-10'd305};
ram[62099] = {9'd98,-10'd302};
ram[62100] = {-9'd99,-10'd299};
ram[62101] = {-9'd96,-10'd296};
ram[62102] = {-9'd92,-10'd293};
ram[62103] = {-9'd89,-10'd290};
ram[62104] = {-9'd86,-10'd286};
ram[62105] = {-9'd83,-10'd283};
ram[62106] = {-9'd80,-10'd280};
ram[62107] = {-9'd77,-10'd277};
ram[62108] = {-9'd74,-10'd274};
ram[62109] = {-9'd70,-10'd271};
ram[62110] = {-9'd67,-10'd268};
ram[62111] = {-9'd64,-10'd264};
ram[62112] = {-9'd61,-10'd261};
ram[62113] = {-9'd58,-10'd258};
ram[62114] = {-9'd55,-10'd255};
ram[62115] = {-9'd52,-10'd252};
ram[62116] = {-9'd48,-10'd249};
ram[62117] = {-9'd45,-10'd246};
ram[62118] = {-9'd42,-10'd242};
ram[62119] = {-9'd39,-10'd239};
ram[62120] = {-9'd36,-10'd236};
ram[62121] = {-9'd33,-10'd233};
ram[62122] = {-9'd30,-10'd230};
ram[62123] = {-9'd26,-10'd227};
ram[62124] = {-9'd23,-10'd224};
ram[62125] = {-9'd20,-10'd220};
ram[62126] = {-9'd17,-10'd217};
ram[62127] = {-9'd14,-10'd214};
ram[62128] = {-9'd11,-10'd211};
ram[62129] = {-9'd8,-10'd208};
ram[62130] = {-9'd4,-10'd205};
ram[62131] = {-9'd1,-10'd202};
ram[62132] = {9'd2,-10'd198};
ram[62133] = {9'd5,-10'd195};
ram[62134] = {9'd8,-10'd192};
ram[62135] = {9'd11,-10'd189};
ram[62136] = {9'd14,-10'd186};
ram[62137] = {9'd18,-10'd183};
ram[62138] = {9'd21,-10'd180};
ram[62139] = {9'd24,-10'd176};
ram[62140] = {9'd27,-10'd173};
ram[62141] = {9'd30,-10'd170};
ram[62142] = {9'd33,-10'd167};
ram[62143] = {9'd36,-10'd164};
ram[62144] = {9'd40,-10'd161};
ram[62145] = {9'd43,-10'd158};
ram[62146] = {9'd46,-10'd154};
ram[62147] = {9'd49,-10'd151};
ram[62148] = {9'd52,-10'd148};
ram[62149] = {9'd55,-10'd145};
ram[62150] = {9'd58,-10'd142};
ram[62151] = {9'd62,-10'd139};
ram[62152] = {9'd65,-10'd136};
ram[62153] = {9'd68,-10'd132};
ram[62154] = {9'd71,-10'd129};
ram[62155] = {9'd74,-10'd126};
ram[62156] = {9'd77,-10'd123};
ram[62157] = {9'd80,-10'd120};
ram[62158] = {9'd84,-10'd117};
ram[62159] = {9'd87,-10'd114};
ram[62160] = {9'd90,-10'd110};
ram[62161] = {9'd93,-10'd107};
ram[62162] = {9'd96,-10'd104};
ram[62163] = {9'd99,-10'd101};
ram[62164] = {-9'd98,-10'd98};
ram[62165] = {-9'd95,-10'd95};
ram[62166] = {-9'd92,-10'd92};
ram[62167] = {-9'd88,-10'd88};
ram[62168] = {-9'd85,-10'd85};
ram[62169] = {-9'd82,-10'd82};
ram[62170] = {-9'd79,-10'd79};
ram[62171] = {-9'd76,-10'd76};
ram[62172] = {-9'd73,-10'd73};
ram[62173] = {-9'd70,-10'd70};
ram[62174] = {-9'd66,-10'd66};
ram[62175] = {-9'd63,-10'd63};
ram[62176] = {-9'd60,-10'd60};
ram[62177] = {-9'd57,-10'd57};
ram[62178] = {-9'd54,-10'd54};
ram[62179] = {-9'd51,-10'd51};
ram[62180] = {-9'd48,-10'd48};
ram[62181] = {-9'd44,-10'd44};
ram[62182] = {-9'd41,-10'd41};
ram[62183] = {-9'd38,-10'd38};
ram[62184] = {-9'd35,-10'd35};
ram[62185] = {-9'd32,-10'd32};
ram[62186] = {-9'd29,-10'd29};
ram[62187] = {-9'd26,-10'd26};
ram[62188] = {-9'd22,-10'd22};
ram[62189] = {-9'd19,-10'd19};
ram[62190] = {-9'd16,-10'd16};
ram[62191] = {-9'd13,-10'd13};
ram[62192] = {-9'd10,-10'd10};
ram[62193] = {-9'd7,-10'd7};
ram[62194] = {-9'd4,-10'd4};
ram[62195] = {9'd0,10'd0};
ram[62196] = {9'd3,10'd3};
ram[62197] = {9'd6,10'd6};
ram[62198] = {9'd9,10'd9};
ram[62199] = {9'd12,10'd12};
ram[62200] = {9'd15,10'd15};
ram[62201] = {9'd18,10'd18};
ram[62202] = {9'd21,10'd21};
ram[62203] = {9'd25,10'd25};
ram[62204] = {9'd28,10'd28};
ram[62205] = {9'd31,10'd31};
ram[62206] = {9'd34,10'd34};
ram[62207] = {9'd37,10'd37};
ram[62208] = {9'd37,10'd37};
ram[62209] = {9'd40,10'd40};
ram[62210] = {9'd43,10'd43};
ram[62211] = {9'd47,10'd47};
ram[62212] = {9'd50,10'd50};
ram[62213] = {9'd53,10'd53};
ram[62214] = {9'd56,10'd56};
ram[62215] = {9'd59,10'd59};
ram[62216] = {9'd62,10'd62};
ram[62217] = {9'd65,10'd65};
ram[62218] = {9'd69,10'd69};
ram[62219] = {9'd72,10'd72};
ram[62220] = {9'd75,10'd75};
ram[62221] = {9'd78,10'd78};
ram[62222] = {9'd81,10'd81};
ram[62223] = {9'd84,10'd84};
ram[62224] = {9'd87,10'd87};
ram[62225] = {9'd91,10'd91};
ram[62226] = {9'd94,10'd94};
ram[62227] = {9'd97,10'd97};
ram[62228] = {-9'd100,10'd100};
ram[62229] = {-9'd97,10'd103};
ram[62230] = {-9'd94,10'd106};
ram[62231] = {-9'd91,10'd109};
ram[62232] = {-9'd88,10'd113};
ram[62233] = {-9'd85,10'd116};
ram[62234] = {-9'd81,10'd119};
ram[62235] = {-9'd78,10'd122};
ram[62236] = {-9'd75,10'd125};
ram[62237] = {-9'd72,10'd128};
ram[62238] = {-9'd69,10'd131};
ram[62239] = {-9'd66,10'd135};
ram[62240] = {-9'd63,10'd138};
ram[62241] = {-9'd59,10'd141};
ram[62242] = {-9'd56,10'd144};
ram[62243] = {-9'd53,10'd147};
ram[62244] = {-9'd50,10'd150};
ram[62245] = {-9'd47,10'd153};
ram[62246] = {-9'd44,10'd157};
ram[62247] = {-9'd41,10'd160};
ram[62248] = {-9'd37,10'd163};
ram[62249] = {-9'd34,10'd166};
ram[62250] = {-9'd31,10'd169};
ram[62251] = {-9'd28,10'd172};
ram[62252] = {-9'd25,10'd175};
ram[62253] = {-9'd22,10'd179};
ram[62254] = {-9'd19,10'd182};
ram[62255] = {-9'd15,10'd185};
ram[62256] = {-9'd12,10'd188};
ram[62257] = {-9'd9,10'd191};
ram[62258] = {-9'd6,10'd194};
ram[62259] = {-9'd3,10'd197};
ram[62260] = {9'd0,10'd201};
ram[62261] = {9'd3,10'd204};
ram[62262] = {9'd7,10'd207};
ram[62263] = {9'd10,10'd210};
ram[62264] = {9'd13,10'd213};
ram[62265] = {9'd16,10'd216};
ram[62266] = {9'd19,10'd219};
ram[62267] = {9'd22,10'd223};
ram[62268] = {9'd25,10'd226};
ram[62269] = {9'd29,10'd229};
ram[62270] = {9'd32,10'd232};
ram[62271] = {9'd35,10'd235};
ram[62272] = {9'd38,10'd238};
ram[62273] = {9'd41,10'd241};
ram[62274] = {9'd44,10'd245};
ram[62275] = {9'd47,10'd248};
ram[62276] = {9'd51,10'd251};
ram[62277] = {9'd54,10'd254};
ram[62278] = {9'd57,10'd257};
ram[62279] = {9'd60,10'd260};
ram[62280] = {9'd63,10'd263};
ram[62281] = {9'd66,10'd267};
ram[62282] = {9'd69,10'd270};
ram[62283] = {9'd73,10'd273};
ram[62284] = {9'd76,10'd276};
ram[62285] = {9'd79,10'd279};
ram[62286] = {9'd82,10'd282};
ram[62287] = {9'd85,10'd285};
ram[62288] = {9'd88,10'd289};
ram[62289] = {9'd91,10'd292};
ram[62290] = {9'd95,10'd295};
ram[62291] = {9'd98,10'd298};
ram[62292] = {-9'd99,10'd301};
ram[62293] = {-9'd96,10'd304};
ram[62294] = {-9'd93,10'd307};
ram[62295] = {-9'd90,10'd311};
ram[62296] = {-9'd87,10'd314};
ram[62297] = {-9'd84,10'd317};
ram[62298] = {-9'd81,10'd320};
ram[62299] = {-9'd77,10'd323};
ram[62300] = {-9'd74,10'd326};
ram[62301] = {-9'd71,10'd329};
ram[62302] = {-9'd68,10'd333};
ram[62303] = {-9'd65,10'd336};
ram[62304] = {-9'd62,10'd339};
ram[62305] = {-9'd59,10'd342};
ram[62306] = {-9'd55,10'd345};
ram[62307] = {-9'd52,10'd348};
ram[62308] = {-9'd49,10'd351};
ram[62309] = {-9'd46,10'd354};
ram[62310] = {-9'd43,10'd358};
ram[62311] = {-9'd40,10'd361};
ram[62312] = {-9'd37,10'd364};
ram[62313] = {-9'd33,10'd367};
ram[62314] = {-9'd30,10'd370};
ram[62315] = {-9'd27,10'd373};
ram[62316] = {-9'd24,10'd376};
ram[62317] = {-9'd21,10'd380};
ram[62318] = {-9'd18,10'd383};
ram[62319] = {-9'd15,10'd386};
ram[62320] = {-9'd11,10'd389};
ram[62321] = {-9'd8,10'd392};
ram[62322] = {-9'd5,10'd395};
ram[62323] = {-9'd2,10'd398};
ram[62324] = {9'd1,-10'd399};
ram[62325] = {9'd4,-10'd396};
ram[62326] = {9'd7,-10'd393};
ram[62327] = {9'd10,-10'd390};
ram[62328] = {9'd14,-10'd387};
ram[62329] = {9'd17,-10'd384};
ram[62330] = {9'd20,-10'd381};
ram[62331] = {9'd23,-10'd377};
ram[62332] = {9'd26,-10'd374};
ram[62333] = {9'd29,-10'd371};
ram[62334] = {9'd32,-10'd368};
ram[62335] = {9'd36,-10'd365};
ram[62336] = {9'd36,-10'd365};
ram[62337] = {9'd39,-10'd362};
ram[62338] = {9'd42,-10'd359};
ram[62339] = {9'd45,-10'd355};
ram[62340] = {9'd48,-10'd352};
ram[62341] = {9'd51,-10'd349};
ram[62342] = {9'd54,-10'd346};
ram[62343] = {9'd58,-10'd343};
ram[62344] = {9'd61,-10'd340};
ram[62345] = {9'd64,-10'd337};
ram[62346] = {9'd67,-10'd334};
ram[62347] = {9'd70,-10'd330};
ram[62348] = {9'd73,-10'd327};
ram[62349] = {9'd76,-10'd324};
ram[62350] = {9'd80,-10'd321};
ram[62351] = {9'd83,-10'd318};
ram[62352] = {9'd86,-10'd315};
ram[62353] = {9'd89,-10'd312};
ram[62354] = {9'd92,-10'd308};
ram[62355] = {9'd95,-10'd305};
ram[62356] = {9'd98,-10'd302};
ram[62357] = {-9'd99,-10'd299};
ram[62358] = {-9'd96,-10'd296};
ram[62359] = {-9'd92,-10'd293};
ram[62360] = {-9'd89,-10'd290};
ram[62361] = {-9'd86,-10'd286};
ram[62362] = {-9'd83,-10'd283};
ram[62363] = {-9'd80,-10'd280};
ram[62364] = {-9'd77,-10'd277};
ram[62365] = {-9'd74,-10'd274};
ram[62366] = {-9'd70,-10'd271};
ram[62367] = {-9'd67,-10'd268};
ram[62368] = {-9'd64,-10'd264};
ram[62369] = {-9'd61,-10'd261};
ram[62370] = {-9'd58,-10'd258};
ram[62371] = {-9'd55,-10'd255};
ram[62372] = {-9'd52,-10'd252};
ram[62373] = {-9'd48,-10'd249};
ram[62374] = {-9'd45,-10'd246};
ram[62375] = {-9'd42,-10'd242};
ram[62376] = {-9'd39,-10'd239};
ram[62377] = {-9'd36,-10'd236};
ram[62378] = {-9'd33,-10'd233};
ram[62379] = {-9'd30,-10'd230};
ram[62380] = {-9'd26,-10'd227};
ram[62381] = {-9'd23,-10'd224};
ram[62382] = {-9'd20,-10'd220};
ram[62383] = {-9'd17,-10'd217};
ram[62384] = {-9'd14,-10'd214};
ram[62385] = {-9'd11,-10'd211};
ram[62386] = {-9'd8,-10'd208};
ram[62387] = {-9'd4,-10'd205};
ram[62388] = {-9'd1,-10'd202};
ram[62389] = {9'd2,-10'd198};
ram[62390] = {9'd5,-10'd195};
ram[62391] = {9'd8,-10'd192};
ram[62392] = {9'd11,-10'd189};
ram[62393] = {9'd14,-10'd186};
ram[62394] = {9'd18,-10'd183};
ram[62395] = {9'd21,-10'd180};
ram[62396] = {9'd24,-10'd176};
ram[62397] = {9'd27,-10'd173};
ram[62398] = {9'd30,-10'd170};
ram[62399] = {9'd33,-10'd167};
ram[62400] = {9'd36,-10'd164};
ram[62401] = {9'd40,-10'd161};
ram[62402] = {9'd43,-10'd158};
ram[62403] = {9'd46,-10'd154};
ram[62404] = {9'd49,-10'd151};
ram[62405] = {9'd52,-10'd148};
ram[62406] = {9'd55,-10'd145};
ram[62407] = {9'd58,-10'd142};
ram[62408] = {9'd62,-10'd139};
ram[62409] = {9'd65,-10'd136};
ram[62410] = {9'd68,-10'd132};
ram[62411] = {9'd71,-10'd129};
ram[62412] = {9'd74,-10'd126};
ram[62413] = {9'd77,-10'd123};
ram[62414] = {9'd80,-10'd120};
ram[62415] = {9'd84,-10'd117};
ram[62416] = {9'd87,-10'd114};
ram[62417] = {9'd90,-10'd110};
ram[62418] = {9'd93,-10'd107};
ram[62419] = {9'd96,-10'd104};
ram[62420] = {9'd99,-10'd101};
ram[62421] = {-9'd98,-10'd98};
ram[62422] = {-9'd95,-10'd95};
ram[62423] = {-9'd92,-10'd92};
ram[62424] = {-9'd88,-10'd88};
ram[62425] = {-9'd85,-10'd85};
ram[62426] = {-9'd82,-10'd82};
ram[62427] = {-9'd79,-10'd79};
ram[62428] = {-9'd76,-10'd76};
ram[62429] = {-9'd73,-10'd73};
ram[62430] = {-9'd70,-10'd70};
ram[62431] = {-9'd66,-10'd66};
ram[62432] = {-9'd63,-10'd63};
ram[62433] = {-9'd60,-10'd60};
ram[62434] = {-9'd57,-10'd57};
ram[62435] = {-9'd54,-10'd54};
ram[62436] = {-9'd51,-10'd51};
ram[62437] = {-9'd48,-10'd48};
ram[62438] = {-9'd44,-10'd44};
ram[62439] = {-9'd41,-10'd41};
ram[62440] = {-9'd38,-10'd38};
ram[62441] = {-9'd35,-10'd35};
ram[62442] = {-9'd32,-10'd32};
ram[62443] = {-9'd29,-10'd29};
ram[62444] = {-9'd26,-10'd26};
ram[62445] = {-9'd22,-10'd22};
ram[62446] = {-9'd19,-10'd19};
ram[62447] = {-9'd16,-10'd16};
ram[62448] = {-9'd13,-10'd13};
ram[62449] = {-9'd10,-10'd10};
ram[62450] = {-9'd7,-10'd7};
ram[62451] = {-9'd4,-10'd4};
ram[62452] = {9'd0,10'd0};
ram[62453] = {9'd3,10'd3};
ram[62454] = {9'd6,10'd6};
ram[62455] = {9'd9,10'd9};
ram[62456] = {9'd12,10'd12};
ram[62457] = {9'd15,10'd15};
ram[62458] = {9'd18,10'd18};
ram[62459] = {9'd21,10'd21};
ram[62460] = {9'd25,10'd25};
ram[62461] = {9'd28,10'd28};
ram[62462] = {9'd31,10'd31};
ram[62463] = {9'd34,10'd34};
ram[62464] = {9'd34,10'd34};
ram[62465] = {9'd37,10'd37};
ram[62466] = {9'd40,10'd40};
ram[62467] = {9'd43,10'd43};
ram[62468] = {9'd47,10'd47};
ram[62469] = {9'd50,10'd50};
ram[62470] = {9'd53,10'd53};
ram[62471] = {9'd56,10'd56};
ram[62472] = {9'd59,10'd59};
ram[62473] = {9'd62,10'd62};
ram[62474] = {9'd65,10'd65};
ram[62475] = {9'd69,10'd69};
ram[62476] = {9'd72,10'd72};
ram[62477] = {9'd75,10'd75};
ram[62478] = {9'd78,10'd78};
ram[62479] = {9'd81,10'd81};
ram[62480] = {9'd84,10'd84};
ram[62481] = {9'd87,10'd87};
ram[62482] = {9'd91,10'd91};
ram[62483] = {9'd94,10'd94};
ram[62484] = {9'd97,10'd97};
ram[62485] = {-9'd100,10'd100};
ram[62486] = {-9'd97,10'd103};
ram[62487] = {-9'd94,10'd106};
ram[62488] = {-9'd91,10'd109};
ram[62489] = {-9'd88,10'd113};
ram[62490] = {-9'd85,10'd116};
ram[62491] = {-9'd81,10'd119};
ram[62492] = {-9'd78,10'd122};
ram[62493] = {-9'd75,10'd125};
ram[62494] = {-9'd72,10'd128};
ram[62495] = {-9'd69,10'd131};
ram[62496] = {-9'd66,10'd135};
ram[62497] = {-9'd63,10'd138};
ram[62498] = {-9'd59,10'd141};
ram[62499] = {-9'd56,10'd144};
ram[62500] = {-9'd53,10'd147};
ram[62501] = {-9'd50,10'd150};
ram[62502] = {-9'd47,10'd153};
ram[62503] = {-9'd44,10'd157};
ram[62504] = {-9'd41,10'd160};
ram[62505] = {-9'd37,10'd163};
ram[62506] = {-9'd34,10'd166};
ram[62507] = {-9'd31,10'd169};
ram[62508] = {-9'd28,10'd172};
ram[62509] = {-9'd25,10'd175};
ram[62510] = {-9'd22,10'd179};
ram[62511] = {-9'd19,10'd182};
ram[62512] = {-9'd15,10'd185};
ram[62513] = {-9'd12,10'd188};
ram[62514] = {-9'd9,10'd191};
ram[62515] = {-9'd6,10'd194};
ram[62516] = {-9'd3,10'd197};
ram[62517] = {9'd0,10'd201};
ram[62518] = {9'd3,10'd204};
ram[62519] = {9'd7,10'd207};
ram[62520] = {9'd10,10'd210};
ram[62521] = {9'd13,10'd213};
ram[62522] = {9'd16,10'd216};
ram[62523] = {9'd19,10'd219};
ram[62524] = {9'd22,10'd223};
ram[62525] = {9'd25,10'd226};
ram[62526] = {9'd29,10'd229};
ram[62527] = {9'd32,10'd232};
ram[62528] = {9'd35,10'd235};
ram[62529] = {9'd38,10'd238};
ram[62530] = {9'd41,10'd241};
ram[62531] = {9'd44,10'd245};
ram[62532] = {9'd47,10'd248};
ram[62533] = {9'd51,10'd251};
ram[62534] = {9'd54,10'd254};
ram[62535] = {9'd57,10'd257};
ram[62536] = {9'd60,10'd260};
ram[62537] = {9'd63,10'd263};
ram[62538] = {9'd66,10'd267};
ram[62539] = {9'd69,10'd270};
ram[62540] = {9'd73,10'd273};
ram[62541] = {9'd76,10'd276};
ram[62542] = {9'd79,10'd279};
ram[62543] = {9'd82,10'd282};
ram[62544] = {9'd85,10'd285};
ram[62545] = {9'd88,10'd289};
ram[62546] = {9'd91,10'd292};
ram[62547] = {9'd95,10'd295};
ram[62548] = {9'd98,10'd298};
ram[62549] = {-9'd99,10'd301};
ram[62550] = {-9'd96,10'd304};
ram[62551] = {-9'd93,10'd307};
ram[62552] = {-9'd90,10'd311};
ram[62553] = {-9'd87,10'd314};
ram[62554] = {-9'd84,10'd317};
ram[62555] = {-9'd81,10'd320};
ram[62556] = {-9'd77,10'd323};
ram[62557] = {-9'd74,10'd326};
ram[62558] = {-9'd71,10'd329};
ram[62559] = {-9'd68,10'd333};
ram[62560] = {-9'd65,10'd336};
ram[62561] = {-9'd62,10'd339};
ram[62562] = {-9'd59,10'd342};
ram[62563] = {-9'd55,10'd345};
ram[62564] = {-9'd52,10'd348};
ram[62565] = {-9'd49,10'd351};
ram[62566] = {-9'd46,10'd354};
ram[62567] = {-9'd43,10'd358};
ram[62568] = {-9'd40,10'd361};
ram[62569] = {-9'd37,10'd364};
ram[62570] = {-9'd33,10'd367};
ram[62571] = {-9'd30,10'd370};
ram[62572] = {-9'd27,10'd373};
ram[62573] = {-9'd24,10'd376};
ram[62574] = {-9'd21,10'd380};
ram[62575] = {-9'd18,10'd383};
ram[62576] = {-9'd15,10'd386};
ram[62577] = {-9'd11,10'd389};
ram[62578] = {-9'd8,10'd392};
ram[62579] = {-9'd5,10'd395};
ram[62580] = {-9'd2,10'd398};
ram[62581] = {9'd1,-10'd399};
ram[62582] = {9'd4,-10'd396};
ram[62583] = {9'd7,-10'd393};
ram[62584] = {9'd10,-10'd390};
ram[62585] = {9'd14,-10'd387};
ram[62586] = {9'd17,-10'd384};
ram[62587] = {9'd20,-10'd381};
ram[62588] = {9'd23,-10'd377};
ram[62589] = {9'd26,-10'd374};
ram[62590] = {9'd29,-10'd371};
ram[62591] = {9'd32,-10'd368};
ram[62592] = {9'd32,-10'd368};
ram[62593] = {9'd36,-10'd365};
ram[62594] = {9'd39,-10'd362};
ram[62595] = {9'd42,-10'd359};
ram[62596] = {9'd45,-10'd355};
ram[62597] = {9'd48,-10'd352};
ram[62598] = {9'd51,-10'd349};
ram[62599] = {9'd54,-10'd346};
ram[62600] = {9'd58,-10'd343};
ram[62601] = {9'd61,-10'd340};
ram[62602] = {9'd64,-10'd337};
ram[62603] = {9'd67,-10'd334};
ram[62604] = {9'd70,-10'd330};
ram[62605] = {9'd73,-10'd327};
ram[62606] = {9'd76,-10'd324};
ram[62607] = {9'd80,-10'd321};
ram[62608] = {9'd83,-10'd318};
ram[62609] = {9'd86,-10'd315};
ram[62610] = {9'd89,-10'd312};
ram[62611] = {9'd92,-10'd308};
ram[62612] = {9'd95,-10'd305};
ram[62613] = {9'd98,-10'd302};
ram[62614] = {-9'd99,-10'd299};
ram[62615] = {-9'd96,-10'd296};
ram[62616] = {-9'd92,-10'd293};
ram[62617] = {-9'd89,-10'd290};
ram[62618] = {-9'd86,-10'd286};
ram[62619] = {-9'd83,-10'd283};
ram[62620] = {-9'd80,-10'd280};
ram[62621] = {-9'd77,-10'd277};
ram[62622] = {-9'd74,-10'd274};
ram[62623] = {-9'd70,-10'd271};
ram[62624] = {-9'd67,-10'd268};
ram[62625] = {-9'd64,-10'd264};
ram[62626] = {-9'd61,-10'd261};
ram[62627] = {-9'd58,-10'd258};
ram[62628] = {-9'd55,-10'd255};
ram[62629] = {-9'd52,-10'd252};
ram[62630] = {-9'd48,-10'd249};
ram[62631] = {-9'd45,-10'd246};
ram[62632] = {-9'd42,-10'd242};
ram[62633] = {-9'd39,-10'd239};
ram[62634] = {-9'd36,-10'd236};
ram[62635] = {-9'd33,-10'd233};
ram[62636] = {-9'd30,-10'd230};
ram[62637] = {-9'd26,-10'd227};
ram[62638] = {-9'd23,-10'd224};
ram[62639] = {-9'd20,-10'd220};
ram[62640] = {-9'd17,-10'd217};
ram[62641] = {-9'd14,-10'd214};
ram[62642] = {-9'd11,-10'd211};
ram[62643] = {-9'd8,-10'd208};
ram[62644] = {-9'd4,-10'd205};
ram[62645] = {-9'd1,-10'd202};
ram[62646] = {9'd2,-10'd198};
ram[62647] = {9'd5,-10'd195};
ram[62648] = {9'd8,-10'd192};
ram[62649] = {9'd11,-10'd189};
ram[62650] = {9'd14,-10'd186};
ram[62651] = {9'd18,-10'd183};
ram[62652] = {9'd21,-10'd180};
ram[62653] = {9'd24,-10'd176};
ram[62654] = {9'd27,-10'd173};
ram[62655] = {9'd30,-10'd170};
ram[62656] = {9'd33,-10'd167};
ram[62657] = {9'd36,-10'd164};
ram[62658] = {9'd40,-10'd161};
ram[62659] = {9'd43,-10'd158};
ram[62660] = {9'd46,-10'd154};
ram[62661] = {9'd49,-10'd151};
ram[62662] = {9'd52,-10'd148};
ram[62663] = {9'd55,-10'd145};
ram[62664] = {9'd58,-10'd142};
ram[62665] = {9'd62,-10'd139};
ram[62666] = {9'd65,-10'd136};
ram[62667] = {9'd68,-10'd132};
ram[62668] = {9'd71,-10'd129};
ram[62669] = {9'd74,-10'd126};
ram[62670] = {9'd77,-10'd123};
ram[62671] = {9'd80,-10'd120};
ram[62672] = {9'd84,-10'd117};
ram[62673] = {9'd87,-10'd114};
ram[62674] = {9'd90,-10'd110};
ram[62675] = {9'd93,-10'd107};
ram[62676] = {9'd96,-10'd104};
ram[62677] = {9'd99,-10'd101};
ram[62678] = {-9'd98,-10'd98};
ram[62679] = {-9'd95,-10'd95};
ram[62680] = {-9'd92,-10'd92};
ram[62681] = {-9'd88,-10'd88};
ram[62682] = {-9'd85,-10'd85};
ram[62683] = {-9'd82,-10'd82};
ram[62684] = {-9'd79,-10'd79};
ram[62685] = {-9'd76,-10'd76};
ram[62686] = {-9'd73,-10'd73};
ram[62687] = {-9'd70,-10'd70};
ram[62688] = {-9'd66,-10'd66};
ram[62689] = {-9'd63,-10'd63};
ram[62690] = {-9'd60,-10'd60};
ram[62691] = {-9'd57,-10'd57};
ram[62692] = {-9'd54,-10'd54};
ram[62693] = {-9'd51,-10'd51};
ram[62694] = {-9'd48,-10'd48};
ram[62695] = {-9'd44,-10'd44};
ram[62696] = {-9'd41,-10'd41};
ram[62697] = {-9'd38,-10'd38};
ram[62698] = {-9'd35,-10'd35};
ram[62699] = {-9'd32,-10'd32};
ram[62700] = {-9'd29,-10'd29};
ram[62701] = {-9'd26,-10'd26};
ram[62702] = {-9'd22,-10'd22};
ram[62703] = {-9'd19,-10'd19};
ram[62704] = {-9'd16,-10'd16};
ram[62705] = {-9'd13,-10'd13};
ram[62706] = {-9'd10,-10'd10};
ram[62707] = {-9'd7,-10'd7};
ram[62708] = {-9'd4,-10'd4};
ram[62709] = {9'd0,10'd0};
ram[62710] = {9'd3,10'd3};
ram[62711] = {9'd6,10'd6};
ram[62712] = {9'd9,10'd9};
ram[62713] = {9'd12,10'd12};
ram[62714] = {9'd15,10'd15};
ram[62715] = {9'd18,10'd18};
ram[62716] = {9'd21,10'd21};
ram[62717] = {9'd25,10'd25};
ram[62718] = {9'd28,10'd28};
ram[62719] = {9'd31,10'd31};
ram[62720] = {9'd31,10'd31};
ram[62721] = {9'd34,10'd34};
ram[62722] = {9'd37,10'd37};
ram[62723] = {9'd40,10'd40};
ram[62724] = {9'd43,10'd43};
ram[62725] = {9'd47,10'd47};
ram[62726] = {9'd50,10'd50};
ram[62727] = {9'd53,10'd53};
ram[62728] = {9'd56,10'd56};
ram[62729] = {9'd59,10'd59};
ram[62730] = {9'd62,10'd62};
ram[62731] = {9'd65,10'd65};
ram[62732] = {9'd69,10'd69};
ram[62733] = {9'd72,10'd72};
ram[62734] = {9'd75,10'd75};
ram[62735] = {9'd78,10'd78};
ram[62736] = {9'd81,10'd81};
ram[62737] = {9'd84,10'd84};
ram[62738] = {9'd87,10'd87};
ram[62739] = {9'd91,10'd91};
ram[62740] = {9'd94,10'd94};
ram[62741] = {9'd97,10'd97};
ram[62742] = {-9'd100,10'd100};
ram[62743] = {-9'd97,10'd103};
ram[62744] = {-9'd94,10'd106};
ram[62745] = {-9'd91,10'd109};
ram[62746] = {-9'd88,10'd113};
ram[62747] = {-9'd85,10'd116};
ram[62748] = {-9'd81,10'd119};
ram[62749] = {-9'd78,10'd122};
ram[62750] = {-9'd75,10'd125};
ram[62751] = {-9'd72,10'd128};
ram[62752] = {-9'd69,10'd131};
ram[62753] = {-9'd66,10'd135};
ram[62754] = {-9'd63,10'd138};
ram[62755] = {-9'd59,10'd141};
ram[62756] = {-9'd56,10'd144};
ram[62757] = {-9'd53,10'd147};
ram[62758] = {-9'd50,10'd150};
ram[62759] = {-9'd47,10'd153};
ram[62760] = {-9'd44,10'd157};
ram[62761] = {-9'd41,10'd160};
ram[62762] = {-9'd37,10'd163};
ram[62763] = {-9'd34,10'd166};
ram[62764] = {-9'd31,10'd169};
ram[62765] = {-9'd28,10'd172};
ram[62766] = {-9'd25,10'd175};
ram[62767] = {-9'd22,10'd179};
ram[62768] = {-9'd19,10'd182};
ram[62769] = {-9'd15,10'd185};
ram[62770] = {-9'd12,10'd188};
ram[62771] = {-9'd9,10'd191};
ram[62772] = {-9'd6,10'd194};
ram[62773] = {-9'd3,10'd197};
ram[62774] = {9'd0,10'd201};
ram[62775] = {9'd3,10'd204};
ram[62776] = {9'd7,10'd207};
ram[62777] = {9'd10,10'd210};
ram[62778] = {9'd13,10'd213};
ram[62779] = {9'd16,10'd216};
ram[62780] = {9'd19,10'd219};
ram[62781] = {9'd22,10'd223};
ram[62782] = {9'd25,10'd226};
ram[62783] = {9'd29,10'd229};
ram[62784] = {9'd32,10'd232};
ram[62785] = {9'd35,10'd235};
ram[62786] = {9'd38,10'd238};
ram[62787] = {9'd41,10'd241};
ram[62788] = {9'd44,10'd245};
ram[62789] = {9'd47,10'd248};
ram[62790] = {9'd51,10'd251};
ram[62791] = {9'd54,10'd254};
ram[62792] = {9'd57,10'd257};
ram[62793] = {9'd60,10'd260};
ram[62794] = {9'd63,10'd263};
ram[62795] = {9'd66,10'd267};
ram[62796] = {9'd69,10'd270};
ram[62797] = {9'd73,10'd273};
ram[62798] = {9'd76,10'd276};
ram[62799] = {9'd79,10'd279};
ram[62800] = {9'd82,10'd282};
ram[62801] = {9'd85,10'd285};
ram[62802] = {9'd88,10'd289};
ram[62803] = {9'd91,10'd292};
ram[62804] = {9'd95,10'd295};
ram[62805] = {9'd98,10'd298};
ram[62806] = {-9'd99,10'd301};
ram[62807] = {-9'd96,10'd304};
ram[62808] = {-9'd93,10'd307};
ram[62809] = {-9'd90,10'd311};
ram[62810] = {-9'd87,10'd314};
ram[62811] = {-9'd84,10'd317};
ram[62812] = {-9'd81,10'd320};
ram[62813] = {-9'd77,10'd323};
ram[62814] = {-9'd74,10'd326};
ram[62815] = {-9'd71,10'd329};
ram[62816] = {-9'd68,10'd333};
ram[62817] = {-9'd65,10'd336};
ram[62818] = {-9'd62,10'd339};
ram[62819] = {-9'd59,10'd342};
ram[62820] = {-9'd55,10'd345};
ram[62821] = {-9'd52,10'd348};
ram[62822] = {-9'd49,10'd351};
ram[62823] = {-9'd46,10'd354};
ram[62824] = {-9'd43,10'd358};
ram[62825] = {-9'd40,10'd361};
ram[62826] = {-9'd37,10'd364};
ram[62827] = {-9'd33,10'd367};
ram[62828] = {-9'd30,10'd370};
ram[62829] = {-9'd27,10'd373};
ram[62830] = {-9'd24,10'd376};
ram[62831] = {-9'd21,10'd380};
ram[62832] = {-9'd18,10'd383};
ram[62833] = {-9'd15,10'd386};
ram[62834] = {-9'd11,10'd389};
ram[62835] = {-9'd8,10'd392};
ram[62836] = {-9'd5,10'd395};
ram[62837] = {-9'd2,10'd398};
ram[62838] = {9'd1,-10'd399};
ram[62839] = {9'd4,-10'd396};
ram[62840] = {9'd7,-10'd393};
ram[62841] = {9'd10,-10'd390};
ram[62842] = {9'd14,-10'd387};
ram[62843] = {9'd17,-10'd384};
ram[62844] = {9'd20,-10'd381};
ram[62845] = {9'd23,-10'd377};
ram[62846] = {9'd26,-10'd374};
ram[62847] = {9'd29,-10'd371};
ram[62848] = {9'd29,-10'd371};
ram[62849] = {9'd32,-10'd368};
ram[62850] = {9'd36,-10'd365};
ram[62851] = {9'd39,-10'd362};
ram[62852] = {9'd42,-10'd359};
ram[62853] = {9'd45,-10'd355};
ram[62854] = {9'd48,-10'd352};
ram[62855] = {9'd51,-10'd349};
ram[62856] = {9'd54,-10'd346};
ram[62857] = {9'd58,-10'd343};
ram[62858] = {9'd61,-10'd340};
ram[62859] = {9'd64,-10'd337};
ram[62860] = {9'd67,-10'd334};
ram[62861] = {9'd70,-10'd330};
ram[62862] = {9'd73,-10'd327};
ram[62863] = {9'd76,-10'd324};
ram[62864] = {9'd80,-10'd321};
ram[62865] = {9'd83,-10'd318};
ram[62866] = {9'd86,-10'd315};
ram[62867] = {9'd89,-10'd312};
ram[62868] = {9'd92,-10'd308};
ram[62869] = {9'd95,-10'd305};
ram[62870] = {9'd98,-10'd302};
ram[62871] = {-9'd99,-10'd299};
ram[62872] = {-9'd96,-10'd296};
ram[62873] = {-9'd92,-10'd293};
ram[62874] = {-9'd89,-10'd290};
ram[62875] = {-9'd86,-10'd286};
ram[62876] = {-9'd83,-10'd283};
ram[62877] = {-9'd80,-10'd280};
ram[62878] = {-9'd77,-10'd277};
ram[62879] = {-9'd74,-10'd274};
ram[62880] = {-9'd70,-10'd271};
ram[62881] = {-9'd67,-10'd268};
ram[62882] = {-9'd64,-10'd264};
ram[62883] = {-9'd61,-10'd261};
ram[62884] = {-9'd58,-10'd258};
ram[62885] = {-9'd55,-10'd255};
ram[62886] = {-9'd52,-10'd252};
ram[62887] = {-9'd48,-10'd249};
ram[62888] = {-9'd45,-10'd246};
ram[62889] = {-9'd42,-10'd242};
ram[62890] = {-9'd39,-10'd239};
ram[62891] = {-9'd36,-10'd236};
ram[62892] = {-9'd33,-10'd233};
ram[62893] = {-9'd30,-10'd230};
ram[62894] = {-9'd26,-10'd227};
ram[62895] = {-9'd23,-10'd224};
ram[62896] = {-9'd20,-10'd220};
ram[62897] = {-9'd17,-10'd217};
ram[62898] = {-9'd14,-10'd214};
ram[62899] = {-9'd11,-10'd211};
ram[62900] = {-9'd8,-10'd208};
ram[62901] = {-9'd4,-10'd205};
ram[62902] = {-9'd1,-10'd202};
ram[62903] = {9'd2,-10'd198};
ram[62904] = {9'd5,-10'd195};
ram[62905] = {9'd8,-10'd192};
ram[62906] = {9'd11,-10'd189};
ram[62907] = {9'd14,-10'd186};
ram[62908] = {9'd18,-10'd183};
ram[62909] = {9'd21,-10'd180};
ram[62910] = {9'd24,-10'd176};
ram[62911] = {9'd27,-10'd173};
ram[62912] = {9'd30,-10'd170};
ram[62913] = {9'd33,-10'd167};
ram[62914] = {9'd36,-10'd164};
ram[62915] = {9'd40,-10'd161};
ram[62916] = {9'd43,-10'd158};
ram[62917] = {9'd46,-10'd154};
ram[62918] = {9'd49,-10'd151};
ram[62919] = {9'd52,-10'd148};
ram[62920] = {9'd55,-10'd145};
ram[62921] = {9'd58,-10'd142};
ram[62922] = {9'd62,-10'd139};
ram[62923] = {9'd65,-10'd136};
ram[62924] = {9'd68,-10'd132};
ram[62925] = {9'd71,-10'd129};
ram[62926] = {9'd74,-10'd126};
ram[62927] = {9'd77,-10'd123};
ram[62928] = {9'd80,-10'd120};
ram[62929] = {9'd84,-10'd117};
ram[62930] = {9'd87,-10'd114};
ram[62931] = {9'd90,-10'd110};
ram[62932] = {9'd93,-10'd107};
ram[62933] = {9'd96,-10'd104};
ram[62934] = {9'd99,-10'd101};
ram[62935] = {-9'd98,-10'd98};
ram[62936] = {-9'd95,-10'd95};
ram[62937] = {-9'd92,-10'd92};
ram[62938] = {-9'd88,-10'd88};
ram[62939] = {-9'd85,-10'd85};
ram[62940] = {-9'd82,-10'd82};
ram[62941] = {-9'd79,-10'd79};
ram[62942] = {-9'd76,-10'd76};
ram[62943] = {-9'd73,-10'd73};
ram[62944] = {-9'd70,-10'd70};
ram[62945] = {-9'd66,-10'd66};
ram[62946] = {-9'd63,-10'd63};
ram[62947] = {-9'd60,-10'd60};
ram[62948] = {-9'd57,-10'd57};
ram[62949] = {-9'd54,-10'd54};
ram[62950] = {-9'd51,-10'd51};
ram[62951] = {-9'd48,-10'd48};
ram[62952] = {-9'd44,-10'd44};
ram[62953] = {-9'd41,-10'd41};
ram[62954] = {-9'd38,-10'd38};
ram[62955] = {-9'd35,-10'd35};
ram[62956] = {-9'd32,-10'd32};
ram[62957] = {-9'd29,-10'd29};
ram[62958] = {-9'd26,-10'd26};
ram[62959] = {-9'd22,-10'd22};
ram[62960] = {-9'd19,-10'd19};
ram[62961] = {-9'd16,-10'd16};
ram[62962] = {-9'd13,-10'd13};
ram[62963] = {-9'd10,-10'd10};
ram[62964] = {-9'd7,-10'd7};
ram[62965] = {-9'd4,-10'd4};
ram[62966] = {9'd0,10'd0};
ram[62967] = {9'd3,10'd3};
ram[62968] = {9'd6,10'd6};
ram[62969] = {9'd9,10'd9};
ram[62970] = {9'd12,10'd12};
ram[62971] = {9'd15,10'd15};
ram[62972] = {9'd18,10'd18};
ram[62973] = {9'd21,10'd21};
ram[62974] = {9'd25,10'd25};
ram[62975] = {9'd28,10'd28};
ram[62976] = {9'd28,10'd28};
ram[62977] = {9'd31,10'd31};
ram[62978] = {9'd34,10'd34};
ram[62979] = {9'd37,10'd37};
ram[62980] = {9'd40,10'd40};
ram[62981] = {9'd43,10'd43};
ram[62982] = {9'd47,10'd47};
ram[62983] = {9'd50,10'd50};
ram[62984] = {9'd53,10'd53};
ram[62985] = {9'd56,10'd56};
ram[62986] = {9'd59,10'd59};
ram[62987] = {9'd62,10'd62};
ram[62988] = {9'd65,10'd65};
ram[62989] = {9'd69,10'd69};
ram[62990] = {9'd72,10'd72};
ram[62991] = {9'd75,10'd75};
ram[62992] = {9'd78,10'd78};
ram[62993] = {9'd81,10'd81};
ram[62994] = {9'd84,10'd84};
ram[62995] = {9'd87,10'd87};
ram[62996] = {9'd91,10'd91};
ram[62997] = {9'd94,10'd94};
ram[62998] = {9'd97,10'd97};
ram[62999] = {-9'd100,10'd100};
ram[63000] = {-9'd97,10'd103};
ram[63001] = {-9'd94,10'd106};
ram[63002] = {-9'd91,10'd109};
ram[63003] = {-9'd88,10'd113};
ram[63004] = {-9'd85,10'd116};
ram[63005] = {-9'd81,10'd119};
ram[63006] = {-9'd78,10'd122};
ram[63007] = {-9'd75,10'd125};
ram[63008] = {-9'd72,10'd128};
ram[63009] = {-9'd69,10'd131};
ram[63010] = {-9'd66,10'd135};
ram[63011] = {-9'd63,10'd138};
ram[63012] = {-9'd59,10'd141};
ram[63013] = {-9'd56,10'd144};
ram[63014] = {-9'd53,10'd147};
ram[63015] = {-9'd50,10'd150};
ram[63016] = {-9'd47,10'd153};
ram[63017] = {-9'd44,10'd157};
ram[63018] = {-9'd41,10'd160};
ram[63019] = {-9'd37,10'd163};
ram[63020] = {-9'd34,10'd166};
ram[63021] = {-9'd31,10'd169};
ram[63022] = {-9'd28,10'd172};
ram[63023] = {-9'd25,10'd175};
ram[63024] = {-9'd22,10'd179};
ram[63025] = {-9'd19,10'd182};
ram[63026] = {-9'd15,10'd185};
ram[63027] = {-9'd12,10'd188};
ram[63028] = {-9'd9,10'd191};
ram[63029] = {-9'd6,10'd194};
ram[63030] = {-9'd3,10'd197};
ram[63031] = {9'd0,10'd201};
ram[63032] = {9'd3,10'd204};
ram[63033] = {9'd7,10'd207};
ram[63034] = {9'd10,10'd210};
ram[63035] = {9'd13,10'd213};
ram[63036] = {9'd16,10'd216};
ram[63037] = {9'd19,10'd219};
ram[63038] = {9'd22,10'd223};
ram[63039] = {9'd25,10'd226};
ram[63040] = {9'd29,10'd229};
ram[63041] = {9'd32,10'd232};
ram[63042] = {9'd35,10'd235};
ram[63043] = {9'd38,10'd238};
ram[63044] = {9'd41,10'd241};
ram[63045] = {9'd44,10'd245};
ram[63046] = {9'd47,10'd248};
ram[63047] = {9'd51,10'd251};
ram[63048] = {9'd54,10'd254};
ram[63049] = {9'd57,10'd257};
ram[63050] = {9'd60,10'd260};
ram[63051] = {9'd63,10'd263};
ram[63052] = {9'd66,10'd267};
ram[63053] = {9'd69,10'd270};
ram[63054] = {9'd73,10'd273};
ram[63055] = {9'd76,10'd276};
ram[63056] = {9'd79,10'd279};
ram[63057] = {9'd82,10'd282};
ram[63058] = {9'd85,10'd285};
ram[63059] = {9'd88,10'd289};
ram[63060] = {9'd91,10'd292};
ram[63061] = {9'd95,10'd295};
ram[63062] = {9'd98,10'd298};
ram[63063] = {-9'd99,10'd301};
ram[63064] = {-9'd96,10'd304};
ram[63065] = {-9'd93,10'd307};
ram[63066] = {-9'd90,10'd311};
ram[63067] = {-9'd87,10'd314};
ram[63068] = {-9'd84,10'd317};
ram[63069] = {-9'd81,10'd320};
ram[63070] = {-9'd77,10'd323};
ram[63071] = {-9'd74,10'd326};
ram[63072] = {-9'd71,10'd329};
ram[63073] = {-9'd68,10'd333};
ram[63074] = {-9'd65,10'd336};
ram[63075] = {-9'd62,10'd339};
ram[63076] = {-9'd59,10'd342};
ram[63077] = {-9'd55,10'd345};
ram[63078] = {-9'd52,10'd348};
ram[63079] = {-9'd49,10'd351};
ram[63080] = {-9'd46,10'd354};
ram[63081] = {-9'd43,10'd358};
ram[63082] = {-9'd40,10'd361};
ram[63083] = {-9'd37,10'd364};
ram[63084] = {-9'd33,10'd367};
ram[63085] = {-9'd30,10'd370};
ram[63086] = {-9'd27,10'd373};
ram[63087] = {-9'd24,10'd376};
ram[63088] = {-9'd21,10'd380};
ram[63089] = {-9'd18,10'd383};
ram[63090] = {-9'd15,10'd386};
ram[63091] = {-9'd11,10'd389};
ram[63092] = {-9'd8,10'd392};
ram[63093] = {-9'd5,10'd395};
ram[63094] = {-9'd2,10'd398};
ram[63095] = {9'd1,-10'd399};
ram[63096] = {9'd4,-10'd396};
ram[63097] = {9'd7,-10'd393};
ram[63098] = {9'd10,-10'd390};
ram[63099] = {9'd14,-10'd387};
ram[63100] = {9'd17,-10'd384};
ram[63101] = {9'd20,-10'd381};
ram[63102] = {9'd23,-10'd377};
ram[63103] = {9'd26,-10'd374};
ram[63104] = {9'd26,-10'd374};
ram[63105] = {9'd29,-10'd371};
ram[63106] = {9'd32,-10'd368};
ram[63107] = {9'd36,-10'd365};
ram[63108] = {9'd39,-10'd362};
ram[63109] = {9'd42,-10'd359};
ram[63110] = {9'd45,-10'd355};
ram[63111] = {9'd48,-10'd352};
ram[63112] = {9'd51,-10'd349};
ram[63113] = {9'd54,-10'd346};
ram[63114] = {9'd58,-10'd343};
ram[63115] = {9'd61,-10'd340};
ram[63116] = {9'd64,-10'd337};
ram[63117] = {9'd67,-10'd334};
ram[63118] = {9'd70,-10'd330};
ram[63119] = {9'd73,-10'd327};
ram[63120] = {9'd76,-10'd324};
ram[63121] = {9'd80,-10'd321};
ram[63122] = {9'd83,-10'd318};
ram[63123] = {9'd86,-10'd315};
ram[63124] = {9'd89,-10'd312};
ram[63125] = {9'd92,-10'd308};
ram[63126] = {9'd95,-10'd305};
ram[63127] = {9'd98,-10'd302};
ram[63128] = {-9'd99,-10'd299};
ram[63129] = {-9'd96,-10'd296};
ram[63130] = {-9'd92,-10'd293};
ram[63131] = {-9'd89,-10'd290};
ram[63132] = {-9'd86,-10'd286};
ram[63133] = {-9'd83,-10'd283};
ram[63134] = {-9'd80,-10'd280};
ram[63135] = {-9'd77,-10'd277};
ram[63136] = {-9'd74,-10'd274};
ram[63137] = {-9'd70,-10'd271};
ram[63138] = {-9'd67,-10'd268};
ram[63139] = {-9'd64,-10'd264};
ram[63140] = {-9'd61,-10'd261};
ram[63141] = {-9'd58,-10'd258};
ram[63142] = {-9'd55,-10'd255};
ram[63143] = {-9'd52,-10'd252};
ram[63144] = {-9'd48,-10'd249};
ram[63145] = {-9'd45,-10'd246};
ram[63146] = {-9'd42,-10'd242};
ram[63147] = {-9'd39,-10'd239};
ram[63148] = {-9'd36,-10'd236};
ram[63149] = {-9'd33,-10'd233};
ram[63150] = {-9'd30,-10'd230};
ram[63151] = {-9'd26,-10'd227};
ram[63152] = {-9'd23,-10'd224};
ram[63153] = {-9'd20,-10'd220};
ram[63154] = {-9'd17,-10'd217};
ram[63155] = {-9'd14,-10'd214};
ram[63156] = {-9'd11,-10'd211};
ram[63157] = {-9'd8,-10'd208};
ram[63158] = {-9'd4,-10'd205};
ram[63159] = {-9'd1,-10'd202};
ram[63160] = {9'd2,-10'd198};
ram[63161] = {9'd5,-10'd195};
ram[63162] = {9'd8,-10'd192};
ram[63163] = {9'd11,-10'd189};
ram[63164] = {9'd14,-10'd186};
ram[63165] = {9'd18,-10'd183};
ram[63166] = {9'd21,-10'd180};
ram[63167] = {9'd24,-10'd176};
ram[63168] = {9'd27,-10'd173};
ram[63169] = {9'd30,-10'd170};
ram[63170] = {9'd33,-10'd167};
ram[63171] = {9'd36,-10'd164};
ram[63172] = {9'd40,-10'd161};
ram[63173] = {9'd43,-10'd158};
ram[63174] = {9'd46,-10'd154};
ram[63175] = {9'd49,-10'd151};
ram[63176] = {9'd52,-10'd148};
ram[63177] = {9'd55,-10'd145};
ram[63178] = {9'd58,-10'd142};
ram[63179] = {9'd62,-10'd139};
ram[63180] = {9'd65,-10'd136};
ram[63181] = {9'd68,-10'd132};
ram[63182] = {9'd71,-10'd129};
ram[63183] = {9'd74,-10'd126};
ram[63184] = {9'd77,-10'd123};
ram[63185] = {9'd80,-10'd120};
ram[63186] = {9'd84,-10'd117};
ram[63187] = {9'd87,-10'd114};
ram[63188] = {9'd90,-10'd110};
ram[63189] = {9'd93,-10'd107};
ram[63190] = {9'd96,-10'd104};
ram[63191] = {9'd99,-10'd101};
ram[63192] = {-9'd98,-10'd98};
ram[63193] = {-9'd95,-10'd95};
ram[63194] = {-9'd92,-10'd92};
ram[63195] = {-9'd88,-10'd88};
ram[63196] = {-9'd85,-10'd85};
ram[63197] = {-9'd82,-10'd82};
ram[63198] = {-9'd79,-10'd79};
ram[63199] = {-9'd76,-10'd76};
ram[63200] = {-9'd73,-10'd73};
ram[63201] = {-9'd70,-10'd70};
ram[63202] = {-9'd66,-10'd66};
ram[63203] = {-9'd63,-10'd63};
ram[63204] = {-9'd60,-10'd60};
ram[63205] = {-9'd57,-10'd57};
ram[63206] = {-9'd54,-10'd54};
ram[63207] = {-9'd51,-10'd51};
ram[63208] = {-9'd48,-10'd48};
ram[63209] = {-9'd44,-10'd44};
ram[63210] = {-9'd41,-10'd41};
ram[63211] = {-9'd38,-10'd38};
ram[63212] = {-9'd35,-10'd35};
ram[63213] = {-9'd32,-10'd32};
ram[63214] = {-9'd29,-10'd29};
ram[63215] = {-9'd26,-10'd26};
ram[63216] = {-9'd22,-10'd22};
ram[63217] = {-9'd19,-10'd19};
ram[63218] = {-9'd16,-10'd16};
ram[63219] = {-9'd13,-10'd13};
ram[63220] = {-9'd10,-10'd10};
ram[63221] = {-9'd7,-10'd7};
ram[63222] = {-9'd4,-10'd4};
ram[63223] = {9'd0,10'd0};
ram[63224] = {9'd3,10'd3};
ram[63225] = {9'd6,10'd6};
ram[63226] = {9'd9,10'd9};
ram[63227] = {9'd12,10'd12};
ram[63228] = {9'd15,10'd15};
ram[63229] = {9'd18,10'd18};
ram[63230] = {9'd21,10'd21};
ram[63231] = {9'd25,10'd25};
ram[63232] = {9'd25,10'd25};
ram[63233] = {9'd28,10'd28};
ram[63234] = {9'd31,10'd31};
ram[63235] = {9'd34,10'd34};
ram[63236] = {9'd37,10'd37};
ram[63237] = {9'd40,10'd40};
ram[63238] = {9'd43,10'd43};
ram[63239] = {9'd47,10'd47};
ram[63240] = {9'd50,10'd50};
ram[63241] = {9'd53,10'd53};
ram[63242] = {9'd56,10'd56};
ram[63243] = {9'd59,10'd59};
ram[63244] = {9'd62,10'd62};
ram[63245] = {9'd65,10'd65};
ram[63246] = {9'd69,10'd69};
ram[63247] = {9'd72,10'd72};
ram[63248] = {9'd75,10'd75};
ram[63249] = {9'd78,10'd78};
ram[63250] = {9'd81,10'd81};
ram[63251] = {9'd84,10'd84};
ram[63252] = {9'd87,10'd87};
ram[63253] = {9'd91,10'd91};
ram[63254] = {9'd94,10'd94};
ram[63255] = {9'd97,10'd97};
ram[63256] = {-9'd100,10'd100};
ram[63257] = {-9'd97,10'd103};
ram[63258] = {-9'd94,10'd106};
ram[63259] = {-9'd91,10'd109};
ram[63260] = {-9'd88,10'd113};
ram[63261] = {-9'd85,10'd116};
ram[63262] = {-9'd81,10'd119};
ram[63263] = {-9'd78,10'd122};
ram[63264] = {-9'd75,10'd125};
ram[63265] = {-9'd72,10'd128};
ram[63266] = {-9'd69,10'd131};
ram[63267] = {-9'd66,10'd135};
ram[63268] = {-9'd63,10'd138};
ram[63269] = {-9'd59,10'd141};
ram[63270] = {-9'd56,10'd144};
ram[63271] = {-9'd53,10'd147};
ram[63272] = {-9'd50,10'd150};
ram[63273] = {-9'd47,10'd153};
ram[63274] = {-9'd44,10'd157};
ram[63275] = {-9'd41,10'd160};
ram[63276] = {-9'd37,10'd163};
ram[63277] = {-9'd34,10'd166};
ram[63278] = {-9'd31,10'd169};
ram[63279] = {-9'd28,10'd172};
ram[63280] = {-9'd25,10'd175};
ram[63281] = {-9'd22,10'd179};
ram[63282] = {-9'd19,10'd182};
ram[63283] = {-9'd15,10'd185};
ram[63284] = {-9'd12,10'd188};
ram[63285] = {-9'd9,10'd191};
ram[63286] = {-9'd6,10'd194};
ram[63287] = {-9'd3,10'd197};
ram[63288] = {9'd0,10'd201};
ram[63289] = {9'd3,10'd204};
ram[63290] = {9'd7,10'd207};
ram[63291] = {9'd10,10'd210};
ram[63292] = {9'd13,10'd213};
ram[63293] = {9'd16,10'd216};
ram[63294] = {9'd19,10'd219};
ram[63295] = {9'd22,10'd223};
ram[63296] = {9'd25,10'd226};
ram[63297] = {9'd29,10'd229};
ram[63298] = {9'd32,10'd232};
ram[63299] = {9'd35,10'd235};
ram[63300] = {9'd38,10'd238};
ram[63301] = {9'd41,10'd241};
ram[63302] = {9'd44,10'd245};
ram[63303] = {9'd47,10'd248};
ram[63304] = {9'd51,10'd251};
ram[63305] = {9'd54,10'd254};
ram[63306] = {9'd57,10'd257};
ram[63307] = {9'd60,10'd260};
ram[63308] = {9'd63,10'd263};
ram[63309] = {9'd66,10'd267};
ram[63310] = {9'd69,10'd270};
ram[63311] = {9'd73,10'd273};
ram[63312] = {9'd76,10'd276};
ram[63313] = {9'd79,10'd279};
ram[63314] = {9'd82,10'd282};
ram[63315] = {9'd85,10'd285};
ram[63316] = {9'd88,10'd289};
ram[63317] = {9'd91,10'd292};
ram[63318] = {9'd95,10'd295};
ram[63319] = {9'd98,10'd298};
ram[63320] = {-9'd99,10'd301};
ram[63321] = {-9'd96,10'd304};
ram[63322] = {-9'd93,10'd307};
ram[63323] = {-9'd90,10'd311};
ram[63324] = {-9'd87,10'd314};
ram[63325] = {-9'd84,10'd317};
ram[63326] = {-9'd81,10'd320};
ram[63327] = {-9'd77,10'd323};
ram[63328] = {-9'd74,10'd326};
ram[63329] = {-9'd71,10'd329};
ram[63330] = {-9'd68,10'd333};
ram[63331] = {-9'd65,10'd336};
ram[63332] = {-9'd62,10'd339};
ram[63333] = {-9'd59,10'd342};
ram[63334] = {-9'd55,10'd345};
ram[63335] = {-9'd52,10'd348};
ram[63336] = {-9'd49,10'd351};
ram[63337] = {-9'd46,10'd354};
ram[63338] = {-9'd43,10'd358};
ram[63339] = {-9'd40,10'd361};
ram[63340] = {-9'd37,10'd364};
ram[63341] = {-9'd33,10'd367};
ram[63342] = {-9'd30,10'd370};
ram[63343] = {-9'd27,10'd373};
ram[63344] = {-9'd24,10'd376};
ram[63345] = {-9'd21,10'd380};
ram[63346] = {-9'd18,10'd383};
ram[63347] = {-9'd15,10'd386};
ram[63348] = {-9'd11,10'd389};
ram[63349] = {-9'd8,10'd392};
ram[63350] = {-9'd5,10'd395};
ram[63351] = {-9'd2,10'd398};
ram[63352] = {9'd1,-10'd399};
ram[63353] = {9'd4,-10'd396};
ram[63354] = {9'd7,-10'd393};
ram[63355] = {9'd10,-10'd390};
ram[63356] = {9'd14,-10'd387};
ram[63357] = {9'd17,-10'd384};
ram[63358] = {9'd20,-10'd381};
ram[63359] = {9'd23,-10'd377};
ram[63360] = {9'd23,-10'd377};
ram[63361] = {9'd26,-10'd374};
ram[63362] = {9'd29,-10'd371};
ram[63363] = {9'd32,-10'd368};
ram[63364] = {9'd36,-10'd365};
ram[63365] = {9'd39,-10'd362};
ram[63366] = {9'd42,-10'd359};
ram[63367] = {9'd45,-10'd355};
ram[63368] = {9'd48,-10'd352};
ram[63369] = {9'd51,-10'd349};
ram[63370] = {9'd54,-10'd346};
ram[63371] = {9'd58,-10'd343};
ram[63372] = {9'd61,-10'd340};
ram[63373] = {9'd64,-10'd337};
ram[63374] = {9'd67,-10'd334};
ram[63375] = {9'd70,-10'd330};
ram[63376] = {9'd73,-10'd327};
ram[63377] = {9'd76,-10'd324};
ram[63378] = {9'd80,-10'd321};
ram[63379] = {9'd83,-10'd318};
ram[63380] = {9'd86,-10'd315};
ram[63381] = {9'd89,-10'd312};
ram[63382] = {9'd92,-10'd308};
ram[63383] = {9'd95,-10'd305};
ram[63384] = {9'd98,-10'd302};
ram[63385] = {-9'd99,-10'd299};
ram[63386] = {-9'd96,-10'd296};
ram[63387] = {-9'd92,-10'd293};
ram[63388] = {-9'd89,-10'd290};
ram[63389] = {-9'd86,-10'd286};
ram[63390] = {-9'd83,-10'd283};
ram[63391] = {-9'd80,-10'd280};
ram[63392] = {-9'd77,-10'd277};
ram[63393] = {-9'd74,-10'd274};
ram[63394] = {-9'd70,-10'd271};
ram[63395] = {-9'd67,-10'd268};
ram[63396] = {-9'd64,-10'd264};
ram[63397] = {-9'd61,-10'd261};
ram[63398] = {-9'd58,-10'd258};
ram[63399] = {-9'd55,-10'd255};
ram[63400] = {-9'd52,-10'd252};
ram[63401] = {-9'd48,-10'd249};
ram[63402] = {-9'd45,-10'd246};
ram[63403] = {-9'd42,-10'd242};
ram[63404] = {-9'd39,-10'd239};
ram[63405] = {-9'd36,-10'd236};
ram[63406] = {-9'd33,-10'd233};
ram[63407] = {-9'd30,-10'd230};
ram[63408] = {-9'd26,-10'd227};
ram[63409] = {-9'd23,-10'd224};
ram[63410] = {-9'd20,-10'd220};
ram[63411] = {-9'd17,-10'd217};
ram[63412] = {-9'd14,-10'd214};
ram[63413] = {-9'd11,-10'd211};
ram[63414] = {-9'd8,-10'd208};
ram[63415] = {-9'd4,-10'd205};
ram[63416] = {-9'd1,-10'd202};
ram[63417] = {9'd2,-10'd198};
ram[63418] = {9'd5,-10'd195};
ram[63419] = {9'd8,-10'd192};
ram[63420] = {9'd11,-10'd189};
ram[63421] = {9'd14,-10'd186};
ram[63422] = {9'd18,-10'd183};
ram[63423] = {9'd21,-10'd180};
ram[63424] = {9'd24,-10'd176};
ram[63425] = {9'd27,-10'd173};
ram[63426] = {9'd30,-10'd170};
ram[63427] = {9'd33,-10'd167};
ram[63428] = {9'd36,-10'd164};
ram[63429] = {9'd40,-10'd161};
ram[63430] = {9'd43,-10'd158};
ram[63431] = {9'd46,-10'd154};
ram[63432] = {9'd49,-10'd151};
ram[63433] = {9'd52,-10'd148};
ram[63434] = {9'd55,-10'd145};
ram[63435] = {9'd58,-10'd142};
ram[63436] = {9'd62,-10'd139};
ram[63437] = {9'd65,-10'd136};
ram[63438] = {9'd68,-10'd132};
ram[63439] = {9'd71,-10'd129};
ram[63440] = {9'd74,-10'd126};
ram[63441] = {9'd77,-10'd123};
ram[63442] = {9'd80,-10'd120};
ram[63443] = {9'd84,-10'd117};
ram[63444] = {9'd87,-10'd114};
ram[63445] = {9'd90,-10'd110};
ram[63446] = {9'd93,-10'd107};
ram[63447] = {9'd96,-10'd104};
ram[63448] = {9'd99,-10'd101};
ram[63449] = {-9'd98,-10'd98};
ram[63450] = {-9'd95,-10'd95};
ram[63451] = {-9'd92,-10'd92};
ram[63452] = {-9'd88,-10'd88};
ram[63453] = {-9'd85,-10'd85};
ram[63454] = {-9'd82,-10'd82};
ram[63455] = {-9'd79,-10'd79};
ram[63456] = {-9'd76,-10'd76};
ram[63457] = {-9'd73,-10'd73};
ram[63458] = {-9'd70,-10'd70};
ram[63459] = {-9'd66,-10'd66};
ram[63460] = {-9'd63,-10'd63};
ram[63461] = {-9'd60,-10'd60};
ram[63462] = {-9'd57,-10'd57};
ram[63463] = {-9'd54,-10'd54};
ram[63464] = {-9'd51,-10'd51};
ram[63465] = {-9'd48,-10'd48};
ram[63466] = {-9'd44,-10'd44};
ram[63467] = {-9'd41,-10'd41};
ram[63468] = {-9'd38,-10'd38};
ram[63469] = {-9'd35,-10'd35};
ram[63470] = {-9'd32,-10'd32};
ram[63471] = {-9'd29,-10'd29};
ram[63472] = {-9'd26,-10'd26};
ram[63473] = {-9'd22,-10'd22};
ram[63474] = {-9'd19,-10'd19};
ram[63475] = {-9'd16,-10'd16};
ram[63476] = {-9'd13,-10'd13};
ram[63477] = {-9'd10,-10'd10};
ram[63478] = {-9'd7,-10'd7};
ram[63479] = {-9'd4,-10'd4};
ram[63480] = {9'd0,10'd0};
ram[63481] = {9'd3,10'd3};
ram[63482] = {9'd6,10'd6};
ram[63483] = {9'd9,10'd9};
ram[63484] = {9'd12,10'd12};
ram[63485] = {9'd15,10'd15};
ram[63486] = {9'd18,10'd18};
ram[63487] = {9'd21,10'd21};
ram[63488] = {9'd21,10'd21};
ram[63489] = {9'd25,10'd25};
ram[63490] = {9'd28,10'd28};
ram[63491] = {9'd31,10'd31};
ram[63492] = {9'd34,10'd34};
ram[63493] = {9'd37,10'd37};
ram[63494] = {9'd40,10'd40};
ram[63495] = {9'd43,10'd43};
ram[63496] = {9'd47,10'd47};
ram[63497] = {9'd50,10'd50};
ram[63498] = {9'd53,10'd53};
ram[63499] = {9'd56,10'd56};
ram[63500] = {9'd59,10'd59};
ram[63501] = {9'd62,10'd62};
ram[63502] = {9'd65,10'd65};
ram[63503] = {9'd69,10'd69};
ram[63504] = {9'd72,10'd72};
ram[63505] = {9'd75,10'd75};
ram[63506] = {9'd78,10'd78};
ram[63507] = {9'd81,10'd81};
ram[63508] = {9'd84,10'd84};
ram[63509] = {9'd87,10'd87};
ram[63510] = {9'd91,10'd91};
ram[63511] = {9'd94,10'd94};
ram[63512] = {9'd97,10'd97};
ram[63513] = {-9'd100,10'd100};
ram[63514] = {-9'd97,10'd103};
ram[63515] = {-9'd94,10'd106};
ram[63516] = {-9'd91,10'd109};
ram[63517] = {-9'd88,10'd113};
ram[63518] = {-9'd85,10'd116};
ram[63519] = {-9'd81,10'd119};
ram[63520] = {-9'd78,10'd122};
ram[63521] = {-9'd75,10'd125};
ram[63522] = {-9'd72,10'd128};
ram[63523] = {-9'd69,10'd131};
ram[63524] = {-9'd66,10'd135};
ram[63525] = {-9'd63,10'd138};
ram[63526] = {-9'd59,10'd141};
ram[63527] = {-9'd56,10'd144};
ram[63528] = {-9'd53,10'd147};
ram[63529] = {-9'd50,10'd150};
ram[63530] = {-9'd47,10'd153};
ram[63531] = {-9'd44,10'd157};
ram[63532] = {-9'd41,10'd160};
ram[63533] = {-9'd37,10'd163};
ram[63534] = {-9'd34,10'd166};
ram[63535] = {-9'd31,10'd169};
ram[63536] = {-9'd28,10'd172};
ram[63537] = {-9'd25,10'd175};
ram[63538] = {-9'd22,10'd179};
ram[63539] = {-9'd19,10'd182};
ram[63540] = {-9'd15,10'd185};
ram[63541] = {-9'd12,10'd188};
ram[63542] = {-9'd9,10'd191};
ram[63543] = {-9'd6,10'd194};
ram[63544] = {-9'd3,10'd197};
ram[63545] = {9'd0,10'd201};
ram[63546] = {9'd3,10'd204};
ram[63547] = {9'd7,10'd207};
ram[63548] = {9'd10,10'd210};
ram[63549] = {9'd13,10'd213};
ram[63550] = {9'd16,10'd216};
ram[63551] = {9'd19,10'd219};
ram[63552] = {9'd22,10'd223};
ram[63553] = {9'd25,10'd226};
ram[63554] = {9'd29,10'd229};
ram[63555] = {9'd32,10'd232};
ram[63556] = {9'd35,10'd235};
ram[63557] = {9'd38,10'd238};
ram[63558] = {9'd41,10'd241};
ram[63559] = {9'd44,10'd245};
ram[63560] = {9'd47,10'd248};
ram[63561] = {9'd51,10'd251};
ram[63562] = {9'd54,10'd254};
ram[63563] = {9'd57,10'd257};
ram[63564] = {9'd60,10'd260};
ram[63565] = {9'd63,10'd263};
ram[63566] = {9'd66,10'd267};
ram[63567] = {9'd69,10'd270};
ram[63568] = {9'd73,10'd273};
ram[63569] = {9'd76,10'd276};
ram[63570] = {9'd79,10'd279};
ram[63571] = {9'd82,10'd282};
ram[63572] = {9'd85,10'd285};
ram[63573] = {9'd88,10'd289};
ram[63574] = {9'd91,10'd292};
ram[63575] = {9'd95,10'd295};
ram[63576] = {9'd98,10'd298};
ram[63577] = {-9'd99,10'd301};
ram[63578] = {-9'd96,10'd304};
ram[63579] = {-9'd93,10'd307};
ram[63580] = {-9'd90,10'd311};
ram[63581] = {-9'd87,10'd314};
ram[63582] = {-9'd84,10'd317};
ram[63583] = {-9'd81,10'd320};
ram[63584] = {-9'd77,10'd323};
ram[63585] = {-9'd74,10'd326};
ram[63586] = {-9'd71,10'd329};
ram[63587] = {-9'd68,10'd333};
ram[63588] = {-9'd65,10'd336};
ram[63589] = {-9'd62,10'd339};
ram[63590] = {-9'd59,10'd342};
ram[63591] = {-9'd55,10'd345};
ram[63592] = {-9'd52,10'd348};
ram[63593] = {-9'd49,10'd351};
ram[63594] = {-9'd46,10'd354};
ram[63595] = {-9'd43,10'd358};
ram[63596] = {-9'd40,10'd361};
ram[63597] = {-9'd37,10'd364};
ram[63598] = {-9'd33,10'd367};
ram[63599] = {-9'd30,10'd370};
ram[63600] = {-9'd27,10'd373};
ram[63601] = {-9'd24,10'd376};
ram[63602] = {-9'd21,10'd380};
ram[63603] = {-9'd18,10'd383};
ram[63604] = {-9'd15,10'd386};
ram[63605] = {-9'd11,10'd389};
ram[63606] = {-9'd8,10'd392};
ram[63607] = {-9'd5,10'd395};
ram[63608] = {-9'd2,10'd398};
ram[63609] = {9'd1,-10'd399};
ram[63610] = {9'd4,-10'd396};
ram[63611] = {9'd7,-10'd393};
ram[63612] = {9'd10,-10'd390};
ram[63613] = {9'd14,-10'd387};
ram[63614] = {9'd17,-10'd384};
ram[63615] = {9'd20,-10'd381};
ram[63616] = {9'd20,-10'd381};
ram[63617] = {9'd23,-10'd377};
ram[63618] = {9'd26,-10'd374};
ram[63619] = {9'd29,-10'd371};
ram[63620] = {9'd32,-10'd368};
ram[63621] = {9'd36,-10'd365};
ram[63622] = {9'd39,-10'd362};
ram[63623] = {9'd42,-10'd359};
ram[63624] = {9'd45,-10'd355};
ram[63625] = {9'd48,-10'd352};
ram[63626] = {9'd51,-10'd349};
ram[63627] = {9'd54,-10'd346};
ram[63628] = {9'd58,-10'd343};
ram[63629] = {9'd61,-10'd340};
ram[63630] = {9'd64,-10'd337};
ram[63631] = {9'd67,-10'd334};
ram[63632] = {9'd70,-10'd330};
ram[63633] = {9'd73,-10'd327};
ram[63634] = {9'd76,-10'd324};
ram[63635] = {9'd80,-10'd321};
ram[63636] = {9'd83,-10'd318};
ram[63637] = {9'd86,-10'd315};
ram[63638] = {9'd89,-10'd312};
ram[63639] = {9'd92,-10'd308};
ram[63640] = {9'd95,-10'd305};
ram[63641] = {9'd98,-10'd302};
ram[63642] = {-9'd99,-10'd299};
ram[63643] = {-9'd96,-10'd296};
ram[63644] = {-9'd92,-10'd293};
ram[63645] = {-9'd89,-10'd290};
ram[63646] = {-9'd86,-10'd286};
ram[63647] = {-9'd83,-10'd283};
ram[63648] = {-9'd80,-10'd280};
ram[63649] = {-9'd77,-10'd277};
ram[63650] = {-9'd74,-10'd274};
ram[63651] = {-9'd70,-10'd271};
ram[63652] = {-9'd67,-10'd268};
ram[63653] = {-9'd64,-10'd264};
ram[63654] = {-9'd61,-10'd261};
ram[63655] = {-9'd58,-10'd258};
ram[63656] = {-9'd55,-10'd255};
ram[63657] = {-9'd52,-10'd252};
ram[63658] = {-9'd48,-10'd249};
ram[63659] = {-9'd45,-10'd246};
ram[63660] = {-9'd42,-10'd242};
ram[63661] = {-9'd39,-10'd239};
ram[63662] = {-9'd36,-10'd236};
ram[63663] = {-9'd33,-10'd233};
ram[63664] = {-9'd30,-10'd230};
ram[63665] = {-9'd26,-10'd227};
ram[63666] = {-9'd23,-10'd224};
ram[63667] = {-9'd20,-10'd220};
ram[63668] = {-9'd17,-10'd217};
ram[63669] = {-9'd14,-10'd214};
ram[63670] = {-9'd11,-10'd211};
ram[63671] = {-9'd8,-10'd208};
ram[63672] = {-9'd4,-10'd205};
ram[63673] = {-9'd1,-10'd202};
ram[63674] = {9'd2,-10'd198};
ram[63675] = {9'd5,-10'd195};
ram[63676] = {9'd8,-10'd192};
ram[63677] = {9'd11,-10'd189};
ram[63678] = {9'd14,-10'd186};
ram[63679] = {9'd18,-10'd183};
ram[63680] = {9'd21,-10'd180};
ram[63681] = {9'd24,-10'd176};
ram[63682] = {9'd27,-10'd173};
ram[63683] = {9'd30,-10'd170};
ram[63684] = {9'd33,-10'd167};
ram[63685] = {9'd36,-10'd164};
ram[63686] = {9'd40,-10'd161};
ram[63687] = {9'd43,-10'd158};
ram[63688] = {9'd46,-10'd154};
ram[63689] = {9'd49,-10'd151};
ram[63690] = {9'd52,-10'd148};
ram[63691] = {9'd55,-10'd145};
ram[63692] = {9'd58,-10'd142};
ram[63693] = {9'd62,-10'd139};
ram[63694] = {9'd65,-10'd136};
ram[63695] = {9'd68,-10'd132};
ram[63696] = {9'd71,-10'd129};
ram[63697] = {9'd74,-10'd126};
ram[63698] = {9'd77,-10'd123};
ram[63699] = {9'd80,-10'd120};
ram[63700] = {9'd84,-10'd117};
ram[63701] = {9'd87,-10'd114};
ram[63702] = {9'd90,-10'd110};
ram[63703] = {9'd93,-10'd107};
ram[63704] = {9'd96,-10'd104};
ram[63705] = {9'd99,-10'd101};
ram[63706] = {-9'd98,-10'd98};
ram[63707] = {-9'd95,-10'd95};
ram[63708] = {-9'd92,-10'd92};
ram[63709] = {-9'd88,-10'd88};
ram[63710] = {-9'd85,-10'd85};
ram[63711] = {-9'd82,-10'd82};
ram[63712] = {-9'd79,-10'd79};
ram[63713] = {-9'd76,-10'd76};
ram[63714] = {-9'd73,-10'd73};
ram[63715] = {-9'd70,-10'd70};
ram[63716] = {-9'd66,-10'd66};
ram[63717] = {-9'd63,-10'd63};
ram[63718] = {-9'd60,-10'd60};
ram[63719] = {-9'd57,-10'd57};
ram[63720] = {-9'd54,-10'd54};
ram[63721] = {-9'd51,-10'd51};
ram[63722] = {-9'd48,-10'd48};
ram[63723] = {-9'd44,-10'd44};
ram[63724] = {-9'd41,-10'd41};
ram[63725] = {-9'd38,-10'd38};
ram[63726] = {-9'd35,-10'd35};
ram[63727] = {-9'd32,-10'd32};
ram[63728] = {-9'd29,-10'd29};
ram[63729] = {-9'd26,-10'd26};
ram[63730] = {-9'd22,-10'd22};
ram[63731] = {-9'd19,-10'd19};
ram[63732] = {-9'd16,-10'd16};
ram[63733] = {-9'd13,-10'd13};
ram[63734] = {-9'd10,-10'd10};
ram[63735] = {-9'd7,-10'd7};
ram[63736] = {-9'd4,-10'd4};
ram[63737] = {9'd0,10'd0};
ram[63738] = {9'd3,10'd3};
ram[63739] = {9'd6,10'd6};
ram[63740] = {9'd9,10'd9};
ram[63741] = {9'd12,10'd12};
ram[63742] = {9'd15,10'd15};
ram[63743] = {9'd18,10'd18};
ram[63744] = {9'd18,10'd18};
ram[63745] = {9'd21,10'd21};
ram[63746] = {9'd25,10'd25};
ram[63747] = {9'd28,10'd28};
ram[63748] = {9'd31,10'd31};
ram[63749] = {9'd34,10'd34};
ram[63750] = {9'd37,10'd37};
ram[63751] = {9'd40,10'd40};
ram[63752] = {9'd43,10'd43};
ram[63753] = {9'd47,10'd47};
ram[63754] = {9'd50,10'd50};
ram[63755] = {9'd53,10'd53};
ram[63756] = {9'd56,10'd56};
ram[63757] = {9'd59,10'd59};
ram[63758] = {9'd62,10'd62};
ram[63759] = {9'd65,10'd65};
ram[63760] = {9'd69,10'd69};
ram[63761] = {9'd72,10'd72};
ram[63762] = {9'd75,10'd75};
ram[63763] = {9'd78,10'd78};
ram[63764] = {9'd81,10'd81};
ram[63765] = {9'd84,10'd84};
ram[63766] = {9'd87,10'd87};
ram[63767] = {9'd91,10'd91};
ram[63768] = {9'd94,10'd94};
ram[63769] = {9'd97,10'd97};
ram[63770] = {-9'd100,10'd100};
ram[63771] = {-9'd97,10'd103};
ram[63772] = {-9'd94,10'd106};
ram[63773] = {-9'd91,10'd109};
ram[63774] = {-9'd88,10'd113};
ram[63775] = {-9'd85,10'd116};
ram[63776] = {-9'd81,10'd119};
ram[63777] = {-9'd78,10'd122};
ram[63778] = {-9'd75,10'd125};
ram[63779] = {-9'd72,10'd128};
ram[63780] = {-9'd69,10'd131};
ram[63781] = {-9'd66,10'd135};
ram[63782] = {-9'd63,10'd138};
ram[63783] = {-9'd59,10'd141};
ram[63784] = {-9'd56,10'd144};
ram[63785] = {-9'd53,10'd147};
ram[63786] = {-9'd50,10'd150};
ram[63787] = {-9'd47,10'd153};
ram[63788] = {-9'd44,10'd157};
ram[63789] = {-9'd41,10'd160};
ram[63790] = {-9'd37,10'd163};
ram[63791] = {-9'd34,10'd166};
ram[63792] = {-9'd31,10'd169};
ram[63793] = {-9'd28,10'd172};
ram[63794] = {-9'd25,10'd175};
ram[63795] = {-9'd22,10'd179};
ram[63796] = {-9'd19,10'd182};
ram[63797] = {-9'd15,10'd185};
ram[63798] = {-9'd12,10'd188};
ram[63799] = {-9'd9,10'd191};
ram[63800] = {-9'd6,10'd194};
ram[63801] = {-9'd3,10'd197};
ram[63802] = {9'd0,10'd201};
ram[63803] = {9'd3,10'd204};
ram[63804] = {9'd7,10'd207};
ram[63805] = {9'd10,10'd210};
ram[63806] = {9'd13,10'd213};
ram[63807] = {9'd16,10'd216};
ram[63808] = {9'd19,10'd219};
ram[63809] = {9'd22,10'd223};
ram[63810] = {9'd25,10'd226};
ram[63811] = {9'd29,10'd229};
ram[63812] = {9'd32,10'd232};
ram[63813] = {9'd35,10'd235};
ram[63814] = {9'd38,10'd238};
ram[63815] = {9'd41,10'd241};
ram[63816] = {9'd44,10'd245};
ram[63817] = {9'd47,10'd248};
ram[63818] = {9'd51,10'd251};
ram[63819] = {9'd54,10'd254};
ram[63820] = {9'd57,10'd257};
ram[63821] = {9'd60,10'd260};
ram[63822] = {9'd63,10'd263};
ram[63823] = {9'd66,10'd267};
ram[63824] = {9'd69,10'd270};
ram[63825] = {9'd73,10'd273};
ram[63826] = {9'd76,10'd276};
ram[63827] = {9'd79,10'd279};
ram[63828] = {9'd82,10'd282};
ram[63829] = {9'd85,10'd285};
ram[63830] = {9'd88,10'd289};
ram[63831] = {9'd91,10'd292};
ram[63832] = {9'd95,10'd295};
ram[63833] = {9'd98,10'd298};
ram[63834] = {-9'd99,10'd301};
ram[63835] = {-9'd96,10'd304};
ram[63836] = {-9'd93,10'd307};
ram[63837] = {-9'd90,10'd311};
ram[63838] = {-9'd87,10'd314};
ram[63839] = {-9'd84,10'd317};
ram[63840] = {-9'd81,10'd320};
ram[63841] = {-9'd77,10'd323};
ram[63842] = {-9'd74,10'd326};
ram[63843] = {-9'd71,10'd329};
ram[63844] = {-9'd68,10'd333};
ram[63845] = {-9'd65,10'd336};
ram[63846] = {-9'd62,10'd339};
ram[63847] = {-9'd59,10'd342};
ram[63848] = {-9'd55,10'd345};
ram[63849] = {-9'd52,10'd348};
ram[63850] = {-9'd49,10'd351};
ram[63851] = {-9'd46,10'd354};
ram[63852] = {-9'd43,10'd358};
ram[63853] = {-9'd40,10'd361};
ram[63854] = {-9'd37,10'd364};
ram[63855] = {-9'd33,10'd367};
ram[63856] = {-9'd30,10'd370};
ram[63857] = {-9'd27,10'd373};
ram[63858] = {-9'd24,10'd376};
ram[63859] = {-9'd21,10'd380};
ram[63860] = {-9'd18,10'd383};
ram[63861] = {-9'd15,10'd386};
ram[63862] = {-9'd11,10'd389};
ram[63863] = {-9'd8,10'd392};
ram[63864] = {-9'd5,10'd395};
ram[63865] = {-9'd2,10'd398};
ram[63866] = {9'd1,-10'd399};
ram[63867] = {9'd4,-10'd396};
ram[63868] = {9'd7,-10'd393};
ram[63869] = {9'd10,-10'd390};
ram[63870] = {9'd14,-10'd387};
ram[63871] = {9'd17,-10'd384};
ram[63872] = {9'd17,-10'd384};
ram[63873] = {9'd20,-10'd381};
ram[63874] = {9'd23,-10'd377};
ram[63875] = {9'd26,-10'd374};
ram[63876] = {9'd29,-10'd371};
ram[63877] = {9'd32,-10'd368};
ram[63878] = {9'd36,-10'd365};
ram[63879] = {9'd39,-10'd362};
ram[63880] = {9'd42,-10'd359};
ram[63881] = {9'd45,-10'd355};
ram[63882] = {9'd48,-10'd352};
ram[63883] = {9'd51,-10'd349};
ram[63884] = {9'd54,-10'd346};
ram[63885] = {9'd58,-10'd343};
ram[63886] = {9'd61,-10'd340};
ram[63887] = {9'd64,-10'd337};
ram[63888] = {9'd67,-10'd334};
ram[63889] = {9'd70,-10'd330};
ram[63890] = {9'd73,-10'd327};
ram[63891] = {9'd76,-10'd324};
ram[63892] = {9'd80,-10'd321};
ram[63893] = {9'd83,-10'd318};
ram[63894] = {9'd86,-10'd315};
ram[63895] = {9'd89,-10'd312};
ram[63896] = {9'd92,-10'd308};
ram[63897] = {9'd95,-10'd305};
ram[63898] = {9'd98,-10'd302};
ram[63899] = {-9'd99,-10'd299};
ram[63900] = {-9'd96,-10'd296};
ram[63901] = {-9'd92,-10'd293};
ram[63902] = {-9'd89,-10'd290};
ram[63903] = {-9'd86,-10'd286};
ram[63904] = {-9'd83,-10'd283};
ram[63905] = {-9'd80,-10'd280};
ram[63906] = {-9'd77,-10'd277};
ram[63907] = {-9'd74,-10'd274};
ram[63908] = {-9'd70,-10'd271};
ram[63909] = {-9'd67,-10'd268};
ram[63910] = {-9'd64,-10'd264};
ram[63911] = {-9'd61,-10'd261};
ram[63912] = {-9'd58,-10'd258};
ram[63913] = {-9'd55,-10'd255};
ram[63914] = {-9'd52,-10'd252};
ram[63915] = {-9'd48,-10'd249};
ram[63916] = {-9'd45,-10'd246};
ram[63917] = {-9'd42,-10'd242};
ram[63918] = {-9'd39,-10'd239};
ram[63919] = {-9'd36,-10'd236};
ram[63920] = {-9'd33,-10'd233};
ram[63921] = {-9'd30,-10'd230};
ram[63922] = {-9'd26,-10'd227};
ram[63923] = {-9'd23,-10'd224};
ram[63924] = {-9'd20,-10'd220};
ram[63925] = {-9'd17,-10'd217};
ram[63926] = {-9'd14,-10'd214};
ram[63927] = {-9'd11,-10'd211};
ram[63928] = {-9'd8,-10'd208};
ram[63929] = {-9'd4,-10'd205};
ram[63930] = {-9'd1,-10'd202};
ram[63931] = {9'd2,-10'd198};
ram[63932] = {9'd5,-10'd195};
ram[63933] = {9'd8,-10'd192};
ram[63934] = {9'd11,-10'd189};
ram[63935] = {9'd14,-10'd186};
ram[63936] = {9'd18,-10'd183};
ram[63937] = {9'd21,-10'd180};
ram[63938] = {9'd24,-10'd176};
ram[63939] = {9'd27,-10'd173};
ram[63940] = {9'd30,-10'd170};
ram[63941] = {9'd33,-10'd167};
ram[63942] = {9'd36,-10'd164};
ram[63943] = {9'd40,-10'd161};
ram[63944] = {9'd43,-10'd158};
ram[63945] = {9'd46,-10'd154};
ram[63946] = {9'd49,-10'd151};
ram[63947] = {9'd52,-10'd148};
ram[63948] = {9'd55,-10'd145};
ram[63949] = {9'd58,-10'd142};
ram[63950] = {9'd62,-10'd139};
ram[63951] = {9'd65,-10'd136};
ram[63952] = {9'd68,-10'd132};
ram[63953] = {9'd71,-10'd129};
ram[63954] = {9'd74,-10'd126};
ram[63955] = {9'd77,-10'd123};
ram[63956] = {9'd80,-10'd120};
ram[63957] = {9'd84,-10'd117};
ram[63958] = {9'd87,-10'd114};
ram[63959] = {9'd90,-10'd110};
ram[63960] = {9'd93,-10'd107};
ram[63961] = {9'd96,-10'd104};
ram[63962] = {9'd99,-10'd101};
ram[63963] = {-9'd98,-10'd98};
ram[63964] = {-9'd95,-10'd95};
ram[63965] = {-9'd92,-10'd92};
ram[63966] = {-9'd88,-10'd88};
ram[63967] = {-9'd85,-10'd85};
ram[63968] = {-9'd82,-10'd82};
ram[63969] = {-9'd79,-10'd79};
ram[63970] = {-9'd76,-10'd76};
ram[63971] = {-9'd73,-10'd73};
ram[63972] = {-9'd70,-10'd70};
ram[63973] = {-9'd66,-10'd66};
ram[63974] = {-9'd63,-10'd63};
ram[63975] = {-9'd60,-10'd60};
ram[63976] = {-9'd57,-10'd57};
ram[63977] = {-9'd54,-10'd54};
ram[63978] = {-9'd51,-10'd51};
ram[63979] = {-9'd48,-10'd48};
ram[63980] = {-9'd44,-10'd44};
ram[63981] = {-9'd41,-10'd41};
ram[63982] = {-9'd38,-10'd38};
ram[63983] = {-9'd35,-10'd35};
ram[63984] = {-9'd32,-10'd32};
ram[63985] = {-9'd29,-10'd29};
ram[63986] = {-9'd26,-10'd26};
ram[63987] = {-9'd22,-10'd22};
ram[63988] = {-9'd19,-10'd19};
ram[63989] = {-9'd16,-10'd16};
ram[63990] = {-9'd13,-10'd13};
ram[63991] = {-9'd10,-10'd10};
ram[63992] = {-9'd7,-10'd7};
ram[63993] = {-9'd4,-10'd4};
ram[63994] = {9'd0,10'd0};
ram[63995] = {9'd3,10'd3};
ram[63996] = {9'd6,10'd6};
ram[63997] = {9'd9,10'd9};
ram[63998] = {9'd12,10'd12};
ram[63999] = {9'd15,10'd15};
ram[64000] = {9'd15,10'd15};
ram[64001] = {9'd18,10'd18};
ram[64002] = {9'd21,10'd21};
ram[64003] = {9'd25,10'd25};
ram[64004] = {9'd28,10'd28};
ram[64005] = {9'd31,10'd31};
ram[64006] = {9'd34,10'd34};
ram[64007] = {9'd37,10'd37};
ram[64008] = {9'd40,10'd40};
ram[64009] = {9'd43,10'd43};
ram[64010] = {9'd47,10'd47};
ram[64011] = {9'd50,10'd50};
ram[64012] = {9'd53,10'd53};
ram[64013] = {9'd56,10'd56};
ram[64014] = {9'd59,10'd59};
ram[64015] = {9'd62,10'd62};
ram[64016] = {9'd65,10'd65};
ram[64017] = {9'd69,10'd69};
ram[64018] = {9'd72,10'd72};
ram[64019] = {9'd75,10'd75};
ram[64020] = {9'd78,10'd78};
ram[64021] = {9'd81,10'd81};
ram[64022] = {9'd84,10'd84};
ram[64023] = {9'd87,10'd87};
ram[64024] = {9'd91,10'd91};
ram[64025] = {9'd94,10'd94};
ram[64026] = {9'd97,10'd97};
ram[64027] = {-9'd100,10'd100};
ram[64028] = {-9'd97,10'd103};
ram[64029] = {-9'd94,10'd106};
ram[64030] = {-9'd91,10'd109};
ram[64031] = {-9'd88,10'd113};
ram[64032] = {-9'd85,10'd116};
ram[64033] = {-9'd81,10'd119};
ram[64034] = {-9'd78,10'd122};
ram[64035] = {-9'd75,10'd125};
ram[64036] = {-9'd72,10'd128};
ram[64037] = {-9'd69,10'd131};
ram[64038] = {-9'd66,10'd135};
ram[64039] = {-9'd63,10'd138};
ram[64040] = {-9'd59,10'd141};
ram[64041] = {-9'd56,10'd144};
ram[64042] = {-9'd53,10'd147};
ram[64043] = {-9'd50,10'd150};
ram[64044] = {-9'd47,10'd153};
ram[64045] = {-9'd44,10'd157};
ram[64046] = {-9'd41,10'd160};
ram[64047] = {-9'd37,10'd163};
ram[64048] = {-9'd34,10'd166};
ram[64049] = {-9'd31,10'd169};
ram[64050] = {-9'd28,10'd172};
ram[64051] = {-9'd25,10'd175};
ram[64052] = {-9'd22,10'd179};
ram[64053] = {-9'd19,10'd182};
ram[64054] = {-9'd15,10'd185};
ram[64055] = {-9'd12,10'd188};
ram[64056] = {-9'd9,10'd191};
ram[64057] = {-9'd6,10'd194};
ram[64058] = {-9'd3,10'd197};
ram[64059] = {9'd0,10'd201};
ram[64060] = {9'd3,10'd204};
ram[64061] = {9'd7,10'd207};
ram[64062] = {9'd10,10'd210};
ram[64063] = {9'd13,10'd213};
ram[64064] = {9'd16,10'd216};
ram[64065] = {9'd19,10'd219};
ram[64066] = {9'd22,10'd223};
ram[64067] = {9'd25,10'd226};
ram[64068] = {9'd29,10'd229};
ram[64069] = {9'd32,10'd232};
ram[64070] = {9'd35,10'd235};
ram[64071] = {9'd38,10'd238};
ram[64072] = {9'd41,10'd241};
ram[64073] = {9'd44,10'd245};
ram[64074] = {9'd47,10'd248};
ram[64075] = {9'd51,10'd251};
ram[64076] = {9'd54,10'd254};
ram[64077] = {9'd57,10'd257};
ram[64078] = {9'd60,10'd260};
ram[64079] = {9'd63,10'd263};
ram[64080] = {9'd66,10'd267};
ram[64081] = {9'd69,10'd270};
ram[64082] = {9'd73,10'd273};
ram[64083] = {9'd76,10'd276};
ram[64084] = {9'd79,10'd279};
ram[64085] = {9'd82,10'd282};
ram[64086] = {9'd85,10'd285};
ram[64087] = {9'd88,10'd289};
ram[64088] = {9'd91,10'd292};
ram[64089] = {9'd95,10'd295};
ram[64090] = {9'd98,10'd298};
ram[64091] = {-9'd99,10'd301};
ram[64092] = {-9'd96,10'd304};
ram[64093] = {-9'd93,10'd307};
ram[64094] = {-9'd90,10'd311};
ram[64095] = {-9'd87,10'd314};
ram[64096] = {-9'd84,10'd317};
ram[64097] = {-9'd81,10'd320};
ram[64098] = {-9'd77,10'd323};
ram[64099] = {-9'd74,10'd326};
ram[64100] = {-9'd71,10'd329};
ram[64101] = {-9'd68,10'd333};
ram[64102] = {-9'd65,10'd336};
ram[64103] = {-9'd62,10'd339};
ram[64104] = {-9'd59,10'd342};
ram[64105] = {-9'd55,10'd345};
ram[64106] = {-9'd52,10'd348};
ram[64107] = {-9'd49,10'd351};
ram[64108] = {-9'd46,10'd354};
ram[64109] = {-9'd43,10'd358};
ram[64110] = {-9'd40,10'd361};
ram[64111] = {-9'd37,10'd364};
ram[64112] = {-9'd33,10'd367};
ram[64113] = {-9'd30,10'd370};
ram[64114] = {-9'd27,10'd373};
ram[64115] = {-9'd24,10'd376};
ram[64116] = {-9'd21,10'd380};
ram[64117] = {-9'd18,10'd383};
ram[64118] = {-9'd15,10'd386};
ram[64119] = {-9'd11,10'd389};
ram[64120] = {-9'd8,10'd392};
ram[64121] = {-9'd5,10'd395};
ram[64122] = {-9'd2,10'd398};
ram[64123] = {9'd1,-10'd399};
ram[64124] = {9'd4,-10'd396};
ram[64125] = {9'd7,-10'd393};
ram[64126] = {9'd10,-10'd390};
ram[64127] = {9'd14,-10'd387};
ram[64128] = {9'd14,-10'd387};
ram[64129] = {9'd17,-10'd384};
ram[64130] = {9'd20,-10'd381};
ram[64131] = {9'd23,-10'd377};
ram[64132] = {9'd26,-10'd374};
ram[64133] = {9'd29,-10'd371};
ram[64134] = {9'd32,-10'd368};
ram[64135] = {9'd36,-10'd365};
ram[64136] = {9'd39,-10'd362};
ram[64137] = {9'd42,-10'd359};
ram[64138] = {9'd45,-10'd355};
ram[64139] = {9'd48,-10'd352};
ram[64140] = {9'd51,-10'd349};
ram[64141] = {9'd54,-10'd346};
ram[64142] = {9'd58,-10'd343};
ram[64143] = {9'd61,-10'd340};
ram[64144] = {9'd64,-10'd337};
ram[64145] = {9'd67,-10'd334};
ram[64146] = {9'd70,-10'd330};
ram[64147] = {9'd73,-10'd327};
ram[64148] = {9'd76,-10'd324};
ram[64149] = {9'd80,-10'd321};
ram[64150] = {9'd83,-10'd318};
ram[64151] = {9'd86,-10'd315};
ram[64152] = {9'd89,-10'd312};
ram[64153] = {9'd92,-10'd308};
ram[64154] = {9'd95,-10'd305};
ram[64155] = {9'd98,-10'd302};
ram[64156] = {-9'd99,-10'd299};
ram[64157] = {-9'd96,-10'd296};
ram[64158] = {-9'd92,-10'd293};
ram[64159] = {-9'd89,-10'd290};
ram[64160] = {-9'd86,-10'd286};
ram[64161] = {-9'd83,-10'd283};
ram[64162] = {-9'd80,-10'd280};
ram[64163] = {-9'd77,-10'd277};
ram[64164] = {-9'd74,-10'd274};
ram[64165] = {-9'd70,-10'd271};
ram[64166] = {-9'd67,-10'd268};
ram[64167] = {-9'd64,-10'd264};
ram[64168] = {-9'd61,-10'd261};
ram[64169] = {-9'd58,-10'd258};
ram[64170] = {-9'd55,-10'd255};
ram[64171] = {-9'd52,-10'd252};
ram[64172] = {-9'd48,-10'd249};
ram[64173] = {-9'd45,-10'd246};
ram[64174] = {-9'd42,-10'd242};
ram[64175] = {-9'd39,-10'd239};
ram[64176] = {-9'd36,-10'd236};
ram[64177] = {-9'd33,-10'd233};
ram[64178] = {-9'd30,-10'd230};
ram[64179] = {-9'd26,-10'd227};
ram[64180] = {-9'd23,-10'd224};
ram[64181] = {-9'd20,-10'd220};
ram[64182] = {-9'd17,-10'd217};
ram[64183] = {-9'd14,-10'd214};
ram[64184] = {-9'd11,-10'd211};
ram[64185] = {-9'd8,-10'd208};
ram[64186] = {-9'd4,-10'd205};
ram[64187] = {-9'd1,-10'd202};
ram[64188] = {9'd2,-10'd198};
ram[64189] = {9'd5,-10'd195};
ram[64190] = {9'd8,-10'd192};
ram[64191] = {9'd11,-10'd189};
ram[64192] = {9'd14,-10'd186};
ram[64193] = {9'd18,-10'd183};
ram[64194] = {9'd21,-10'd180};
ram[64195] = {9'd24,-10'd176};
ram[64196] = {9'd27,-10'd173};
ram[64197] = {9'd30,-10'd170};
ram[64198] = {9'd33,-10'd167};
ram[64199] = {9'd36,-10'd164};
ram[64200] = {9'd40,-10'd161};
ram[64201] = {9'd43,-10'd158};
ram[64202] = {9'd46,-10'd154};
ram[64203] = {9'd49,-10'd151};
ram[64204] = {9'd52,-10'd148};
ram[64205] = {9'd55,-10'd145};
ram[64206] = {9'd58,-10'd142};
ram[64207] = {9'd62,-10'd139};
ram[64208] = {9'd65,-10'd136};
ram[64209] = {9'd68,-10'd132};
ram[64210] = {9'd71,-10'd129};
ram[64211] = {9'd74,-10'd126};
ram[64212] = {9'd77,-10'd123};
ram[64213] = {9'd80,-10'd120};
ram[64214] = {9'd84,-10'd117};
ram[64215] = {9'd87,-10'd114};
ram[64216] = {9'd90,-10'd110};
ram[64217] = {9'd93,-10'd107};
ram[64218] = {9'd96,-10'd104};
ram[64219] = {9'd99,-10'd101};
ram[64220] = {-9'd98,-10'd98};
ram[64221] = {-9'd95,-10'd95};
ram[64222] = {-9'd92,-10'd92};
ram[64223] = {-9'd88,-10'd88};
ram[64224] = {-9'd85,-10'd85};
ram[64225] = {-9'd82,-10'd82};
ram[64226] = {-9'd79,-10'd79};
ram[64227] = {-9'd76,-10'd76};
ram[64228] = {-9'd73,-10'd73};
ram[64229] = {-9'd70,-10'd70};
ram[64230] = {-9'd66,-10'd66};
ram[64231] = {-9'd63,-10'd63};
ram[64232] = {-9'd60,-10'd60};
ram[64233] = {-9'd57,-10'd57};
ram[64234] = {-9'd54,-10'd54};
ram[64235] = {-9'd51,-10'd51};
ram[64236] = {-9'd48,-10'd48};
ram[64237] = {-9'd44,-10'd44};
ram[64238] = {-9'd41,-10'd41};
ram[64239] = {-9'd38,-10'd38};
ram[64240] = {-9'd35,-10'd35};
ram[64241] = {-9'd32,-10'd32};
ram[64242] = {-9'd29,-10'd29};
ram[64243] = {-9'd26,-10'd26};
ram[64244] = {-9'd22,-10'd22};
ram[64245] = {-9'd19,-10'd19};
ram[64246] = {-9'd16,-10'd16};
ram[64247] = {-9'd13,-10'd13};
ram[64248] = {-9'd10,-10'd10};
ram[64249] = {-9'd7,-10'd7};
ram[64250] = {-9'd4,-10'd4};
ram[64251] = {9'd0,10'd0};
ram[64252] = {9'd3,10'd3};
ram[64253] = {9'd6,10'd6};
ram[64254] = {9'd9,10'd9};
ram[64255] = {9'd12,10'd12};
ram[64256] = {9'd12,10'd12};
ram[64257] = {9'd15,10'd15};
ram[64258] = {9'd18,10'd18};
ram[64259] = {9'd21,10'd21};
ram[64260] = {9'd25,10'd25};
ram[64261] = {9'd28,10'd28};
ram[64262] = {9'd31,10'd31};
ram[64263] = {9'd34,10'd34};
ram[64264] = {9'd37,10'd37};
ram[64265] = {9'd40,10'd40};
ram[64266] = {9'd43,10'd43};
ram[64267] = {9'd47,10'd47};
ram[64268] = {9'd50,10'd50};
ram[64269] = {9'd53,10'd53};
ram[64270] = {9'd56,10'd56};
ram[64271] = {9'd59,10'd59};
ram[64272] = {9'd62,10'd62};
ram[64273] = {9'd65,10'd65};
ram[64274] = {9'd69,10'd69};
ram[64275] = {9'd72,10'd72};
ram[64276] = {9'd75,10'd75};
ram[64277] = {9'd78,10'd78};
ram[64278] = {9'd81,10'd81};
ram[64279] = {9'd84,10'd84};
ram[64280] = {9'd87,10'd87};
ram[64281] = {9'd91,10'd91};
ram[64282] = {9'd94,10'd94};
ram[64283] = {9'd97,10'd97};
ram[64284] = {-9'd100,10'd100};
ram[64285] = {-9'd97,10'd103};
ram[64286] = {-9'd94,10'd106};
ram[64287] = {-9'd91,10'd109};
ram[64288] = {-9'd88,10'd113};
ram[64289] = {-9'd85,10'd116};
ram[64290] = {-9'd81,10'd119};
ram[64291] = {-9'd78,10'd122};
ram[64292] = {-9'd75,10'd125};
ram[64293] = {-9'd72,10'd128};
ram[64294] = {-9'd69,10'd131};
ram[64295] = {-9'd66,10'd135};
ram[64296] = {-9'd63,10'd138};
ram[64297] = {-9'd59,10'd141};
ram[64298] = {-9'd56,10'd144};
ram[64299] = {-9'd53,10'd147};
ram[64300] = {-9'd50,10'd150};
ram[64301] = {-9'd47,10'd153};
ram[64302] = {-9'd44,10'd157};
ram[64303] = {-9'd41,10'd160};
ram[64304] = {-9'd37,10'd163};
ram[64305] = {-9'd34,10'd166};
ram[64306] = {-9'd31,10'd169};
ram[64307] = {-9'd28,10'd172};
ram[64308] = {-9'd25,10'd175};
ram[64309] = {-9'd22,10'd179};
ram[64310] = {-9'd19,10'd182};
ram[64311] = {-9'd15,10'd185};
ram[64312] = {-9'd12,10'd188};
ram[64313] = {-9'd9,10'd191};
ram[64314] = {-9'd6,10'd194};
ram[64315] = {-9'd3,10'd197};
ram[64316] = {9'd0,10'd201};
ram[64317] = {9'd3,10'd204};
ram[64318] = {9'd7,10'd207};
ram[64319] = {9'd10,10'd210};
ram[64320] = {9'd13,10'd213};
ram[64321] = {9'd16,10'd216};
ram[64322] = {9'd19,10'd219};
ram[64323] = {9'd22,10'd223};
ram[64324] = {9'd25,10'd226};
ram[64325] = {9'd29,10'd229};
ram[64326] = {9'd32,10'd232};
ram[64327] = {9'd35,10'd235};
ram[64328] = {9'd38,10'd238};
ram[64329] = {9'd41,10'd241};
ram[64330] = {9'd44,10'd245};
ram[64331] = {9'd47,10'd248};
ram[64332] = {9'd51,10'd251};
ram[64333] = {9'd54,10'd254};
ram[64334] = {9'd57,10'd257};
ram[64335] = {9'd60,10'd260};
ram[64336] = {9'd63,10'd263};
ram[64337] = {9'd66,10'd267};
ram[64338] = {9'd69,10'd270};
ram[64339] = {9'd73,10'd273};
ram[64340] = {9'd76,10'd276};
ram[64341] = {9'd79,10'd279};
ram[64342] = {9'd82,10'd282};
ram[64343] = {9'd85,10'd285};
ram[64344] = {9'd88,10'd289};
ram[64345] = {9'd91,10'd292};
ram[64346] = {9'd95,10'd295};
ram[64347] = {9'd98,10'd298};
ram[64348] = {-9'd99,10'd301};
ram[64349] = {-9'd96,10'd304};
ram[64350] = {-9'd93,10'd307};
ram[64351] = {-9'd90,10'd311};
ram[64352] = {-9'd87,10'd314};
ram[64353] = {-9'd84,10'd317};
ram[64354] = {-9'd81,10'd320};
ram[64355] = {-9'd77,10'd323};
ram[64356] = {-9'd74,10'd326};
ram[64357] = {-9'd71,10'd329};
ram[64358] = {-9'd68,10'd333};
ram[64359] = {-9'd65,10'd336};
ram[64360] = {-9'd62,10'd339};
ram[64361] = {-9'd59,10'd342};
ram[64362] = {-9'd55,10'd345};
ram[64363] = {-9'd52,10'd348};
ram[64364] = {-9'd49,10'd351};
ram[64365] = {-9'd46,10'd354};
ram[64366] = {-9'd43,10'd358};
ram[64367] = {-9'd40,10'd361};
ram[64368] = {-9'd37,10'd364};
ram[64369] = {-9'd33,10'd367};
ram[64370] = {-9'd30,10'd370};
ram[64371] = {-9'd27,10'd373};
ram[64372] = {-9'd24,10'd376};
ram[64373] = {-9'd21,10'd380};
ram[64374] = {-9'd18,10'd383};
ram[64375] = {-9'd15,10'd386};
ram[64376] = {-9'd11,10'd389};
ram[64377] = {-9'd8,10'd392};
ram[64378] = {-9'd5,10'd395};
ram[64379] = {-9'd2,10'd398};
ram[64380] = {9'd1,-10'd399};
ram[64381] = {9'd4,-10'd396};
ram[64382] = {9'd7,-10'd393};
ram[64383] = {9'd10,-10'd390};
ram[64384] = {9'd10,-10'd390};
ram[64385] = {9'd14,-10'd387};
ram[64386] = {9'd17,-10'd384};
ram[64387] = {9'd20,-10'd381};
ram[64388] = {9'd23,-10'd377};
ram[64389] = {9'd26,-10'd374};
ram[64390] = {9'd29,-10'd371};
ram[64391] = {9'd32,-10'd368};
ram[64392] = {9'd36,-10'd365};
ram[64393] = {9'd39,-10'd362};
ram[64394] = {9'd42,-10'd359};
ram[64395] = {9'd45,-10'd355};
ram[64396] = {9'd48,-10'd352};
ram[64397] = {9'd51,-10'd349};
ram[64398] = {9'd54,-10'd346};
ram[64399] = {9'd58,-10'd343};
ram[64400] = {9'd61,-10'd340};
ram[64401] = {9'd64,-10'd337};
ram[64402] = {9'd67,-10'd334};
ram[64403] = {9'd70,-10'd330};
ram[64404] = {9'd73,-10'd327};
ram[64405] = {9'd76,-10'd324};
ram[64406] = {9'd80,-10'd321};
ram[64407] = {9'd83,-10'd318};
ram[64408] = {9'd86,-10'd315};
ram[64409] = {9'd89,-10'd312};
ram[64410] = {9'd92,-10'd308};
ram[64411] = {9'd95,-10'd305};
ram[64412] = {9'd98,-10'd302};
ram[64413] = {-9'd99,-10'd299};
ram[64414] = {-9'd96,-10'd296};
ram[64415] = {-9'd92,-10'd293};
ram[64416] = {-9'd89,-10'd290};
ram[64417] = {-9'd86,-10'd286};
ram[64418] = {-9'd83,-10'd283};
ram[64419] = {-9'd80,-10'd280};
ram[64420] = {-9'd77,-10'd277};
ram[64421] = {-9'd74,-10'd274};
ram[64422] = {-9'd70,-10'd271};
ram[64423] = {-9'd67,-10'd268};
ram[64424] = {-9'd64,-10'd264};
ram[64425] = {-9'd61,-10'd261};
ram[64426] = {-9'd58,-10'd258};
ram[64427] = {-9'd55,-10'd255};
ram[64428] = {-9'd52,-10'd252};
ram[64429] = {-9'd48,-10'd249};
ram[64430] = {-9'd45,-10'd246};
ram[64431] = {-9'd42,-10'd242};
ram[64432] = {-9'd39,-10'd239};
ram[64433] = {-9'd36,-10'd236};
ram[64434] = {-9'd33,-10'd233};
ram[64435] = {-9'd30,-10'd230};
ram[64436] = {-9'd26,-10'd227};
ram[64437] = {-9'd23,-10'd224};
ram[64438] = {-9'd20,-10'd220};
ram[64439] = {-9'd17,-10'd217};
ram[64440] = {-9'd14,-10'd214};
ram[64441] = {-9'd11,-10'd211};
ram[64442] = {-9'd8,-10'd208};
ram[64443] = {-9'd4,-10'd205};
ram[64444] = {-9'd1,-10'd202};
ram[64445] = {9'd2,-10'd198};
ram[64446] = {9'd5,-10'd195};
ram[64447] = {9'd8,-10'd192};
ram[64448] = {9'd11,-10'd189};
ram[64449] = {9'd14,-10'd186};
ram[64450] = {9'd18,-10'd183};
ram[64451] = {9'd21,-10'd180};
ram[64452] = {9'd24,-10'd176};
ram[64453] = {9'd27,-10'd173};
ram[64454] = {9'd30,-10'd170};
ram[64455] = {9'd33,-10'd167};
ram[64456] = {9'd36,-10'd164};
ram[64457] = {9'd40,-10'd161};
ram[64458] = {9'd43,-10'd158};
ram[64459] = {9'd46,-10'd154};
ram[64460] = {9'd49,-10'd151};
ram[64461] = {9'd52,-10'd148};
ram[64462] = {9'd55,-10'd145};
ram[64463] = {9'd58,-10'd142};
ram[64464] = {9'd62,-10'd139};
ram[64465] = {9'd65,-10'd136};
ram[64466] = {9'd68,-10'd132};
ram[64467] = {9'd71,-10'd129};
ram[64468] = {9'd74,-10'd126};
ram[64469] = {9'd77,-10'd123};
ram[64470] = {9'd80,-10'd120};
ram[64471] = {9'd84,-10'd117};
ram[64472] = {9'd87,-10'd114};
ram[64473] = {9'd90,-10'd110};
ram[64474] = {9'd93,-10'd107};
ram[64475] = {9'd96,-10'd104};
ram[64476] = {9'd99,-10'd101};
ram[64477] = {-9'd98,-10'd98};
ram[64478] = {-9'd95,-10'd95};
ram[64479] = {-9'd92,-10'd92};
ram[64480] = {-9'd88,-10'd88};
ram[64481] = {-9'd85,-10'd85};
ram[64482] = {-9'd82,-10'd82};
ram[64483] = {-9'd79,-10'd79};
ram[64484] = {-9'd76,-10'd76};
ram[64485] = {-9'd73,-10'd73};
ram[64486] = {-9'd70,-10'd70};
ram[64487] = {-9'd66,-10'd66};
ram[64488] = {-9'd63,-10'd63};
ram[64489] = {-9'd60,-10'd60};
ram[64490] = {-9'd57,-10'd57};
ram[64491] = {-9'd54,-10'd54};
ram[64492] = {-9'd51,-10'd51};
ram[64493] = {-9'd48,-10'd48};
ram[64494] = {-9'd44,-10'd44};
ram[64495] = {-9'd41,-10'd41};
ram[64496] = {-9'd38,-10'd38};
ram[64497] = {-9'd35,-10'd35};
ram[64498] = {-9'd32,-10'd32};
ram[64499] = {-9'd29,-10'd29};
ram[64500] = {-9'd26,-10'd26};
ram[64501] = {-9'd22,-10'd22};
ram[64502] = {-9'd19,-10'd19};
ram[64503] = {-9'd16,-10'd16};
ram[64504] = {-9'd13,-10'd13};
ram[64505] = {-9'd10,-10'd10};
ram[64506] = {-9'd7,-10'd7};
ram[64507] = {-9'd4,-10'd4};
ram[64508] = {9'd0,10'd0};
ram[64509] = {9'd3,10'd3};
ram[64510] = {9'd6,10'd6};
ram[64511] = {9'd9,10'd9};
ram[64512] = {9'd9,10'd9};
ram[64513] = {9'd12,10'd12};
ram[64514] = {9'd15,10'd15};
ram[64515] = {9'd18,10'd18};
ram[64516] = {9'd21,10'd21};
ram[64517] = {9'd25,10'd25};
ram[64518] = {9'd28,10'd28};
ram[64519] = {9'd31,10'd31};
ram[64520] = {9'd34,10'd34};
ram[64521] = {9'd37,10'd37};
ram[64522] = {9'd40,10'd40};
ram[64523] = {9'd43,10'd43};
ram[64524] = {9'd47,10'd47};
ram[64525] = {9'd50,10'd50};
ram[64526] = {9'd53,10'd53};
ram[64527] = {9'd56,10'd56};
ram[64528] = {9'd59,10'd59};
ram[64529] = {9'd62,10'd62};
ram[64530] = {9'd65,10'd65};
ram[64531] = {9'd69,10'd69};
ram[64532] = {9'd72,10'd72};
ram[64533] = {9'd75,10'd75};
ram[64534] = {9'd78,10'd78};
ram[64535] = {9'd81,10'd81};
ram[64536] = {9'd84,10'd84};
ram[64537] = {9'd87,10'd87};
ram[64538] = {9'd91,10'd91};
ram[64539] = {9'd94,10'd94};
ram[64540] = {9'd97,10'd97};
ram[64541] = {-9'd100,10'd100};
ram[64542] = {-9'd97,10'd103};
ram[64543] = {-9'd94,10'd106};
ram[64544] = {-9'd91,10'd109};
ram[64545] = {-9'd88,10'd113};
ram[64546] = {-9'd85,10'd116};
ram[64547] = {-9'd81,10'd119};
ram[64548] = {-9'd78,10'd122};
ram[64549] = {-9'd75,10'd125};
ram[64550] = {-9'd72,10'd128};
ram[64551] = {-9'd69,10'd131};
ram[64552] = {-9'd66,10'd135};
ram[64553] = {-9'd63,10'd138};
ram[64554] = {-9'd59,10'd141};
ram[64555] = {-9'd56,10'd144};
ram[64556] = {-9'd53,10'd147};
ram[64557] = {-9'd50,10'd150};
ram[64558] = {-9'd47,10'd153};
ram[64559] = {-9'd44,10'd157};
ram[64560] = {-9'd41,10'd160};
ram[64561] = {-9'd37,10'd163};
ram[64562] = {-9'd34,10'd166};
ram[64563] = {-9'd31,10'd169};
ram[64564] = {-9'd28,10'd172};
ram[64565] = {-9'd25,10'd175};
ram[64566] = {-9'd22,10'd179};
ram[64567] = {-9'd19,10'd182};
ram[64568] = {-9'd15,10'd185};
ram[64569] = {-9'd12,10'd188};
ram[64570] = {-9'd9,10'd191};
ram[64571] = {-9'd6,10'd194};
ram[64572] = {-9'd3,10'd197};
ram[64573] = {9'd0,10'd201};
ram[64574] = {9'd3,10'd204};
ram[64575] = {9'd7,10'd207};
ram[64576] = {9'd10,10'd210};
ram[64577] = {9'd13,10'd213};
ram[64578] = {9'd16,10'd216};
ram[64579] = {9'd19,10'd219};
ram[64580] = {9'd22,10'd223};
ram[64581] = {9'd25,10'd226};
ram[64582] = {9'd29,10'd229};
ram[64583] = {9'd32,10'd232};
ram[64584] = {9'd35,10'd235};
ram[64585] = {9'd38,10'd238};
ram[64586] = {9'd41,10'd241};
ram[64587] = {9'd44,10'd245};
ram[64588] = {9'd47,10'd248};
ram[64589] = {9'd51,10'd251};
ram[64590] = {9'd54,10'd254};
ram[64591] = {9'd57,10'd257};
ram[64592] = {9'd60,10'd260};
ram[64593] = {9'd63,10'd263};
ram[64594] = {9'd66,10'd267};
ram[64595] = {9'd69,10'd270};
ram[64596] = {9'd73,10'd273};
ram[64597] = {9'd76,10'd276};
ram[64598] = {9'd79,10'd279};
ram[64599] = {9'd82,10'd282};
ram[64600] = {9'd85,10'd285};
ram[64601] = {9'd88,10'd289};
ram[64602] = {9'd91,10'd292};
ram[64603] = {9'd95,10'd295};
ram[64604] = {9'd98,10'd298};
ram[64605] = {-9'd99,10'd301};
ram[64606] = {-9'd96,10'd304};
ram[64607] = {-9'd93,10'd307};
ram[64608] = {-9'd90,10'd311};
ram[64609] = {-9'd87,10'd314};
ram[64610] = {-9'd84,10'd317};
ram[64611] = {-9'd81,10'd320};
ram[64612] = {-9'd77,10'd323};
ram[64613] = {-9'd74,10'd326};
ram[64614] = {-9'd71,10'd329};
ram[64615] = {-9'd68,10'd333};
ram[64616] = {-9'd65,10'd336};
ram[64617] = {-9'd62,10'd339};
ram[64618] = {-9'd59,10'd342};
ram[64619] = {-9'd55,10'd345};
ram[64620] = {-9'd52,10'd348};
ram[64621] = {-9'd49,10'd351};
ram[64622] = {-9'd46,10'd354};
ram[64623] = {-9'd43,10'd358};
ram[64624] = {-9'd40,10'd361};
ram[64625] = {-9'd37,10'd364};
ram[64626] = {-9'd33,10'd367};
ram[64627] = {-9'd30,10'd370};
ram[64628] = {-9'd27,10'd373};
ram[64629] = {-9'd24,10'd376};
ram[64630] = {-9'd21,10'd380};
ram[64631] = {-9'd18,10'd383};
ram[64632] = {-9'd15,10'd386};
ram[64633] = {-9'd11,10'd389};
ram[64634] = {-9'd8,10'd392};
ram[64635] = {-9'd5,10'd395};
ram[64636] = {-9'd2,10'd398};
ram[64637] = {9'd1,-10'd399};
ram[64638] = {9'd4,-10'd396};
ram[64639] = {9'd7,-10'd393};
ram[64640] = {9'd7,-10'd393};
ram[64641] = {9'd10,-10'd390};
ram[64642] = {9'd14,-10'd387};
ram[64643] = {9'd17,-10'd384};
ram[64644] = {9'd20,-10'd381};
ram[64645] = {9'd23,-10'd377};
ram[64646] = {9'd26,-10'd374};
ram[64647] = {9'd29,-10'd371};
ram[64648] = {9'd32,-10'd368};
ram[64649] = {9'd36,-10'd365};
ram[64650] = {9'd39,-10'd362};
ram[64651] = {9'd42,-10'd359};
ram[64652] = {9'd45,-10'd355};
ram[64653] = {9'd48,-10'd352};
ram[64654] = {9'd51,-10'd349};
ram[64655] = {9'd54,-10'd346};
ram[64656] = {9'd58,-10'd343};
ram[64657] = {9'd61,-10'd340};
ram[64658] = {9'd64,-10'd337};
ram[64659] = {9'd67,-10'd334};
ram[64660] = {9'd70,-10'd330};
ram[64661] = {9'd73,-10'd327};
ram[64662] = {9'd76,-10'd324};
ram[64663] = {9'd80,-10'd321};
ram[64664] = {9'd83,-10'd318};
ram[64665] = {9'd86,-10'd315};
ram[64666] = {9'd89,-10'd312};
ram[64667] = {9'd92,-10'd308};
ram[64668] = {9'd95,-10'd305};
ram[64669] = {9'd98,-10'd302};
ram[64670] = {-9'd99,-10'd299};
ram[64671] = {-9'd96,-10'd296};
ram[64672] = {-9'd92,-10'd293};
ram[64673] = {-9'd89,-10'd290};
ram[64674] = {-9'd86,-10'd286};
ram[64675] = {-9'd83,-10'd283};
ram[64676] = {-9'd80,-10'd280};
ram[64677] = {-9'd77,-10'd277};
ram[64678] = {-9'd74,-10'd274};
ram[64679] = {-9'd70,-10'd271};
ram[64680] = {-9'd67,-10'd268};
ram[64681] = {-9'd64,-10'd264};
ram[64682] = {-9'd61,-10'd261};
ram[64683] = {-9'd58,-10'd258};
ram[64684] = {-9'd55,-10'd255};
ram[64685] = {-9'd52,-10'd252};
ram[64686] = {-9'd48,-10'd249};
ram[64687] = {-9'd45,-10'd246};
ram[64688] = {-9'd42,-10'd242};
ram[64689] = {-9'd39,-10'd239};
ram[64690] = {-9'd36,-10'd236};
ram[64691] = {-9'd33,-10'd233};
ram[64692] = {-9'd30,-10'd230};
ram[64693] = {-9'd26,-10'd227};
ram[64694] = {-9'd23,-10'd224};
ram[64695] = {-9'd20,-10'd220};
ram[64696] = {-9'd17,-10'd217};
ram[64697] = {-9'd14,-10'd214};
ram[64698] = {-9'd11,-10'd211};
ram[64699] = {-9'd8,-10'd208};
ram[64700] = {-9'd4,-10'd205};
ram[64701] = {-9'd1,-10'd202};
ram[64702] = {9'd2,-10'd198};
ram[64703] = {9'd5,-10'd195};
ram[64704] = {9'd8,-10'd192};
ram[64705] = {9'd11,-10'd189};
ram[64706] = {9'd14,-10'd186};
ram[64707] = {9'd18,-10'd183};
ram[64708] = {9'd21,-10'd180};
ram[64709] = {9'd24,-10'd176};
ram[64710] = {9'd27,-10'd173};
ram[64711] = {9'd30,-10'd170};
ram[64712] = {9'd33,-10'd167};
ram[64713] = {9'd36,-10'd164};
ram[64714] = {9'd40,-10'd161};
ram[64715] = {9'd43,-10'd158};
ram[64716] = {9'd46,-10'd154};
ram[64717] = {9'd49,-10'd151};
ram[64718] = {9'd52,-10'd148};
ram[64719] = {9'd55,-10'd145};
ram[64720] = {9'd58,-10'd142};
ram[64721] = {9'd62,-10'd139};
ram[64722] = {9'd65,-10'd136};
ram[64723] = {9'd68,-10'd132};
ram[64724] = {9'd71,-10'd129};
ram[64725] = {9'd74,-10'd126};
ram[64726] = {9'd77,-10'd123};
ram[64727] = {9'd80,-10'd120};
ram[64728] = {9'd84,-10'd117};
ram[64729] = {9'd87,-10'd114};
ram[64730] = {9'd90,-10'd110};
ram[64731] = {9'd93,-10'd107};
ram[64732] = {9'd96,-10'd104};
ram[64733] = {9'd99,-10'd101};
ram[64734] = {-9'd98,-10'd98};
ram[64735] = {-9'd95,-10'd95};
ram[64736] = {-9'd92,-10'd92};
ram[64737] = {-9'd88,-10'd88};
ram[64738] = {-9'd85,-10'd85};
ram[64739] = {-9'd82,-10'd82};
ram[64740] = {-9'd79,-10'd79};
ram[64741] = {-9'd76,-10'd76};
ram[64742] = {-9'd73,-10'd73};
ram[64743] = {-9'd70,-10'd70};
ram[64744] = {-9'd66,-10'd66};
ram[64745] = {-9'd63,-10'd63};
ram[64746] = {-9'd60,-10'd60};
ram[64747] = {-9'd57,-10'd57};
ram[64748] = {-9'd54,-10'd54};
ram[64749] = {-9'd51,-10'd51};
ram[64750] = {-9'd48,-10'd48};
ram[64751] = {-9'd44,-10'd44};
ram[64752] = {-9'd41,-10'd41};
ram[64753] = {-9'd38,-10'd38};
ram[64754] = {-9'd35,-10'd35};
ram[64755] = {-9'd32,-10'd32};
ram[64756] = {-9'd29,-10'd29};
ram[64757] = {-9'd26,-10'd26};
ram[64758] = {-9'd22,-10'd22};
ram[64759] = {-9'd19,-10'd19};
ram[64760] = {-9'd16,-10'd16};
ram[64761] = {-9'd13,-10'd13};
ram[64762] = {-9'd10,-10'd10};
ram[64763] = {-9'd7,-10'd7};
ram[64764] = {-9'd4,-10'd4};
ram[64765] = {9'd0,10'd0};
ram[64766] = {9'd3,10'd3};
ram[64767] = {9'd6,10'd6};
ram[64768] = {9'd6,10'd6};
ram[64769] = {9'd9,10'd9};
ram[64770] = {9'd12,10'd12};
ram[64771] = {9'd15,10'd15};
ram[64772] = {9'd18,10'd18};
ram[64773] = {9'd21,10'd21};
ram[64774] = {9'd25,10'd25};
ram[64775] = {9'd28,10'd28};
ram[64776] = {9'd31,10'd31};
ram[64777] = {9'd34,10'd34};
ram[64778] = {9'd37,10'd37};
ram[64779] = {9'd40,10'd40};
ram[64780] = {9'd43,10'd43};
ram[64781] = {9'd47,10'd47};
ram[64782] = {9'd50,10'd50};
ram[64783] = {9'd53,10'd53};
ram[64784] = {9'd56,10'd56};
ram[64785] = {9'd59,10'd59};
ram[64786] = {9'd62,10'd62};
ram[64787] = {9'd65,10'd65};
ram[64788] = {9'd69,10'd69};
ram[64789] = {9'd72,10'd72};
ram[64790] = {9'd75,10'd75};
ram[64791] = {9'd78,10'd78};
ram[64792] = {9'd81,10'd81};
ram[64793] = {9'd84,10'd84};
ram[64794] = {9'd87,10'd87};
ram[64795] = {9'd91,10'd91};
ram[64796] = {9'd94,10'd94};
ram[64797] = {9'd97,10'd97};
ram[64798] = {-9'd100,10'd100};
ram[64799] = {-9'd97,10'd103};
ram[64800] = {-9'd94,10'd106};
ram[64801] = {-9'd91,10'd109};
ram[64802] = {-9'd88,10'd113};
ram[64803] = {-9'd85,10'd116};
ram[64804] = {-9'd81,10'd119};
ram[64805] = {-9'd78,10'd122};
ram[64806] = {-9'd75,10'd125};
ram[64807] = {-9'd72,10'd128};
ram[64808] = {-9'd69,10'd131};
ram[64809] = {-9'd66,10'd135};
ram[64810] = {-9'd63,10'd138};
ram[64811] = {-9'd59,10'd141};
ram[64812] = {-9'd56,10'd144};
ram[64813] = {-9'd53,10'd147};
ram[64814] = {-9'd50,10'd150};
ram[64815] = {-9'd47,10'd153};
ram[64816] = {-9'd44,10'd157};
ram[64817] = {-9'd41,10'd160};
ram[64818] = {-9'd37,10'd163};
ram[64819] = {-9'd34,10'd166};
ram[64820] = {-9'd31,10'd169};
ram[64821] = {-9'd28,10'd172};
ram[64822] = {-9'd25,10'd175};
ram[64823] = {-9'd22,10'd179};
ram[64824] = {-9'd19,10'd182};
ram[64825] = {-9'd15,10'd185};
ram[64826] = {-9'd12,10'd188};
ram[64827] = {-9'd9,10'd191};
ram[64828] = {-9'd6,10'd194};
ram[64829] = {-9'd3,10'd197};
ram[64830] = {9'd0,10'd201};
ram[64831] = {9'd3,10'd204};
ram[64832] = {9'd7,10'd207};
ram[64833] = {9'd10,10'd210};
ram[64834] = {9'd13,10'd213};
ram[64835] = {9'd16,10'd216};
ram[64836] = {9'd19,10'd219};
ram[64837] = {9'd22,10'd223};
ram[64838] = {9'd25,10'd226};
ram[64839] = {9'd29,10'd229};
ram[64840] = {9'd32,10'd232};
ram[64841] = {9'd35,10'd235};
ram[64842] = {9'd38,10'd238};
ram[64843] = {9'd41,10'd241};
ram[64844] = {9'd44,10'd245};
ram[64845] = {9'd47,10'd248};
ram[64846] = {9'd51,10'd251};
ram[64847] = {9'd54,10'd254};
ram[64848] = {9'd57,10'd257};
ram[64849] = {9'd60,10'd260};
ram[64850] = {9'd63,10'd263};
ram[64851] = {9'd66,10'd267};
ram[64852] = {9'd69,10'd270};
ram[64853] = {9'd73,10'd273};
ram[64854] = {9'd76,10'd276};
ram[64855] = {9'd79,10'd279};
ram[64856] = {9'd82,10'd282};
ram[64857] = {9'd85,10'd285};
ram[64858] = {9'd88,10'd289};
ram[64859] = {9'd91,10'd292};
ram[64860] = {9'd95,10'd295};
ram[64861] = {9'd98,10'd298};
ram[64862] = {-9'd99,10'd301};
ram[64863] = {-9'd96,10'd304};
ram[64864] = {-9'd93,10'd307};
ram[64865] = {-9'd90,10'd311};
ram[64866] = {-9'd87,10'd314};
ram[64867] = {-9'd84,10'd317};
ram[64868] = {-9'd81,10'd320};
ram[64869] = {-9'd77,10'd323};
ram[64870] = {-9'd74,10'd326};
ram[64871] = {-9'd71,10'd329};
ram[64872] = {-9'd68,10'd333};
ram[64873] = {-9'd65,10'd336};
ram[64874] = {-9'd62,10'd339};
ram[64875] = {-9'd59,10'd342};
ram[64876] = {-9'd55,10'd345};
ram[64877] = {-9'd52,10'd348};
ram[64878] = {-9'd49,10'd351};
ram[64879] = {-9'd46,10'd354};
ram[64880] = {-9'd43,10'd358};
ram[64881] = {-9'd40,10'd361};
ram[64882] = {-9'd37,10'd364};
ram[64883] = {-9'd33,10'd367};
ram[64884] = {-9'd30,10'd370};
ram[64885] = {-9'd27,10'd373};
ram[64886] = {-9'd24,10'd376};
ram[64887] = {-9'd21,10'd380};
ram[64888] = {-9'd18,10'd383};
ram[64889] = {-9'd15,10'd386};
ram[64890] = {-9'd11,10'd389};
ram[64891] = {-9'd8,10'd392};
ram[64892] = {-9'd5,10'd395};
ram[64893] = {-9'd2,10'd398};
ram[64894] = {9'd1,-10'd399};
ram[64895] = {9'd4,-10'd396};
ram[64896] = {9'd4,-10'd396};
ram[64897] = {9'd7,-10'd393};
ram[64898] = {9'd10,-10'd390};
ram[64899] = {9'd14,-10'd387};
ram[64900] = {9'd17,-10'd384};
ram[64901] = {9'd20,-10'd381};
ram[64902] = {9'd23,-10'd377};
ram[64903] = {9'd26,-10'd374};
ram[64904] = {9'd29,-10'd371};
ram[64905] = {9'd32,-10'd368};
ram[64906] = {9'd36,-10'd365};
ram[64907] = {9'd39,-10'd362};
ram[64908] = {9'd42,-10'd359};
ram[64909] = {9'd45,-10'd355};
ram[64910] = {9'd48,-10'd352};
ram[64911] = {9'd51,-10'd349};
ram[64912] = {9'd54,-10'd346};
ram[64913] = {9'd58,-10'd343};
ram[64914] = {9'd61,-10'd340};
ram[64915] = {9'd64,-10'd337};
ram[64916] = {9'd67,-10'd334};
ram[64917] = {9'd70,-10'd330};
ram[64918] = {9'd73,-10'd327};
ram[64919] = {9'd76,-10'd324};
ram[64920] = {9'd80,-10'd321};
ram[64921] = {9'd83,-10'd318};
ram[64922] = {9'd86,-10'd315};
ram[64923] = {9'd89,-10'd312};
ram[64924] = {9'd92,-10'd308};
ram[64925] = {9'd95,-10'd305};
ram[64926] = {9'd98,-10'd302};
ram[64927] = {-9'd99,-10'd299};
ram[64928] = {-9'd96,-10'd296};
ram[64929] = {-9'd92,-10'd293};
ram[64930] = {-9'd89,-10'd290};
ram[64931] = {-9'd86,-10'd286};
ram[64932] = {-9'd83,-10'd283};
ram[64933] = {-9'd80,-10'd280};
ram[64934] = {-9'd77,-10'd277};
ram[64935] = {-9'd74,-10'd274};
ram[64936] = {-9'd70,-10'd271};
ram[64937] = {-9'd67,-10'd268};
ram[64938] = {-9'd64,-10'd264};
ram[64939] = {-9'd61,-10'd261};
ram[64940] = {-9'd58,-10'd258};
ram[64941] = {-9'd55,-10'd255};
ram[64942] = {-9'd52,-10'd252};
ram[64943] = {-9'd48,-10'd249};
ram[64944] = {-9'd45,-10'd246};
ram[64945] = {-9'd42,-10'd242};
ram[64946] = {-9'd39,-10'd239};
ram[64947] = {-9'd36,-10'd236};
ram[64948] = {-9'd33,-10'd233};
ram[64949] = {-9'd30,-10'd230};
ram[64950] = {-9'd26,-10'd227};
ram[64951] = {-9'd23,-10'd224};
ram[64952] = {-9'd20,-10'd220};
ram[64953] = {-9'd17,-10'd217};
ram[64954] = {-9'd14,-10'd214};
ram[64955] = {-9'd11,-10'd211};
ram[64956] = {-9'd8,-10'd208};
ram[64957] = {-9'd4,-10'd205};
ram[64958] = {-9'd1,-10'd202};
ram[64959] = {9'd2,-10'd198};
ram[64960] = {9'd5,-10'd195};
ram[64961] = {9'd8,-10'd192};
ram[64962] = {9'd11,-10'd189};
ram[64963] = {9'd14,-10'd186};
ram[64964] = {9'd18,-10'd183};
ram[64965] = {9'd21,-10'd180};
ram[64966] = {9'd24,-10'd176};
ram[64967] = {9'd27,-10'd173};
ram[64968] = {9'd30,-10'd170};
ram[64969] = {9'd33,-10'd167};
ram[64970] = {9'd36,-10'd164};
ram[64971] = {9'd40,-10'd161};
ram[64972] = {9'd43,-10'd158};
ram[64973] = {9'd46,-10'd154};
ram[64974] = {9'd49,-10'd151};
ram[64975] = {9'd52,-10'd148};
ram[64976] = {9'd55,-10'd145};
ram[64977] = {9'd58,-10'd142};
ram[64978] = {9'd62,-10'd139};
ram[64979] = {9'd65,-10'd136};
ram[64980] = {9'd68,-10'd132};
ram[64981] = {9'd71,-10'd129};
ram[64982] = {9'd74,-10'd126};
ram[64983] = {9'd77,-10'd123};
ram[64984] = {9'd80,-10'd120};
ram[64985] = {9'd84,-10'd117};
ram[64986] = {9'd87,-10'd114};
ram[64987] = {9'd90,-10'd110};
ram[64988] = {9'd93,-10'd107};
ram[64989] = {9'd96,-10'd104};
ram[64990] = {9'd99,-10'd101};
ram[64991] = {-9'd98,-10'd98};
ram[64992] = {-9'd95,-10'd95};
ram[64993] = {-9'd92,-10'd92};
ram[64994] = {-9'd88,-10'd88};
ram[64995] = {-9'd85,-10'd85};
ram[64996] = {-9'd82,-10'd82};
ram[64997] = {-9'd79,-10'd79};
ram[64998] = {-9'd76,-10'd76};
ram[64999] = {-9'd73,-10'd73};
ram[65000] = {-9'd70,-10'd70};
ram[65001] = {-9'd66,-10'd66};
ram[65002] = {-9'd63,-10'd63};
ram[65003] = {-9'd60,-10'd60};
ram[65004] = {-9'd57,-10'd57};
ram[65005] = {-9'd54,-10'd54};
ram[65006] = {-9'd51,-10'd51};
ram[65007] = {-9'd48,-10'd48};
ram[65008] = {-9'd44,-10'd44};
ram[65009] = {-9'd41,-10'd41};
ram[65010] = {-9'd38,-10'd38};
ram[65011] = {-9'd35,-10'd35};
ram[65012] = {-9'd32,-10'd32};
ram[65013] = {-9'd29,-10'd29};
ram[65014] = {-9'd26,-10'd26};
ram[65015] = {-9'd22,-10'd22};
ram[65016] = {-9'd19,-10'd19};
ram[65017] = {-9'd16,-10'd16};
ram[65018] = {-9'd13,-10'd13};
ram[65019] = {-9'd10,-10'd10};
ram[65020] = {-9'd7,-10'd7};
ram[65021] = {-9'd4,-10'd4};
ram[65022] = {9'd0,10'd0};
ram[65023] = {9'd3,10'd3};
ram[65024] = {9'd3,10'd3};
ram[65025] = {9'd6,10'd6};
ram[65026] = {9'd9,10'd9};
ram[65027] = {9'd12,10'd12};
ram[65028] = {9'd15,10'd15};
ram[65029] = {9'd18,10'd18};
ram[65030] = {9'd21,10'd21};
ram[65031] = {9'd25,10'd25};
ram[65032] = {9'd28,10'd28};
ram[65033] = {9'd31,10'd31};
ram[65034] = {9'd34,10'd34};
ram[65035] = {9'd37,10'd37};
ram[65036] = {9'd40,10'd40};
ram[65037] = {9'd43,10'd43};
ram[65038] = {9'd47,10'd47};
ram[65039] = {9'd50,10'd50};
ram[65040] = {9'd53,10'd53};
ram[65041] = {9'd56,10'd56};
ram[65042] = {9'd59,10'd59};
ram[65043] = {9'd62,10'd62};
ram[65044] = {9'd65,10'd65};
ram[65045] = {9'd69,10'd69};
ram[65046] = {9'd72,10'd72};
ram[65047] = {9'd75,10'd75};
ram[65048] = {9'd78,10'd78};
ram[65049] = {9'd81,10'd81};
ram[65050] = {9'd84,10'd84};
ram[65051] = {9'd87,10'd87};
ram[65052] = {9'd91,10'd91};
ram[65053] = {9'd94,10'd94};
ram[65054] = {9'd97,10'd97};
ram[65055] = {-9'd100,10'd100};
ram[65056] = {-9'd97,10'd103};
ram[65057] = {-9'd94,10'd106};
ram[65058] = {-9'd91,10'd109};
ram[65059] = {-9'd88,10'd113};
ram[65060] = {-9'd85,10'd116};
ram[65061] = {-9'd81,10'd119};
ram[65062] = {-9'd78,10'd122};
ram[65063] = {-9'd75,10'd125};
ram[65064] = {-9'd72,10'd128};
ram[65065] = {-9'd69,10'd131};
ram[65066] = {-9'd66,10'd135};
ram[65067] = {-9'd63,10'd138};
ram[65068] = {-9'd59,10'd141};
ram[65069] = {-9'd56,10'd144};
ram[65070] = {-9'd53,10'd147};
ram[65071] = {-9'd50,10'd150};
ram[65072] = {-9'd47,10'd153};
ram[65073] = {-9'd44,10'd157};
ram[65074] = {-9'd41,10'd160};
ram[65075] = {-9'd37,10'd163};
ram[65076] = {-9'd34,10'd166};
ram[65077] = {-9'd31,10'd169};
ram[65078] = {-9'd28,10'd172};
ram[65079] = {-9'd25,10'd175};
ram[65080] = {-9'd22,10'd179};
ram[65081] = {-9'd19,10'd182};
ram[65082] = {-9'd15,10'd185};
ram[65083] = {-9'd12,10'd188};
ram[65084] = {-9'd9,10'd191};
ram[65085] = {-9'd6,10'd194};
ram[65086] = {-9'd3,10'd197};
ram[65087] = {9'd0,10'd201};
ram[65088] = {9'd3,10'd204};
ram[65089] = {9'd7,10'd207};
ram[65090] = {9'd10,10'd210};
ram[65091] = {9'd13,10'd213};
ram[65092] = {9'd16,10'd216};
ram[65093] = {9'd19,10'd219};
ram[65094] = {9'd22,10'd223};
ram[65095] = {9'd25,10'd226};
ram[65096] = {9'd29,10'd229};
ram[65097] = {9'd32,10'd232};
ram[65098] = {9'd35,10'd235};
ram[65099] = {9'd38,10'd238};
ram[65100] = {9'd41,10'd241};
ram[65101] = {9'd44,10'd245};
ram[65102] = {9'd47,10'd248};
ram[65103] = {9'd51,10'd251};
ram[65104] = {9'd54,10'd254};
ram[65105] = {9'd57,10'd257};
ram[65106] = {9'd60,10'd260};
ram[65107] = {9'd63,10'd263};
ram[65108] = {9'd66,10'd267};
ram[65109] = {9'd69,10'd270};
ram[65110] = {9'd73,10'd273};
ram[65111] = {9'd76,10'd276};
ram[65112] = {9'd79,10'd279};
ram[65113] = {9'd82,10'd282};
ram[65114] = {9'd85,10'd285};
ram[65115] = {9'd88,10'd289};
ram[65116] = {9'd91,10'd292};
ram[65117] = {9'd95,10'd295};
ram[65118] = {9'd98,10'd298};
ram[65119] = {-9'd99,10'd301};
ram[65120] = {-9'd96,10'd304};
ram[65121] = {-9'd93,10'd307};
ram[65122] = {-9'd90,10'd311};
ram[65123] = {-9'd87,10'd314};
ram[65124] = {-9'd84,10'd317};
ram[65125] = {-9'd81,10'd320};
ram[65126] = {-9'd77,10'd323};
ram[65127] = {-9'd74,10'd326};
ram[65128] = {-9'd71,10'd329};
ram[65129] = {-9'd68,10'd333};
ram[65130] = {-9'd65,10'd336};
ram[65131] = {-9'd62,10'd339};
ram[65132] = {-9'd59,10'd342};
ram[65133] = {-9'd55,10'd345};
ram[65134] = {-9'd52,10'd348};
ram[65135] = {-9'd49,10'd351};
ram[65136] = {-9'd46,10'd354};
ram[65137] = {-9'd43,10'd358};
ram[65138] = {-9'd40,10'd361};
ram[65139] = {-9'd37,10'd364};
ram[65140] = {-9'd33,10'd367};
ram[65141] = {-9'd30,10'd370};
ram[65142] = {-9'd27,10'd373};
ram[65143] = {-9'd24,10'd376};
ram[65144] = {-9'd21,10'd380};
ram[65145] = {-9'd18,10'd383};
ram[65146] = {-9'd15,10'd386};
ram[65147] = {-9'd11,10'd389};
ram[65148] = {-9'd8,10'd392};
ram[65149] = {-9'd5,10'd395};
ram[65150] = {-9'd2,10'd398};
ram[65151] = {9'd1,-10'd399};
ram[65152] = {9'd1,-10'd399};
ram[65153] = {9'd4,-10'd396};
ram[65154] = {9'd7,-10'd393};
ram[65155] = {9'd10,-10'd390};
ram[65156] = {9'd14,-10'd387};
ram[65157] = {9'd17,-10'd384};
ram[65158] = {9'd20,-10'd381};
ram[65159] = {9'd23,-10'd377};
ram[65160] = {9'd26,-10'd374};
ram[65161] = {9'd29,-10'd371};
ram[65162] = {9'd32,-10'd368};
ram[65163] = {9'd36,-10'd365};
ram[65164] = {9'd39,-10'd362};
ram[65165] = {9'd42,-10'd359};
ram[65166] = {9'd45,-10'd355};
ram[65167] = {9'd48,-10'd352};
ram[65168] = {9'd51,-10'd349};
ram[65169] = {9'd54,-10'd346};
ram[65170] = {9'd58,-10'd343};
ram[65171] = {9'd61,-10'd340};
ram[65172] = {9'd64,-10'd337};
ram[65173] = {9'd67,-10'd334};
ram[65174] = {9'd70,-10'd330};
ram[65175] = {9'd73,-10'd327};
ram[65176] = {9'd76,-10'd324};
ram[65177] = {9'd80,-10'd321};
ram[65178] = {9'd83,-10'd318};
ram[65179] = {9'd86,-10'd315};
ram[65180] = {9'd89,-10'd312};
ram[65181] = {9'd92,-10'd308};
ram[65182] = {9'd95,-10'd305};
ram[65183] = {9'd98,-10'd302};
ram[65184] = {-9'd99,-10'd299};
ram[65185] = {-9'd96,-10'd296};
ram[65186] = {-9'd92,-10'd293};
ram[65187] = {-9'd89,-10'd290};
ram[65188] = {-9'd86,-10'd286};
ram[65189] = {-9'd83,-10'd283};
ram[65190] = {-9'd80,-10'd280};
ram[65191] = {-9'd77,-10'd277};
ram[65192] = {-9'd74,-10'd274};
ram[65193] = {-9'd70,-10'd271};
ram[65194] = {-9'd67,-10'd268};
ram[65195] = {-9'd64,-10'd264};
ram[65196] = {-9'd61,-10'd261};
ram[65197] = {-9'd58,-10'd258};
ram[65198] = {-9'd55,-10'd255};
ram[65199] = {-9'd52,-10'd252};
ram[65200] = {-9'd48,-10'd249};
ram[65201] = {-9'd45,-10'd246};
ram[65202] = {-9'd42,-10'd242};
ram[65203] = {-9'd39,-10'd239};
ram[65204] = {-9'd36,-10'd236};
ram[65205] = {-9'd33,-10'd233};
ram[65206] = {-9'd30,-10'd230};
ram[65207] = {-9'd26,-10'd227};
ram[65208] = {-9'd23,-10'd224};
ram[65209] = {-9'd20,-10'd220};
ram[65210] = {-9'd17,-10'd217};
ram[65211] = {-9'd14,-10'd214};
ram[65212] = {-9'd11,-10'd211};
ram[65213] = {-9'd8,-10'd208};
ram[65214] = {-9'd4,-10'd205};
ram[65215] = {-9'd1,-10'd202};
ram[65216] = {9'd2,-10'd198};
ram[65217] = {9'd5,-10'd195};
ram[65218] = {9'd8,-10'd192};
ram[65219] = {9'd11,-10'd189};
ram[65220] = {9'd14,-10'd186};
ram[65221] = {9'd18,-10'd183};
ram[65222] = {9'd21,-10'd180};
ram[65223] = {9'd24,-10'd176};
ram[65224] = {9'd27,-10'd173};
ram[65225] = {9'd30,-10'd170};
ram[65226] = {9'd33,-10'd167};
ram[65227] = {9'd36,-10'd164};
ram[65228] = {9'd40,-10'd161};
ram[65229] = {9'd43,-10'd158};
ram[65230] = {9'd46,-10'd154};
ram[65231] = {9'd49,-10'd151};
ram[65232] = {9'd52,-10'd148};
ram[65233] = {9'd55,-10'd145};
ram[65234] = {9'd58,-10'd142};
ram[65235] = {9'd62,-10'd139};
ram[65236] = {9'd65,-10'd136};
ram[65237] = {9'd68,-10'd132};
ram[65238] = {9'd71,-10'd129};
ram[65239] = {9'd74,-10'd126};
ram[65240] = {9'd77,-10'd123};
ram[65241] = {9'd80,-10'd120};
ram[65242] = {9'd84,-10'd117};
ram[65243] = {9'd87,-10'd114};
ram[65244] = {9'd90,-10'd110};
ram[65245] = {9'd93,-10'd107};
ram[65246] = {9'd96,-10'd104};
ram[65247] = {9'd99,-10'd101};
ram[65248] = {-9'd98,-10'd98};
ram[65249] = {-9'd95,-10'd95};
ram[65250] = {-9'd92,-10'd92};
ram[65251] = {-9'd88,-10'd88};
ram[65252] = {-9'd85,-10'd85};
ram[65253] = {-9'd82,-10'd82};
ram[65254] = {-9'd79,-10'd79};
ram[65255] = {-9'd76,-10'd76};
ram[65256] = {-9'd73,-10'd73};
ram[65257] = {-9'd70,-10'd70};
ram[65258] = {-9'd66,-10'd66};
ram[65259] = {-9'd63,-10'd63};
ram[65260] = {-9'd60,-10'd60};
ram[65261] = {-9'd57,-10'd57};
ram[65262] = {-9'd54,-10'd54};
ram[65263] = {-9'd51,-10'd51};
ram[65264] = {-9'd48,-10'd48};
ram[65265] = {-9'd44,-10'd44};
ram[65266] = {-9'd41,-10'd41};
ram[65267] = {-9'd38,-10'd38};
ram[65268] = {-9'd35,-10'd35};
ram[65269] = {-9'd32,-10'd32};
ram[65270] = {-9'd29,-10'd29};
ram[65271] = {-9'd26,-10'd26};
ram[65272] = {-9'd22,-10'd22};
ram[65273] = {-9'd19,-10'd19};
ram[65274] = {-9'd16,-10'd16};
ram[65275] = {-9'd13,-10'd13};
ram[65276] = {-9'd10,-10'd10};
ram[65277] = {-9'd7,-10'd7};
ram[65278] = {-9'd4,-10'd4};
ram[65279] = {9'd0,10'd0};
ram[65280] = {9'd0,10'd0};
ram[65281] = {9'd3,10'd3};
ram[65282] = {9'd6,10'd6};
ram[65283] = {9'd9,10'd9};
ram[65284] = {9'd12,10'd12};
ram[65285] = {9'd15,10'd15};
ram[65286] = {9'd18,10'd18};
ram[65287] = {9'd21,10'd21};
ram[65288] = {9'd25,10'd25};
ram[65289] = {9'd28,10'd28};
ram[65290] = {9'd31,10'd31};
ram[65291] = {9'd34,10'd34};
ram[65292] = {9'd37,10'd37};
ram[65293] = {9'd40,10'd40};
ram[65294] = {9'd43,10'd43};
ram[65295] = {9'd47,10'd47};
ram[65296] = {9'd50,10'd50};
ram[65297] = {9'd53,10'd53};
ram[65298] = {9'd56,10'd56};
ram[65299] = {9'd59,10'd59};
ram[65300] = {9'd62,10'd62};
ram[65301] = {9'd65,10'd65};
ram[65302] = {9'd69,10'd69};
ram[65303] = {9'd72,10'd72};
ram[65304] = {9'd75,10'd75};
ram[65305] = {9'd78,10'd78};
ram[65306] = {9'd81,10'd81};
ram[65307] = {9'd84,10'd84};
ram[65308] = {9'd87,10'd87};
ram[65309] = {9'd91,10'd91};
ram[65310] = {9'd94,10'd94};
ram[65311] = {9'd97,10'd97};
ram[65312] = {-9'd100,10'd100};
ram[65313] = {-9'd97,10'd103};
ram[65314] = {-9'd94,10'd106};
ram[65315] = {-9'd91,10'd109};
ram[65316] = {-9'd88,10'd113};
ram[65317] = {-9'd85,10'd116};
ram[65318] = {-9'd81,10'd119};
ram[65319] = {-9'd78,10'd122};
ram[65320] = {-9'd75,10'd125};
ram[65321] = {-9'd72,10'd128};
ram[65322] = {-9'd69,10'd131};
ram[65323] = {-9'd66,10'd135};
ram[65324] = {-9'd63,10'd138};
ram[65325] = {-9'd59,10'd141};
ram[65326] = {-9'd56,10'd144};
ram[65327] = {-9'd53,10'd147};
ram[65328] = {-9'd50,10'd150};
ram[65329] = {-9'd47,10'd153};
ram[65330] = {-9'd44,10'd157};
ram[65331] = {-9'd41,10'd160};
ram[65332] = {-9'd37,10'd163};
ram[65333] = {-9'd34,10'd166};
ram[65334] = {-9'd31,10'd169};
ram[65335] = {-9'd28,10'd172};
ram[65336] = {-9'd25,10'd175};
ram[65337] = {-9'd22,10'd179};
ram[65338] = {-9'd19,10'd182};
ram[65339] = {-9'd15,10'd185};
ram[65340] = {-9'd12,10'd188};
ram[65341] = {-9'd9,10'd191};
ram[65342] = {-9'd6,10'd194};
ram[65343] = {-9'd3,10'd197};
ram[65344] = {9'd0,10'd201};
ram[65345] = {9'd3,10'd204};
ram[65346] = {9'd7,10'd207};
ram[65347] = {9'd10,10'd210};
ram[65348] = {9'd13,10'd213};
ram[65349] = {9'd16,10'd216};
ram[65350] = {9'd19,10'd219};
ram[65351] = {9'd22,10'd223};
ram[65352] = {9'd25,10'd226};
ram[65353] = {9'd29,10'd229};
ram[65354] = {9'd32,10'd232};
ram[65355] = {9'd35,10'd235};
ram[65356] = {9'd38,10'd238};
ram[65357] = {9'd41,10'd241};
ram[65358] = {9'd44,10'd245};
ram[65359] = {9'd47,10'd248};
ram[65360] = {9'd51,10'd251};
ram[65361] = {9'd54,10'd254};
ram[65362] = {9'd57,10'd257};
ram[65363] = {9'd60,10'd260};
ram[65364] = {9'd63,10'd263};
ram[65365] = {9'd66,10'd267};
ram[65366] = {9'd69,10'd270};
ram[65367] = {9'd73,10'd273};
ram[65368] = {9'd76,10'd276};
ram[65369] = {9'd79,10'd279};
ram[65370] = {9'd82,10'd282};
ram[65371] = {9'd85,10'd285};
ram[65372] = {9'd88,10'd289};
ram[65373] = {9'd91,10'd292};
ram[65374] = {9'd95,10'd295};
ram[65375] = {9'd98,10'd298};
ram[65376] = {-9'd99,10'd301};
ram[65377] = {-9'd96,10'd304};
ram[65378] = {-9'd93,10'd307};
ram[65379] = {-9'd90,10'd311};
ram[65380] = {-9'd87,10'd314};
ram[65381] = {-9'd84,10'd317};
ram[65382] = {-9'd81,10'd320};
ram[65383] = {-9'd77,10'd323};
ram[65384] = {-9'd74,10'd326};
ram[65385] = {-9'd71,10'd329};
ram[65386] = {-9'd68,10'd333};
ram[65387] = {-9'd65,10'd336};
ram[65388] = {-9'd62,10'd339};
ram[65389] = {-9'd59,10'd342};
ram[65390] = {-9'd55,10'd345};
ram[65391] = {-9'd52,10'd348};
ram[65392] = {-9'd49,10'd351};
ram[65393] = {-9'd46,10'd354};
ram[65394] = {-9'd43,10'd358};
ram[65395] = {-9'd40,10'd361};
ram[65396] = {-9'd37,10'd364};
ram[65397] = {-9'd33,10'd367};
ram[65398] = {-9'd30,10'd370};
ram[65399] = {-9'd27,10'd373};
ram[65400] = {-9'd24,10'd376};
ram[65401] = {-9'd21,10'd380};
ram[65402] = {-9'd18,10'd383};
ram[65403] = {-9'd15,10'd386};
ram[65404] = {-9'd11,10'd389};
ram[65405] = {-9'd8,10'd392};
ram[65406] = {-9'd5,10'd395};
ram[65407] = {-9'd2,10'd398};
ram[65408] = {-9'd2,10'd398};
ram[65409] = {9'd1,-10'd399};
ram[65410] = {9'd4,-10'd396};
ram[65411] = {9'd7,-10'd393};
ram[65412] = {9'd10,-10'd390};
ram[65413] = {9'd14,-10'd387};
ram[65414] = {9'd17,-10'd384};
ram[65415] = {9'd20,-10'd381};
ram[65416] = {9'd23,-10'd377};
ram[65417] = {9'd26,-10'd374};
ram[65418] = {9'd29,-10'd371};
ram[65419] = {9'd32,-10'd368};
ram[65420] = {9'd36,-10'd365};
ram[65421] = {9'd39,-10'd362};
ram[65422] = {9'd42,-10'd359};
ram[65423] = {9'd45,-10'd355};
ram[65424] = {9'd48,-10'd352};
ram[65425] = {9'd51,-10'd349};
ram[65426] = {9'd54,-10'd346};
ram[65427] = {9'd58,-10'd343};
ram[65428] = {9'd61,-10'd340};
ram[65429] = {9'd64,-10'd337};
ram[65430] = {9'd67,-10'd334};
ram[65431] = {9'd70,-10'd330};
ram[65432] = {9'd73,-10'd327};
ram[65433] = {9'd76,-10'd324};
ram[65434] = {9'd80,-10'd321};
ram[65435] = {9'd83,-10'd318};
ram[65436] = {9'd86,-10'd315};
ram[65437] = {9'd89,-10'd312};
ram[65438] = {9'd92,-10'd308};
ram[65439] = {9'd95,-10'd305};
ram[65440] = {9'd98,-10'd302};
ram[65441] = {-9'd99,-10'd299};
ram[65442] = {-9'd96,-10'd296};
ram[65443] = {-9'd92,-10'd293};
ram[65444] = {-9'd89,-10'd290};
ram[65445] = {-9'd86,-10'd286};
ram[65446] = {-9'd83,-10'd283};
ram[65447] = {-9'd80,-10'd280};
ram[65448] = {-9'd77,-10'd277};
ram[65449] = {-9'd74,-10'd274};
ram[65450] = {-9'd70,-10'd271};
ram[65451] = {-9'd67,-10'd268};
ram[65452] = {-9'd64,-10'd264};
ram[65453] = {-9'd61,-10'd261};
ram[65454] = {-9'd58,-10'd258};
ram[65455] = {-9'd55,-10'd255};
ram[65456] = {-9'd52,-10'd252};
ram[65457] = {-9'd48,-10'd249};
ram[65458] = {-9'd45,-10'd246};
ram[65459] = {-9'd42,-10'd242};
ram[65460] = {-9'd39,-10'd239};
ram[65461] = {-9'd36,-10'd236};
ram[65462] = {-9'd33,-10'd233};
ram[65463] = {-9'd30,-10'd230};
ram[65464] = {-9'd26,-10'd227};
ram[65465] = {-9'd23,-10'd224};
ram[65466] = {-9'd20,-10'd220};
ram[65467] = {-9'd17,-10'd217};
ram[65468] = {-9'd14,-10'd214};
ram[65469] = {-9'd11,-10'd211};
ram[65470] = {-9'd8,-10'd208};
ram[65471] = {-9'd4,-10'd205};
ram[65472] = {-9'd1,-10'd202};
ram[65473] = {9'd2,-10'd198};
ram[65474] = {9'd5,-10'd195};
ram[65475] = {9'd8,-10'd192};
ram[65476] = {9'd11,-10'd189};
ram[65477] = {9'd14,-10'd186};
ram[65478] = {9'd18,-10'd183};
ram[65479] = {9'd21,-10'd180};
ram[65480] = {9'd24,-10'd176};
ram[65481] = {9'd27,-10'd173};
ram[65482] = {9'd30,-10'd170};
ram[65483] = {9'd33,-10'd167};
ram[65484] = {9'd36,-10'd164};
ram[65485] = {9'd40,-10'd161};
ram[65486] = {9'd43,-10'd158};
ram[65487] = {9'd46,-10'd154};
ram[65488] = {9'd49,-10'd151};
ram[65489] = {9'd52,-10'd148};
ram[65490] = {9'd55,-10'd145};
ram[65491] = {9'd58,-10'd142};
ram[65492] = {9'd62,-10'd139};
ram[65493] = {9'd65,-10'd136};
ram[65494] = {9'd68,-10'd132};
ram[65495] = {9'd71,-10'd129};
ram[65496] = {9'd74,-10'd126};
ram[65497] = {9'd77,-10'd123};
ram[65498] = {9'd80,-10'd120};
ram[65499] = {9'd84,-10'd117};
ram[65500] = {9'd87,-10'd114};
ram[65501] = {9'd90,-10'd110};
ram[65502] = {9'd93,-10'd107};
ram[65503] = {9'd96,-10'd104};
ram[65504] = {9'd99,-10'd101};
ram[65505] = {-9'd98,-10'd98};
ram[65506] = {-9'd95,-10'd95};
ram[65507] = {-9'd92,-10'd92};
ram[65508] = {-9'd88,-10'd88};
ram[65509] = {-9'd85,-10'd85};
ram[65510] = {-9'd82,-10'd82};
ram[65511] = {-9'd79,-10'd79};
ram[65512] = {-9'd76,-10'd76};
ram[65513] = {-9'd73,-10'd73};
ram[65514] = {-9'd70,-10'd70};
ram[65515] = {-9'd66,-10'd66};
ram[65516] = {-9'd63,-10'd63};
ram[65517] = {-9'd60,-10'd60};
ram[65518] = {-9'd57,-10'd57};
ram[65519] = {-9'd54,-10'd54};
ram[65520] = {-9'd51,-10'd51};
ram[65521] = {-9'd48,-10'd48};
ram[65522] = {-9'd44,-10'd44};
ram[65523] = {-9'd41,-10'd41};
ram[65524] = {-9'd38,-10'd38};
ram[65525] = {-9'd35,-10'd35};
ram[65526] = {-9'd32,-10'd32};
ram[65527] = {-9'd29,-10'd29};
ram[65528] = {-9'd26,-10'd26};
ram[65529] = {-9'd22,-10'd22};
ram[65530] = {-9'd19,-10'd19};
ram[65531] = {-9'd16,-10'd16};
ram[65532] = {-9'd13,-10'd13};
ram[65533] = {-9'd10,-10'd10};
ram[65534] = {-9'd7,-10'd7};
ram[65535] = {-9'd4,-10'd4};

end

assign test_pos={phase_acum_mod[8:1],input_angles[8:1]};
//assign test_pos={phase_acum_mod[8-1:1-1],input_angles[8:1]};

always @ ( posedge clk ) begin
	begin
		{phi_error,val_engle}<=ram[{phase_acum_mod[8:1],input_angles[8:1]}];		
	end
			
end

endmodule 
