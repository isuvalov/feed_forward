library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
entity table_demod is
	generic(
		BIT_IN:integer:=8;
		BIT_OUT:integer:=8 
	);
	 port(
		  clk : in std_logic;
		  i_ce: in std_logic;
	      sample_in_re: in std_logic_vector(BIT_IN-1 downto 0);
	      sample_in_im: in std_logic_vector(BIT_IN-1 downto 0);
		  o_ce: out std_logic;
	      sample_out_re: out std_logic_vector(BIT_OUT-1 downto 0);
	      sample_out_im: out std_logic_vector(BIT_OUT-1 downto 0)
		 );
    end table_demod;
architecture table_demod of table_demod is
type Tmem is array (0 to 65535) of std_logic_vector(7 downto 0);
constant mem_re:Tmem:=  (
"01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01011010", "01110010", "01111000", "01111011", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111011", "01111000", "01110010", "01011010", "01111111", "01110010", "01011010", "01101010", "01110010", "01110110", "01111000", "01111010", "01111011", 
"01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111011", 
"01111010", "01111000", "01110110", "01110010", "01101010", "01011010", "01110010", "01111111", "01111000", "01101010", "01011010", "01100110", "01101101", "01110010", "01110101", "01110111", "01111000", "01111010", "01111011", "01111011", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111000", "01110111", "01110101", "01110010", "01101101", "01100110", 
"01011010", "01101010", "01111000", "01111111", "01111011", "01110010", "01100110", "01011010", "01100011", "01101010", "01101110", "01110010", "01110100", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111011", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110100", "01110010", "01101110", "01101010", "01100011", "01011010", "01100110", "01110010", "01111011", "01111111", 
"01111101", "01110110", "01101101", "01100011", "01011010", "01100010", "01100111", "01101100", "01101111", "01110010", "01110100", "01110101", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", 
"01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", 
"01111000", "01111000", "01110111", "01110101", "01110100", "01110010", "01101111", "01101100", "01100111", "01100010", "01011010", "01100011", "01101101", "01110110", "01111101", "01111111", "01111101", "01111000", "01110010", "01101010", 
"01100010", "01011010", "01100000", "01100110", "01101010", "01101101", "01101111", "01110010", "01110011", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110011", "01110010", 
"01101111", "01101101", "01101010", "01100110", "01100000", "01011010", "01100010", "01101010", "01110010", "01111000", "01111101", "01111111", "01111110", "01111010", "01110101", "01101110", "01100111", "01100000", "01011010", "01100000", 
"01100100", "01101000", "01101011", "01101110", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", 
"01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101110", "01101011", "01101000", "01100100", "01100000", 
"01011010", "01100000", "01100111", "01101110", "01110101", "01111010", "01111110", "01111111", "01111110", "01111011", "01110111", "01110010", "01101100", "01100110", "01100000", "01011010", "01011111", "01100011", "01100111", "01101010", 
"01101100", "01101110", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101110", "01101100", "01101010", "01100111", "01100011", "01011111", "01011010", "01100000", "01100110", "01101100", "01110010", 
"01110111", "01111011", "01111110", "01111111", "01111110", "01111100", "01111000", "01110100", "01101111", "01101010", "01100100", "01011111", "01011010", "01011110", "01100010", "01100110", "01101000", "01101011", "01101101", "01101111", 
"01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", 
"01110011", "01110010", "01110000", "01101111", "01101101", "01101011", "01101000", "01100110", "01100010", "01011110", "01011010", "01011111", "01100100", "01101010", "01101111", "01110100", "01111000", "01111100", "01111110", "01111111", 
"01111110", "01111101", "01111010", "01110110", "01110010", "01101101", "01101000", "01100011", "01011110", "01011010", "01011110", "01100010", "01100101", "01100111", "01101010", "01101100", "01101101", "01101111", "01110000", "01110010", 
"01110011", "01110100", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110000", "01101111", "01101101", "01101100", 
"01101010", "01100111", "01100101", "01100010", "01011110", "01011010", "01011110", "01100011", "01101000", "01101101", "01110010", "01110110", "01111010", "01111101", "01111110", "01111111", "01111110", "01111101", "01111011", "01110111", 
"01110100", "01101111", "01101011", "01100111", "01100010", "01011110", "01011010", "01011110", "01100001", "01100100", "01100110", "01101001", "01101011", "01101100", "01101110", "01101111", "01110001", "01110010", "01110011", "01110011", 
"01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01101111", "01101110", "01101100", "01101011", "01101001", "01100110", "01100100", "01100001", "01011110", 
"01011010", "01011110", "01100010", "01100111", "01101011", "01101111", "01110100", "01110111", "01111011", "01111101", "01111110", "01111111", "01111111", "01111101", "01111011", "01111000", "01110101", "01110010", "01101110", "01101010", 
"01100110", "01100010", "01011110", "01011010", "01011101", "01100000", "01100011", "01100110", "01101000", "01101010", "01101011", "01101101", "01101110", "01101111", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", 
"01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", 
"01110100", "01110011", "01110010", "01110010", "01110001", "01101111", "01101110", "01101101", "01101011", "01101010", "01101000", "01100110", "01100011", "01100000", "01011101", "01011010", "01011110", "01100010", "01100110", "01101010", 
"01101110", "01110010", "01110101", "01111000", "01111011", "01111101", "01111111", "01111111", "01111111", "01111110", "01111100", "01111001", "01110111", "01110011", "01110000", "01101100", "01101000", "01100101", "01100001", "01011101", 
"01011010", "01011101", "01100000", "01100011", "01100101", "01100111", "01101001", "01101010", "01101100", "01101101", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", 
"01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", 
"01101111", "01101101", "01101100", "01101010", "01101001", "01100111", "01100101", "01100011", "01100000", "01011101", "01011010", "01011101", "01100001", "01100101", "01101000", "01101100", "01110000", "01110011", "01110111", "01111001", 
"01111100", "01111110", "01111111", "01111111", "01111111", "01111110", "01111100", "01111010", "01111000", "01110101", "01110010", "01101110", "01101011", "01100111", "01100100", "01100000", "01011101", "01011010", "01011101", "01100000", 
"01100010", "01100100", "01100110", "01101000", "01101010", "01101011", "01101100", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", 
"01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101100", "01101011", "01101010", "01101000", 
"01100110", "01100100", "01100010", "01100000", "01011101", "01011010", "01011101", "01100000", "01100100", "01100111", "01101011", "01101110", "01110010", "01110101", "01111000", "01111010", "01111100", "01111110", "01111111", "01111111", 
"01111111", "01111110", "01111101", "01111011", "01111000", "01110110", "01110011", "01110000", "01101101", "01101010", "01100110", "01100011", "01100000", "01011101", "01011010", "01011101", "01011111", "01100010", "01100100", "01100110", 
"01100111", "01101001", "01101010", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", 
"01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", 
"01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101010", "01101001", "01100111", "01100110", "01100100", "01100010", "01011111", "01011101", 
"01011010", "01011101", "01100000", "01100011", "01100110", "01101010", "01101101", "01110000", "01110011", "01110110", "01111000", "01111011", "01111101", "01111110", "01111111", "01111111", "01111111", "01111110", "01111101", "01111011", 
"01111001", "01110111", "01110100", "01110010", "01101111", "01101100", "01101001", "01100110", "01100011", "01100000", "01011101", "01011010", "01011100", "01011111", "01100001", "01100011", "01100101", "01100111", "01101000", "01101010", 
"01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", 
"01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", 
"01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101000", "01100111", "01100101", "01100011", "01100001", "01011111", "01011100", "01011010", "01011101", "01100000", "01100011", "01100110", 
"01101001", "01101100", "01101111", "01110010", "01110100", "01110111", "01111001", "01111011", "01111101", "01111110", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111010", "01111000", "01110101", "01110011", 
"01110000", "01101101", "01101011", "01101000", "01100101", "01100010", "01011111", "01011100", "01011010", "01011100", "01011111", "01100001", "01100011", "01100100", "01100110", "01101000", "01101001", "01101010", "01101011", "01101101", 
"01101110", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", 
"01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101110", "01101101", 
"01101011", "01101010", "01101001", "01101000", "01100110", "01100100", "01100011", "01100001", "01011111", "01011100", "01011010", "01011100", "01011111", "01100010", "01100101", "01101000", "01101011", "01101101", "01110000", "01110011", 
"01110101", "01111000", "01111010", "01111100", "01111101", "01111110", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111010", "01111000", "01110110", "01110100", "01110010", "01101111", "01101100", "01101010", 
"01100111", "01100100", "01100010", "01011111", "01011100", "01011010", "01011100", "01011110", "01100000", "01100010", "01100100", "01100110", "01100111", "01101000", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", 
"01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", 
"01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", 
"01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101000", "01100111", "01100110", 
"01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011111", "01100010", "01100100", "01100111", "01101010", "01101100", "01101111", "01110010", "01110100", "01110110", "01111000", "01111010", "01111100", 
"01111101", "01111110", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111011", "01111001", "01110111", "01110101", "01110011", "01110000", "01101110", "01101011", "01101001", "01100110", "01100100", "01100001", 
"01011111", "01011100", "01011010", "01011100", "01011110", "01100000", "01100010", "01100100", "01100101", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110000", 
"01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", 
"01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100101", "01100100", "01100010", "01100000", "01011110", "01011100", 
"01011010", "01011100", "01011111", "01100001", "01100100", "01100110", "01101001", "01101011", "01101110", "01110000", "01110011", "01110101", "01110111", "01111001", "01111011", "01111100", "01111101", "01111110", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111101", "01111011", "01111010", "01111000", "01110110", "01110100", "01110010", "01101111", "01101101", "01101010", "01101000", "01100110", "01100011", "01100001", "01011110", "01011100", "01011010", 
"01011100", "01011110", "01100000", "01100010", "01100011", "01100101", "01100110", "01100111", "01101001", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", 
"01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", 
"01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101001", "01100111", "01100110", "01100101", "01100011", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011110", "01100001", "01100011", 
"01100110", "01101000", "01101010", "01101101", "01101111", "01110010", "01110100", "01110110", "01111000", "01111010", "01111011", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", 
"01111100", "01111010", "01111000", "01110111", "01110101", "01110011", "01110001", "01101110", "01101100", "01101010", "01100111", "01100101", "01100011", "01100000", "01011110", "01011100", "01011010", "01011100", "01011110", "01100000", 
"01100001", "01100011", "01100100", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", 
"01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101011", "01101010", 
"01101001", "01101000", "01100111", "01100110", "01100100", "01100011", "01100001", "01100000", "01011110", "01011100", "01011010", "01011100", "01011110", "01100000", "01100011", "01100101", "01100111", "01101010", "01101100", "01101110", 
"01110001", "01110011", "01110101", "01110111", "01111000", "01111010", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111001", "01110111", 
"01110110", "01110100", "01110010", "01101111", "01101101", "01101011", "01101001", "01100111", "01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011110", "01011111", "01100001", "01100010", "01100100", 
"01100101", "01100110", "01101000", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", 
"01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101000", "01100110", "01100101", "01100100", 
"01100010", "01100001", "01011111", "01011110", "01011100", "01011010", "01011100", "01011110", "01100000", "01100010", "01100100", "01100111", "01101001", "01101011", "01101101", "01101111", "01110010", "01110100", "01110110", "01110111", 
"01111001", "01111011", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111011", "01111001", "01111000", "01110110", "01110100", "01110011", "01110001", 
"01101111", "01101100", "01101010", "01101000", "01100110", "01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011101", "01011111", "01100001", "01100010", "01100100", "01100101", "01100110", "01100111", 
"01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", 
"01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", 
"01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100010", "01100001", "01011111", "01011101", "01011100", 
"01011010", "01011100", "01011110", "01100000", "01100010", "01100100", "01100110", "01101000", "01101010", "01101100", "01101111", "01110001", "01110011", "01110100", "01110110", "01111000", "01111001", "01111011", "01111100", "01111101", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111011", "01111010", "01111000", "01110111", "01110101", "01110011", "01110010", "01110000", "01101110", "01101100", "01101010", 
"01101000", "01100110", "01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011101", "01011111", "01100000", "01100010", "01100011", "01100100", "01100110", "01100111", "01101000", "01101001", "01101010", 
"01101011", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", 
"01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", 
"01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", 
"01101100", "01101011", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100100", "01100011", "01100010", "01100000", "01011111", "01011101", "01011100", "01011010", "01011100", "01011110", "01100000", "01100010", 
"01100100", "01100110", "01101000", "01101010", "01101100", "01101110", "01110000", "01110010", "01110011", "01110101", "01110111", "01111000", "01111010", "01111011", "01111100", "01111101", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111101", "01111101", "01111011", "01111010", "01111001", "01110111", "01110110", "01110100", "01110010", "01110001", "01101111", "01101101", "01101011", "01101001", "01100111", "01100101", "01100011", 
"01100001", "01011111", "01011101", "01011100", "01011010", "01011100", "01011101", "01011111", "01100000", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", 
"01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", 
"01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", 
"01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101000", 
"01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100000", "01011111", "01011101", "01011100", "01011010", "01011100", "01011101", "01011111", "01100001", "01100011", "01100101", "01100111", "01101001", "01101011", 
"01101101", "01101111", "01110001", "01110010", "01110100", "01110110", "01110111", "01111001", "01111010", "01111011", "01111101", "01111101", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111101", "01111100", "01111011", "01111001", "01111000", "01110111", "01110101", "01110011", "01110010", "01110000", "01101110", "01101100", "01101010", "01101000", "01100111", "01100101", "01100011", "01100001", "01011111", "01011101", 
"01011100", "01011010", "01011011", "01011101", "01011111", "01100000", "01100001", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101101", "01101101", 
"01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", 
"01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", 
"01100001", "01100000", "01011111", "01011101", "01011011", "01011010", "01011100", "01011101", "01011111", "01100001", "01100011", "01100101", "01100111", "01101000", "01101010", "01101100", "01101110", "01110000", "01110010", "01110011", 
"01110101", "01110111", "01111000", "01111001", "01111011", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111010", 
"01111000", "01110111", "01110110", "01110100", "01110010", "01110001", "01101111", "01101101", "01101011", "01101010", "01101000", "01100110", "01100100", "01100010", "01100001", "01011111", "01011101", "01011011", "01011010", "01011011", 
"01011101", "01011110", "01100000", "01100001", "01100010", "01100011", "01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", 
"01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", 
"01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", 
"01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", 
"01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100101", "01100011", "01100010", "01100001", "01100000", "01011110", "01011101", "01011011", 
"01011010", "01011011", "01011101", "01011111", "01100001", "01100010", "01100100", "01100110", "01101000", "01101010", "01101011", "01101101", "01101111", "01110001", "01110010", "01110100", "01110110", "01110111", "01111000", "01111010", 
"01111011", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110110", "01110101", 
"01110011", "01110010", "01110000", "01101110", "01101101", "01101011", "01101001", "01100111", "01100110", "01100100", "01100010", "01100000", "01011111", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01100000", 
"01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", 
"01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", 
"01101010", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011111", "01100000", 
"01100010", "01100100", "01100110", "01100111", "01101001", "01101011", "01101101", "01101110", "01110000", "01110010", "01110011", "01110101", "01110110", "01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110111", "01110101", "01110100", "01110010", "01110001", "01101111", 
"01101110", "01101100", "01101010", "01101001", "01100111", "01100101", "01100100", "01100010", "01100000", "01011111", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01011111", "01100001", "01100010", "01100011", 
"01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", 
"01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01011111", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011111", "01100000", "01100010", "01100100", "01100101", "01100111", "01101001", 
"01101010", "01101100", "01101110", "01101111", "01110001", "01110010", "01110100", "01110101", "01110111", "01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111000", "01110111", "01110110", "01110101", "01110011", "01110010", "01110000", "01101110", "01101101", "01101011", "01101010", 
"01101000", "01100110", "01100101", "01100011", "01100010", "01100000", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01011111", "01100000", "01100010", "01100011", "01100100", "01100101", "01100110", 
"01100110", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", 
"01101111", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100011", "01100010", 
"01100000", "01011111", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01100000", "01100010", "01100011", "01100101", "01100110", "01101000", "01101010", "01101011", "01101101", "01101110", "01110000", 
"01110010", "01110011", "01110101", "01110110", "01110111", "01111000", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111101", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110110", "01110101", "01110100", "01110010", "01110001", "01101111", "01101110", "01101100", "01101011", "01101001", "01101000", "01100110", "01100100", 
"01100011", "01100001", "01100000", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", 
"01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", 
"01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", 
"01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", 
"01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011011", 
"01011010", "01011011", "01011101", "01011110", "01100000", "01100001", "01100011", "01100100", "01100110", "01101000", "01101001", "01101011", "01101100", "01101110", "01101111", "01110001", "01110010", "01110100", "01110101", "01110110", 
"01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", 
"01111010", "01111001", "01111000", "01110111", "01110110", "01110100", "01110011", "01110010", "01110000", "01101111", "01101101", "01101100", "01101010", "01101001", "01100111", "01100110", "01100100", "01100011", "01100001", "01100000", 
"01011110", "01011101", "01011011", "01011010", "01011011", "01011100", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101010", 
"01101010", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", 
"01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", 
"01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", 
"01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011101", "01011110", "01100000", 
"01100001", "01100011", "01100100", "01100110", "01100111", "01101001", "01101010", "01101100", "01101101", "01101111", "01110000", "01110010", "01110011", "01110100", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", 
"01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111100", "01111011", "01111011", "01111010", "01111000", "01110111", 
"01110110", "01110101", "01110100", "01110010", "01110001", "01101111", "01101110", "01101101", "01101011", "01101010", "01101000", "01100111", "01100101", "01100100", "01100010", "01100001", "01011111", "01011110", "01011101", "01011011", 
"01011010", "01011011", "01011100", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", 
"01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", 
"01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100110", 
"01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011101", "01011110", "01011111", "01100001", "01100010", "01100100", "01100101", "01100111", 
"01101000", "01101010", "01101011", "01101101", "01101110", "01101111", "01110001", "01110010", "01110100", "01110101", "01110110", "01110111", "01111000", "01111010", "01111011", "01111011", "01111100", "01111101", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111100", "01111011", "01111010", "01111001", "01111000", "01110111", "01110101", "01110100", "01110011", 
"01110010", "01110000", "01101111", "01101101", "01101100", "01101011", "01101001", "01101000", "01100110", "01100101", "01100011", "01100010", "01100001", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", 
"01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101101", 
"01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", 
"01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", 
"01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", "01011110", "01011111", "01100001", "01100010", "01100011", "01100101", "01100110", "01101000", "01101001", "01101011", "01101100", "01101101", 
"01101111", "01110000", "01110010", "01110011", "01110100", "01110101", "01110111", "01111000", "01111001", "01111010", "01111011", "01111100", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110010", "01110001", "01110000", "01101110", 
"01101101", "01101100", "01101010", "01101001", "01100111", "01100110", "01100101", "01100011", "01100010", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011111", "01100000", 
"01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", 
"01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011101", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011110", "01011111", "01100000", "01100010", "01100011", "01100101", "01100110", "01100111", "01101001", "01101010", "01101100", "01101101", "01101110", "01110000", "01110001", "01110010", "01110100", 
"01110101", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101111", "01101110", "01101100", "01101011", "01101010", 
"01101000", "01100111", "01100110", "01100100", "01100011", "01100010", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", 
"01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", 
"01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", 
"01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", 
"01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011110", "01011111", 
"01100000", "01100010", "01100011", "01100100", "01100110", "01100111", "01101000", "01101010", "01101011", "01101100", "01101110", "01101111", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", 
"01111001", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", 
"01111011", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110011", "01110010", "01110001", "01110000", "01101110", "01101101", "01101100", "01101011", "01101001", "01101000", "01100111", "01100101", 
"01100100", "01100011", "01100001", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", 
"01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", 
"01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", 
"01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", 
"01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", 
"01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", 
"01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011110", "01011111", "01100000", "01100001", "01100011", "01100100", "01100101", 
"01100111", "01101000", "01101001", "01101011", "01101100", "01101101", "01101110", "01110000", "01110001", "01110010", "01110011", "01110101", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111011", "01111100", 
"01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", "01111001", 
"01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101111", "01101110", "01101101", "01101011", "01101010", "01101001", "01101000", "01100110", "01100101", "01100100", "01100010", "01100001", 
"01100000", "01011111", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100111", 
"01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", 
"01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", 
"01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", 
"01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011111", "01100000", "01100001", "01100010", "01100100", "01100101", "01100110", "01101000", "01101001", "01101010", "01101011", 
"01101101", "01101110", "01101111", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111100", "01111100", "01111011", "01111010", "01111001", "01111000", "01111000", "01110111", "01110101", 
"01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101101", "01101100", "01101011", "01101010", "01101000", "01100111", "01100110", "01100101", "01100011", "01100010", "01100001", "01100000", "01011111", "01011101", 
"01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", 
"01101001", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101010", 
"01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011101", "01011111", "01100000", "01100001", "01100010", "01100011", "01100101", "01100110", "01100111", "01101000", "01101010", "01101011", "01101100", "01101101", "01101111", "01110000", "01110001", 
"01110010", "01110011", "01110100", "01110101", "01110111", "01111000", "01111000", "01111001", "01111010", "01111011", "01111100", "01111100", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", 
"01110000", "01101111", "01101110", "01101101", "01101100", "01101010", "01101001", "01101000", "01100111", "01100110", "01100100", "01100011", "01100010", "01100001", "01100000", "01011110", "01011101", "01011100", "01011011", "01011010", 
"01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", 
"01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", 
"01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", 
"01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01100111", 
"01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", 
"01100000", "01100001", "01100010", "01100011", "01100100", "01100110", "01100111", "01101000", "01101001", "01101010", "01101100", "01101101", "01101110", "01101111", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", 
"01110111", "01111000", "01111001", "01111010", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", 
"01101100", "01101011", "01101010", "01101001", "01101000", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", 
"01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", 
"01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", 
"01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", 
"01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", 
"01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100001", "01100010", "01100011", "01100100", 
"01100101", "01100110", "01101000", "01101001", "01101010", "01101011", "01101100", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111001", "01111010", 
"01111011", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111100", "01111100", "01111011", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", 
"01101001", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", 
"01100000", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", 
"01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", 
"01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", 
"01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", 
"01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", "01100000", 
"01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101001", "01101010", 
"01101011", "01101100", "01101101", "01101110", "01101111", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111011", "01111100", "01111100", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", 
"01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101010", "01101001", "01101000", "01100111", "01100110", 
"01100101", "01100100", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", 
"01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", 
"01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", 
"01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", 
"01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101100", "01101101", "01101110", "01101111", 
"01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111001", "01111010", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01110111", 
"01110110", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100100", "01100011", "01100010", 
"01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", 
"01100101", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", 
"01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", 
"01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", 
"01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", 
"01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", 
"01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110001", "01110010", "01110011", "01110100", 
"01110101", "01110110", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110100", 
"01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", 
"01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", 
"01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", 
"01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", 
"01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", 
"01100010", "01100010", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", 
"01100100", "01100101", "01100110", "01100111", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", 
"01111000", "01111001", "01111010", "01111011", "01111011", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", "01111001", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110001", 
"01110000", "01101111", "01101110", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", 
"01011011", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", 
"01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", 
"01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", 
"01011110", "01011101", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", 
"01101001", "01101010", "01101011", "01101100", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110100", "01110101", "01110110", "01110111", "01111000", "01111001", "01111001", "01111010", "01111011", 
"01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111100", "01111100", "01111011", "01111010", "01111010", "01111001", "01111000", "01110111", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", 
"01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", 
"01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", 
"01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", 
"01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", 
"01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", 
"01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111001", "01111010", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", 
"01111011", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", 
"01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", 
"01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", 
"01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", 
"01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", 
"01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", 
"01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", 
"01110011", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111001", 
"01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", 
"01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01100000", 
"01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", 
"01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", 
"01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", 
"01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100010", 
"01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", 
"01110110", "01110111", "01111000", "01111001", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01110111", "01110111", "01110110", 
"01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", 
"01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", 
"01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", 
"01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", 
"01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", 
"01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", 
"01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", 
"01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011111", 
"01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", 
"01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111001", 
"01111010", "01111010", "01111011", "01111011", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", 
"01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", 
"01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", 
"01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", 
"01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", 
"01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", 
"01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", 
"01101101", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111001", "01111000", "01110111", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", 
"01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", 
"01011100", "01011100", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", 
"01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", 
"01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", 
"01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", 
"01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", 
"01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", 
"01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", 
"01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111001", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", 
"01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", 
"01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", 
"01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", 
"01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", 
"01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", 
"01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", 
"01100011", "01100100", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", 
"01110101", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", 
"01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101011", "01101010", 
"01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", 
"01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", 
"01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", 
"01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", 
"01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", 
"01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", 
"01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100110", 
"01100111", "01101000", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", 
"01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111001", "01111000", "01110111", 
"01110111", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01101000", "01100111", 
"01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", 
"01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", 
"01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", 
"01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", 
"01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", 
"01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", 
"01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", 
"01101011", "01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111001", "01111001", "01111010", 
"01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110101", 
"01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", 
"01100011", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", 
"01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", 
"01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", 
"01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", 
"01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", 
"01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", 
"01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", 
"01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100001", 
"01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", 
"01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", 
"01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", 
"01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", 
"01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", 
"01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", 
"01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", 
"01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", 
"01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", 
"01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", 
"01101110", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011111", 
"01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", 
"01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", 
"01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", 
"01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", 
"01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", 
"01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", 
"01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", 
"01110110", "01110111", "01110111", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", 
"01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101100", 
"01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", 
"01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", 
"01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", 
"01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", 
"01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", 
"01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", 
"01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", 
"01111001", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101011", "01101010", "01101010", 
"01101001", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", 
"01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", 
"01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", 
"01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", 
"01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", 
"01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", 
"01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", 
"01011110", "01011110", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101101", 
"01101110", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", 
"01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01110111", "01110111", "01110110", 
"01110110", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", 
"01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", 
"01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", 
"01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110010", "01110010", "01110010", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01110000", 
"01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", 
"01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", 
"01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", 
"01100001", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01110000", "01110000", 
"01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", 
"01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100101", "01100100", 
"01100100", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", 
"01011110", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", 
"01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", 
"01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", 
"01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", 
"01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100100", 
"01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", 
"01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", 
"01110001", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100011", "01100010", 
"01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", 
"01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", 
"01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", 
"01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", 
"01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", 
"01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", 
"01101001", "01101010", "01101010", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", 
"01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", 
"01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101111", 
"01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100000", "01100000", 
"01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", 
"01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", 
"01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", 
"01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", 
"01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", 
"01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", 
"01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", 
"01011101", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", 
"01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", 
"01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", 
"01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", 
"01101011", "01101011", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", 
"01011101", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", 
"01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", 
"01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01110000", 
"01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", 
"01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", 
"01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", 
"01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", 
"01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", 
"01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101010", 
"01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", 
"01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", 
"01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", 
"01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", 
"01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", 
"01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", 
"01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", 
"01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110010", "01110010", 
"01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", 
"01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", 
"01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011010", "01011010", "01011010", 
"01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", 
"01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", 
"01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", 
"01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", 
"01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100111", "01100111", 
"01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", 
"01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", 
"01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", 
"01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", 
"01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", 
"01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", 
"01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", 
"01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101011", 
"01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", 
"01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110001", "01110001", 
"01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", 
"01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", 
"01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", 
"01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", 
"01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", 
"01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", 
"01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", 
"01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", 
"01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", 
"01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", 
"01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", 
"01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", 
"01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", 
"01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", 
"01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", 
"01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", 
"01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", 
"01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", 
"01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", 
"01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100001", 
"01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", 
"01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", 
"01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", 
"01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", 
"01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", 
"01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", 
"01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", 
"01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", 
"01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", 
"01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", 
"01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101110", "01101111", 
"01101110", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", 
"01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", 
"01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", 
"01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110110", 
"01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", 
"01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", 
"01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", 
"01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", 
"01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", 
"01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", 
"01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", 
"01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", 
"01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", 
"01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", 
"01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", 
"01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", 
"01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01110000", 
"01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", 
"01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", 
"01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", 
"01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", 
"01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", 
"01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", 
"01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", 
"01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", 
"01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", 
"01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", 
"01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", 
"01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", 
"01101101", "01101101", "01101101", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", 
"01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", 
"01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", 
"01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", 
"01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", 
"01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", 
"01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", 
"01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", 
"01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", 
"01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", 
"01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", 
"01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", 
"01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", 
"01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", 
"01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", 
"01101001", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", 
"01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", 
"01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", 
"01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101111", 
"01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", 
"01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", 
"01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", 
"01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", 
"01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", 
"01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", 
"01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", 
"01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", 
"01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", 
"01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110001", 
"01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", 
"01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100110", 
"01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", 
"01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", 
"01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101001", "01101010", 
"01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101001", 
"01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", 
"01101001", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", 
"01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", 
"01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100100", 
"01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", 
"01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", 
"01101011", "01101011", "01101011", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", 
"01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", 
"01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", 
"01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", 
"01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", 
"01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", 
"01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", 
"01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", 
"01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", 
"01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", 
"01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101110", 
"01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", 
"01111001", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101100", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", 
"01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101010", "01101010", "01101010", "01101010", 
"01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", 
"01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110000", 
"01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", 
"01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", 
"01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", 
"01101000", "01100111", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", 
"01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", 
"01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111100", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", 
"01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", 
"01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", 
"01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", 
"01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", 
"01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", 
"01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", 
"01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", 
"01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", 
"01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", 
"01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", 
"01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011011", 
"01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", 
"01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", 
"01101001", "01101001", "01101001", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", 
"01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", 
"01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", 
"01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", 
"01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", 
"01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", 
"01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", 
"01100100", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", 
"01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", 
"01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", 
"01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", 
"01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", 
"01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", 
"01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", 
"01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", 
"01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", 
"01100100", "01100101", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", "01101000", "01101000", "01101000", "01101000", 
"01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", 
"01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", 
"01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", 
"01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", 
"01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", 
"01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100111", "01100110", "01100110", 
"01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", 
"01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", 
"01101010", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", 
"01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", 
"01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", 
"01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", 
"01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", 
"01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", 
"01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", 
"01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", 
"01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", 
"01100111", "01100111", "01100111", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", 
"01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", 
"01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", 
"01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", 
"01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", 
"01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", 
"01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", 
"01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", 
"01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100110", 
"01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", 
"01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", 
"01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", 
"01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", 
"01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", 
"01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100110", "01100111", "01100110", "01100110", "01100110", "01100110", 
"01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", 
"01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", 
"01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", 
"01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", 
"01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", 
"01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", 
"01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", 
"01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", 
"01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", 
"01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", 
"01100100", "01100100", "01100101", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", 
"01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", 
"01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", 
"01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", 
"01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", 
"01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", 
"01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", 
"01100101", "01100101", "01100101", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", 
"01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", 
"01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", 
"01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", 
"01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", 
"01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", 
"01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", 
"01101000", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", 
"01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", 
"01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", 
"01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", 
"01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", 
"01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", 
"01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", 
"01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", 
"01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", 
"01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", 
"01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100100", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", 
"01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", 
"01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", 
"01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", 
"01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", 
"01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", 
"01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", 
"01100010", "01100010", "01100011", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", 
"01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", 
"01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", 
"01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", 
"01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", 
"01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", 
"01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", 
"01100011", "01100011", "01100011", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", 
"01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", 
"01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", 
"01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", 
"01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", 
"01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", 
"01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", 
"01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", 
"01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", 
"01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", 
"01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", 
"01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", 
"01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", 
"01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", 
"01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", 
"01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", 
"01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", 
"01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", 
"01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", 
"01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", 
"01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", 
"01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", 
"01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", 
"01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", 
"01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", 
"01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", 
"01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", 
"01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", 
"01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", 
"01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", 
"01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100001", "01100001", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", 
"01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", 
"01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", 
"01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", 
"01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", 
"01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", 
"01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", 
"01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", 
"01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", 
"01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", 
"01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", 
"01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", 
"01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", 
"01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", 
"01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", 
"01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", 
"01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", 
"01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", 
"01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", 
"01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", 
"01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", 
"01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", 
"01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", 
"01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", 
"01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", 
"01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", 
"01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", 
"01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", 
"01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", 
"01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", 
"01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", 
"01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", 
"01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", 
"01011111", "01011111", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", 
"01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", 
"01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", 
"01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", 
"01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", 
"01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", 
"01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", 
"01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", 
"01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", 
"01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", 
"01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", 
"01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", 
"01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01011111", "01011111", "01011110", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", 
"01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", 
"01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", 
"01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", 
"01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", 
"01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", 
"01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", 
"01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", 
"01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", 
"01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", 
"01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", 
"01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", 
"01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", 
"01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", 
"01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", 
"01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", 
"01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", 
"01011101", "01011101", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", 
"01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", 
"01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", 
"01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", 
"01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", 
"01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", 
"01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", 
"01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", 
"01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", 
"01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", 
"01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011101", "01011101", "01011100", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", 
"01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", 
"01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", 
"01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", 
"01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", 
"01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", 
"01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", 
"01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", 
"01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", 
"01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", 
"01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", 
"01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", 
"01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", 
"01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", 
"01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", 
"01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", 
"01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", 
"01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", 
"01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", 
"01011011", "01011100", "01011100", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", 
"01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", 
"01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", 
"01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", 
"01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", 
"01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", 
"01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", 
"01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", 
"01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", 
"01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", 
"01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", 
"01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", 
"01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", 
"01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", 
"01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", 
"01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", 
"01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", 
"01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", 
"01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", 
"01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", 
"01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", 
"01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", 
"01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", 
"01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", 
"01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", 
"01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", 
"01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", 
"01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", 
"01011010", "01011010", "01011010", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", 
"01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", 
"01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", 
"01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", 
"01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", 
"01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", 
"01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", 
"01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", 
"01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110111", 
"01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", 
"01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", 
"01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", 
"01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", 
"01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", 
"01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", 
"01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", 
"01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", 
"01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", 
"01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", 
"01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", 
"01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", 
"01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", 
"01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", 
"01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", 
"01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", 
"01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", 
"01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", 
"01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", 
"01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", 
"01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", 
"01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", 
"01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", 
"01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", 
"01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", 
"01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", 
"01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", 
"01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", 
"01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", 
"01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", 
"01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", 
"01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", 
"01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", 
"01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", 
"01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", 
"01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", 
"01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", 
"01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", 
"01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", 
"01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", 
"01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", 
"01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", 
"01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011100", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", 
"01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", 
"01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", 
"01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", 
"01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", 
"01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", 
"01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", 
"01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", 
"01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", 
"01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", 
"01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", 
"01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", 
"01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011101", "01011101", "01011100", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", 
"01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", 
"01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", 
"01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", 
"01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", 
"01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", 
"01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", 
"01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", 
"01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", 
"01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", 
"01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", 
"01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", 
"01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", 
"01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", 
"01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", 
"01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", 
"01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", 
"01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", 
"01011101", "01011110", "01011110", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", 
"01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", 
"01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", 
"01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", 
"01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", 
"01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", 
"01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", 
"01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", 
"01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", 
"01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", 
"01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", 
"01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01011111", "01011111", "01011110", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", 
"01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", 
"01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", 
"01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", 
"01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", 
"01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", 
"01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", 
"01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", 
"01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", 
"01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", 
"01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", 
"01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", 
"01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", 
"01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", 
"01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", 
"01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", 
"01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", 
"01011111", "01100000", "01100000", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", 
"01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", 
"01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", 
"01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", 
"01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", 
"01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", 
"01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", 
"01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", 
"01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", 
"01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", 
"01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", 
"01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", 
"01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", 
"01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", 
"01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", 
"01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", 
"01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", 
"01011110", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", 
"01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", 
"01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", 
"01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", 
"01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", 
"01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", 
"01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", 
"01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", 
"01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", 
"01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", 
"01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", 
"01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", 
"01100001", "01100010", "01100010", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", 
"01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", 
"01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", 
"01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", 
"01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", 
"01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", 
"01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", 
"01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", 
"01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", 
"01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", 
"01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", 
"01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", 
"01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", 
"01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", 
"01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", 
"01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", 
"01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", 
"01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", 
"01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", 
"01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", 
"01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", 
"01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", 
"01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", 
"01011111", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", 
"01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", 
"01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", 
"01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", 
"01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", 
"01100011", "01100011", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", 
"01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", 
"01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", 
"01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", 
"01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", 
"01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", 
"01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100100", 
"01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", 
"01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", 
"01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", 
"01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", 
"01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", 
"01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", 
"01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", 
"01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", 
"01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", 
"01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", 
"01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", 
"01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", 
"01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", 
"01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", 
"01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", 
"01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", 
"01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", 
"01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", 
"01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", 
"01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", 
"01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", 
"01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", 
"01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", 
"01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", 
"01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", 
"01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", 
"01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", 
"01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", 
"01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", 
"01100101", "01100101", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", 
"01100000", "01100000", "01100000", "01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", 
"01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", 
"01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", 
"01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", 
"01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", 
"01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100110", 
"01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", 
"01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", 
"01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", 
"01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", 
"01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", 
"01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", 
"01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100110", "01100111", "01100110", "01100110", "01100110", "01100110", 
"01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", 
"01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", 
"01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", 
"01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", 
"01100100", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", 
"01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", 
"01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", 
"01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", 
"01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100101", "01100100", "01100100", 
"01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", 
"01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", 
"01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", 
"01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", 
"01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01100111", 
"01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", 
"01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100110", "01100111", 
"01100111", "01100111", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", 
"01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", 
"01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", 
"01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", 
"01101110", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", 
"01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", 
"01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", 
"01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", 
"01101000", "01101000", "01100111", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", 
"01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", 
"01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", 
"01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", 
"01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", 
"01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", 
"01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", 
"01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", 
"01100100", "01100101", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", "01101000", "01101000", "01101000", "01101000", 
"01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", 
"01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", 
"01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101011", 
"01101010", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", 
"01100110", "01100110", "01100111", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", 
"01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", 
"01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", 
"01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01011111", "01100000", "01100000", 
"01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", 
"01101000", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", 
"01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", 
"01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", 
"01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", 
"01110000", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", 
"01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", 
"01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", 
"01101001", "01101001", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", 
"01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", 
"01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", 
"01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", 
"01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", 
"01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", 
"01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100011", 
"01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", 
"01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", 
"01101010", "01101010", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", 
"01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", 
"01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", 
"01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", 
"01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101100", 
"01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01011111", "01100000", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", 
"01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101010", "01101010", "01101010", "01101010", 
"01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", 
"01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110000", 
"01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", 
"01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", 
"01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", 
"01101000", "01101000", "01101001", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", 
"01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", 
"01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", 
"01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", 
"01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", 
"01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", 
"01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", 
"01110001", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", 
"01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", 
"01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", 
"01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", 
"01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", 
"01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", 
"01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", 
"01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", 
"01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", 
"01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", 
"01101011", "01101011", "01101011", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", 
"01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", 
"01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", 
"01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", 
"01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101101", 
"01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", 
"01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", 
"01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100111", 
"01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011111", 
"01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", 
"01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", 
"01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", 
"01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", 
"01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", 
"01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", 
"01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100000", "01100001", 
"01100001", "01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", 
"01101001", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", 
"01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", 
"01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", 
"01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", 
"01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101111", 
"01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", 
"01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", 
"01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", 
"01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", 
"01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", 
"01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", 
"01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", 
"01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", 
"01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", 
"01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", 
"01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", 
"01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", 
"01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", 
"01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100100", 
"01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", 
"01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", 
"01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", 
"01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", 
"01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", 
"01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", 
"01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", 
"01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", 
"01101101", "01101101", "01101101", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", 
"01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", 
"01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", 
"01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", 
"01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", 
"01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", 
"01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", 
"01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", 
"01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", 
"01100010", "01100010", "01100011", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", 
"01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", 
"01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", 
"01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", 
"01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", 
"01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", 
"01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100011", 
"01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", 
"01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", 
"01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", 
"01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", 
"01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", 
"01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110010", 
"01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", 
"01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", 
"01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", 
"01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101110", "01101111", "01101110", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", 
"01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", 
"01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", 
"01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", 
"01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", 
"01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", 
"01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", 
"01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", 
"01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", 
"01100000", "01100000", "01100001", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", 
"01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", 
"01101110", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", 
"01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", 
"01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", 
"01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", 
"01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", 
"01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", 
"01111000", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", 
"01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", 
"01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", 
"01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", 
"01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", 
"01101111", "01101111", "01101111", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", 
"01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", 
"01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", 
"01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", 
"01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", 
"01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", 
"01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", 
"01101000", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", 
"01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", 
"01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", 
"01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", 
"01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", 
"01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", 
"01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01101000", "01101000", 
"01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110110", 
"01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", 
"01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", 
"01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", 
"01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", 
"01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", 
"01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", 
"01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101011", 
"01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", 
"01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", 
"01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", 
"01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", 
"01100000", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", 
"01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", 
"01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", 
"01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", 
"01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", 
"01101110", "01101110", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", 
"01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", 
"01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011111", "01011110", 
"01011101", "01011101", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", 
"01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", 
"01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", 
"01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", 
"01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", 
"01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", 
"01011111", "01011111", "01011110", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", 
"01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", 
"01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", 
"01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110001", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", 
"01101000", "01101000", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011010", 
"01011010", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100100", 
"01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", 
"01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", 
"01110001", "01110001", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", 
"01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", 
"01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", 
"01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011010", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", 
"01100100", "01100101", "01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110001", "01110001", "01110010", 
"01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", 
"01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100110", 
"01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011010", "01011011", "01011100", "01011100", 
"01011101", "01011110", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100101", "01100110", "01100110", "01100111", 
"01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", 
"01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", 
"01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", 
"01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011110", "01011101", "01011100", 
"01011100", "01011011", "01011010", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100110", 
"01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", 
"01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", 
"01110001", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100011", "01100010", 
"01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01100000", 
"01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", 
"01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", 
"01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", 
"01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", 
"01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", 
"01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100011", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", 
"01101001", "01101010", "01101010", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110001", "01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", 
"01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", 
"01111010", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", 
"01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", 
"01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100010", 
"01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", 
"01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", 
"01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", 
"01110001", "01110000", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", 
"01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", 
"01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", 
"01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101011", 
"01101100", "01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", 
"01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", 
"01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", 
"01101001", "01101001", "01101000", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", 
"01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", 
"01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101100", 
"01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", 
"01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101100", "01101011", 
"01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100101", "01100100", "01100100", "01100011", 
"01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", 
"01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101101", "01101101", 
"01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", 
"01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110111", "01110110", 
"01110101", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", "01100110", 
"01100110", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", 
"01011101", "01011110", "01011111", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100110", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", 
"01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", 
"01110000", "01101111", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", 
"01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", 
"01100001", "01100000", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", 
"01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", 
"01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110011", 
"01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100011", 
"01100010", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", 
"01100001", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101001", 
"01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", 
"01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", 
"01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", 
"01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", 
"01011111", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", 
"01100011", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110011", 
"01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01110111", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", 
"01101110", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011111", 
"01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", 
"01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", 
"01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", 
"01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101001", 
"01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", 
"01011101", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", 
"01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", 
"01110110", "01110111", "01110111", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", 
"01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", 
"01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", 
"01011010", "01011011", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", 
"01100110", "01100111", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", 
"01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", 
"01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", 
"01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011101", "01011100", 
"01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01101000", 
"01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110011", "01110100", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", 
"01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", 
"01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", 
"01100110", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", 
"01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", 
"01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", 
"01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", 
"01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", 
"01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", 
"01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", 
"01011011", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", 
"01101100", "01101101", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", 
"01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111001", "01111000", "01110111", "01110111", "01110110", "01110101", "01110100", 
"01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", 
"01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", 
"01100001", "01100010", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", 
"01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", 
"01110001", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", 
"01110100", "01110100", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", 
"01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", 
"01100100", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", 
"01011101", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", 
"01101111", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111001", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", 
"01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", 
"01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100011", 
"01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", 
"01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", 
"01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", 
"01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", 
"01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011111", 
"01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", 
"01110010", "01110010", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", 
"01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", 
"01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", 
"01011010", "01011011", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", 
"01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", 
"01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", 
"01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", 
"01100001", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", 
"01100011", "01100100", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", 
"01110101", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", 
"01111001", "01111000", "01110111", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", 
"01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011011", "01011011", "01011100", "01011101", 
"01011110", "01011111", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", 
"01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", 
"01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", 
"01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", 
"01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", 
"01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", 
"01011111", "01011111", "01011110", "01011101", "01011100", "01011011", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", 
"01100110", "01100111", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", 
"01110111", "01111000", "01111001", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", 
"01110101", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", 
"01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", 
"01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", 
"01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", 
"01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", 
"01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", 
"01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", 
"01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011111", "01011110", 
"01011101", "01011100", "01011100", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", 
"01101001", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", 
"01111010", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01110111", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", 
"01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", 
"01011110", "01011101", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100011", "01100100", 
"01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", 
"01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", 
"01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", 
"01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", 
"01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011100", 
"01011011", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", 
"01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", 
"01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111001", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", 
"01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011110", "01011101", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011100", "01011101", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", 
"01101000", "01101000", "01101001", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", 
"01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", 
"01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", 
"01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101001", "01101000", "01101000", "01100111", 
"01100111", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011011", 
"01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", 
"01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111001", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", 
"01111011", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", 
"01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011100", "01011101", 
"01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", 
"01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", 
"01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", 
"01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", 
"01100101", "01100100", "01100100", "01100011", "01100011", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011100", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", 
"01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", 
"01110011", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", "01111010", "01111001", "01111000", 
"01110111", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", 
"01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100001", "01100001", 
"01100010", "01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", 
"01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", 
"01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", 
"01100011", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", 
"01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", 
"01110110", "01110111", "01110111", "01111000", "01111001", "01111010", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", "01111001", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", 
"01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", 
"01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011101", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", 
"01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", 
"01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", 
"01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", 
"01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", 
"01101100", "01101100", "01101011", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100100", "01100011", "01100010", 
"01100001", "01100001", "01100000", "01011111", "01011110", "01011101", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", 
"01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110100", "01110101", "01110110", "01110111", "01111000", 
"01111001", "01111001", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", 
"01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011101", "01011110", "01011110", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01100111", "01101000", 
"01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", 
"01110000", "01110001", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", 
"01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", 
"01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", 
"01011111", "01011110", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", 
"01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111011", 
"01111011", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", 
"01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01101111", "01101110", "01101101", "01101100", "01101011", 
"01101010", "01101001", "01101000", "01100111", "01100110", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", 
"01011110", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", 
"01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", 
"01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011110", "01011110", 
"01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", 
"01101100", "01101101", "01101110", "01101111", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", 
"01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101010", "01101001", "01101000", "01100111", "01100110", 
"01100101", "01100100", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01011111", "01100000", "01100001", "01100010", 
"01100011", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", 
"01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", 
"01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", 
"01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110000", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", 
"01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100011", "01100010", "01100001", "01100000", "01011111", "01011111", "01011110", "01011101", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101100", "01101101", "01101110", "01101111", 
"01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111001", "01111010", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", "01111001", "01111000", "01111000", "01110111", 
"01110110", "01110101", "01110100", "01110011", "01110010", "01110001", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100000", 
"01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100000", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", 
"01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", 
"01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", 
"01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", 
"01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", 
"01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", 
"01100111", "01100111", "01100110", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", 
"01011101", "01011110", "01011111", "01100000", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110001", "01110010", "01110011", 
"01110100", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", 
"01110001", "01110000", "01101111", "01101110", "01101100", "01101011", "01101010", "01101001", "01101000", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01011111", "01011110", "01011101", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", 
"01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", 
"01101111", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", 
"01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", 
"01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01101000", "01101001", "01101010", "01101011", "01101100", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", 
"01110111", "01111000", "01111001", "01111010", "01111011", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101111", "01101110", "01101101", 
"01101100", "01101010", "01101001", "01101000", "01100111", "01100110", "01100100", "01100011", "01100010", "01100001", "01100000", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", 
"01011111", "01100000", "01100001", "01100010", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", 
"01101100", "01101101", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", 
"01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", 
"01101111", "01101110", "01101110", "01101101", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", 
"01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01100000", "01100001", "01100010", "01100011", 
"01100100", "01100110", "01100111", "01101000", "01101001", "01101010", "01101100", "01101101", "01101110", "01101111", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111001", "01111010", 
"01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111100", 
"01111100", "01111011", "01111010", "01111001", "01111000", "01111000", "01110111", "01110101", "01110100", "01110011", "01110010", "01110001", "01110000", "01101111", "01101101", "01101100", "01101011", "01101010", "01101000", "01100111", 
"01100110", "01100101", "01100011", "01100010", "01100001", "01100000", "01011111", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", 
"01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", 
"01101111", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", 
"01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", 
"01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", 
"01101110", "01101101", "01101101", "01101100", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100011", "01100011", 
"01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011111", "01100000", "01100001", "01100010", "01100011", "01100101", "01100110", "01100111", 
"01101000", "01101010", "01101011", "01101100", "01101101", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110111", "01111000", "01111000", "01111001", "01111010", "01111011", "01111100", "01111100", 
"01111101", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111100", "01111011", "01111010", "01111001", 
"01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101111", "01101110", "01101101", "01101011", "01101010", "01101001", "01101000", "01100110", "01100101", "01100100", "01100010", "01100001", 
"01100000", "01011111", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100111", 
"01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", 
"01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", 
"01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", 
"01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", 
"01011111", "01011110", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011111", "01100000", "01100001", "01100010", "01100100", "01100101", "01100110", "01101000", "01101001", "01101010", "01101011", 
"01101101", "01101110", "01101111", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111100", "01111100", "01111101", "01111101", "01111110", "01111110", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", 
"01110011", "01110010", "01110001", "01110000", "01101110", "01101101", "01101100", "01101011", "01101001", "01101000", "01100111", "01100101", "01100100", "01100011", "01100001", "01100000", "01011111", "01011110", "01011100", "01011011", 
"01011010", "01011011", "01011100", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", 
"01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", 
"01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110100", "01110011", 
"01110011", "01110011", "01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", 
"01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", 
"01011100", "01011011", "01011010", "01011011", "01011100", "01011110", "01011111", "01100000", "01100001", "01100011", "01100100", "01100101", "01100111", "01101000", "01101001", "01101011", "01101100", "01101101", "01101110", "01110000", 
"01110001", "01110010", "01110011", "01110101", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101111", 
"01101110", "01101100", "01101011", "01101010", "01101000", "01100111", "01100110", "01100100", "01100011", "01100010", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011110", 
"01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101000", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", 
"01101101", "01101110", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", 
"01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", 
"01110010", "01110010", "01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", 
"01101010", "01101010", "01101001", "01101000", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011101", "01011100", "01011011", "01011010", 
"01011011", "01011100", "01011110", "01011111", "01100000", "01100010", "01100011", "01100100", "01100110", "01100111", "01101000", "01101010", "01101011", "01101100", "01101110", "01101111", "01110000", "01110010", "01110011", "01110100", 
"01110101", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110101", "01110100", "01110010", "01110001", "01110000", "01101110", "01101101", "01101100", "01101010", "01101001", 
"01100111", "01100110", "01100101", "01100011", "01100010", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", "01011101", "01011111", "01100000", "01100001", "01100010", "01100010", "01100011", 
"01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01101111", 
"01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", 
"01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", 
"01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", 
"01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100010", "01100001", "01100000", "01011111", "01011101", "01011100", "01011011", "01011010", "01011011", "01011100", "01011110", 
"01011111", "01100000", "01100010", "01100011", "01100101", "01100110", "01100111", "01101001", "01101010", "01101100", "01101101", "01101110", "01110000", "01110001", "01110010", "01110100", "01110101", "01110110", "01110111", "01111000", 
"01111001", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111100", 
"01111011", "01111010", "01111001", "01111000", "01110111", "01110101", "01110100", "01110011", "01110010", "01110000", "01101111", "01101101", "01101100", "01101011", "01101001", "01101000", "01100110", "01100101", "01100011", "01100010", 
"01100001", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100100", "01100101", "01100110", "01100111", "01101000", 
"01101000", "01101001", "01101010", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110011", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", 
"01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101010", "01101001", "01101000", "01101000", 
"01100111", "01100110", "01100101", "01100100", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011100", "01011110", "01011111", "01100001", "01100010", 
"01100011", "01100101", "01100110", "01101000", "01101001", "01101011", "01101100", "01101101", "01101111", "01110000", "01110010", "01110011", "01110100", "01110101", "01110111", "01111000", "01111001", "01111010", "01111011", "01111100", 
"01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111101", "01111100", "01111011", "01111011", "01111010", "01111000", "01110111", 
"01110110", "01110101", "01110100", "01110010", "01110001", "01101111", "01101110", "01101101", "01101011", "01101010", "01101000", "01100111", "01100101", "01100100", "01100010", "01100001", "01011111", "01011110", "01011101", "01011011", 
"01011010", "01011011", "01011100", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", 
"01101100", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110011", 
"01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", 
"01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100110", 
"01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011101", "01011110", "01011111", "01100001", "01100010", "01100100", "01100101", "01100111", 
"01101000", "01101010", "01101011", "01101101", "01101110", "01101111", "01110001", "01110010", "01110100", "01110101", "01110110", "01110111", "01111000", "01111010", "01111011", "01111011", "01111100", "01111101", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110100", "01110011", "01110010", 
"01110000", "01101111", "01101101", "01101100", "01101010", "01101001", "01100111", "01100110", "01100100", "01100011", "01100001", "01100000", "01011110", "01011101", "01011011", "01011010", "01011011", "01011100", "01011110", "01011111", 
"01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101110", 
"01101111", "01101111", "01110000", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", 
"01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", 
"01110110", "01110101", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", 
"01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", "01100111", "01100110", "01100101", "01100100", "01100011", 
"01100010", "01100001", "01100000", "01011111", "01011110", "01011100", "01011011", "01011010", "01011011", "01011101", "01011110", "01100000", "01100001", "01100011", "01100100", "01100110", "01100111", "01101001", "01101010", "01101100", 
"01101101", "01101111", "01110000", "01110010", "01110011", "01110100", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111101", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110110", "01110101", "01110100", "01110010", "01110001", "01101111", "01101110", "01101100", "01101011", 
"01101001", "01101000", "01100110", "01100100", "01100011", "01100001", "01100000", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01011111", "01100000", "01100001", "01100010", "01100011", "01100100", 
"01100101", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110000", "01110001", 
"01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", 
"01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01110000", "01101111", 
"01101111", "01101110", "01101110", "01101101", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", 
"01011111", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01100000", "01100001", "01100011", "01100100", "01100110", "01101000", "01101001", "01101011", "01101100", "01101110", "01101111", "01110001", 
"01110010", "01110100", "01110101", "01110110", "01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", 
"01111101", "01111101", "01111100", "01111011", "01111010", "01111000", "01110111", "01110110", "01110101", "01110011", "01110010", "01110000", "01101110", "01101101", "01101011", "01101010", "01101000", "01100110", "01100101", "01100011", 
"01100010", "01100000", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01011111", "01100000", "01100010", "01100011", "01100100", "01100101", "01100110", "01100110", "01100111", "01101000", "01101001", 
"01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", 
"01110011", "01110100", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", 
"01110101", "01110101", "01110100", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101111", "01101110", 
"01101101", "01101101", "01101100", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", "01100110", "01100110", "01100101", "01100100", "01100011", "01100010", "01100000", "01011111", "01011110", "01011101", 
"01011011", "01011010", "01011011", "01011101", "01011110", "01100000", "01100010", "01100011", "01100101", "01100110", "01101000", "01101010", "01101011", "01101101", "01101110", "01110000", "01110010", "01110011", "01110101", "01110110", 
"01110111", "01111000", "01111010", "01111011", "01111100", "01111101", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111010", 
"01111001", "01111000", "01110111", "01110101", "01110100", "01110010", "01110001", "01101111", "01101110", "01101100", "01101010", "01101001", "01100111", "01100101", "01100100", "01100010", "01100000", "01011111", "01011101", "01011011", 
"01011010", "01011011", "01011101", "01011110", "01011111", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", 
"01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", 
"01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", 
"01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101101", 
"01101100", "01101011", "01101011", "01101010", "01101001", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01011111", "01011110", "01011101", "01011011", "01011010", "01011011", 
"01011101", "01011111", "01100000", "01100010", "01100100", "01100101", "01100111", "01101001", "01101010", "01101100", "01101110", "01101111", "01110001", "01110010", "01110100", "01110101", "01110111", "01111000", "01111001", "01111010", 
"01111011", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111010", "01111001", "01111000", "01110110", "01110101", 
"01110011", "01110010", "01110000", "01101110", "01101101", "01101011", "01101001", "01100111", "01100110", "01100100", "01100010", "01100000", "01011111", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01100000", 
"01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", 
"01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", 
"01101010", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100011", "01100010", "01100001", "01100000", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011111", "01100000", 
"01100010", "01100100", "01100110", "01100111", "01101001", "01101011", "01101101", "01101110", "01110000", "01110010", "01110011", "01110101", "01110110", "01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111010", "01111000", "01110111", "01110110", "01110100", "01110010", "01110001", "01101111", "01101101", 
"01101011", "01101010", "01101000", "01100110", "01100100", "01100010", "01100001", "01011111", "01011101", "01011011", "01011010", "01011011", "01011101", "01011110", "01100000", "01100001", "01100010", "01100011", "01100101", "01100110", 
"01100111", "01101000", "01101000", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", 
"01110011", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", 
"01110011", "01110011", "01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", 
"01101000", "01101000", "01100111", "01100110", "01100101", "01100011", "01100010", "01100001", "01100000", "01011110", "01011101", "01011011", "01011010", "01011011", "01011101", "01011111", "01100001", "01100010", "01100100", "01100110", 
"01101000", "01101010", "01101011", "01101101", "01101111", "01110001", "01110010", "01110100", "01110110", "01110111", "01111000", "01111010", "01111011", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111001", "01111000", "01110111", "01110101", "01110011", "01110010", "01110000", "01101110", "01101100", "01101010", "01101000", "01100111", "01100101", 
"01100011", "01100001", "01011111", "01011101", "01011100", "01011010", "01011011", "01011101", "01011111", "01100000", "01100001", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101010", 
"01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", 
"01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", 
"01110011", "01110010", "01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101010", "01101001", "01101000", "01100111", 
"01100110", "01100101", "01100100", "01100011", "01100001", "01100000", "01011111", "01011101", "01011011", "01011010", "01011100", "01011101", "01011111", "01100001", "01100011", "01100101", "01100111", "01101000", "01101010", "01101100", 
"01101110", "01110000", "01110010", "01110011", "01110101", "01110111", "01111000", "01111001", "01111011", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111101", 
"01111101", "01111011", "01111010", "01111001", "01110111", "01110110", "01110100", "01110010", "01110001", "01101111", "01101101", "01101011", "01101001", "01100111", "01100101", "01100011", "01100001", "01011111", "01011101", "01011100", 
"01011010", "01011100", "01011101", "01011111", "01100000", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101100", "01101101", "01101110", "01101110", 
"01101111", "01110000", "01110000", "01110001", "01110001", "01110010", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", 
"01110111", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", 
"01110010", "01110010", "01110001", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", 
"01100011", "01100010", "01100000", "01011111", "01011101", "01011100", "01011010", "01011100", "01011101", "01011111", "01100001", "01100011", "01100101", "01100111", "01101001", "01101011", "01101101", "01101111", "01110001", "01110010", 
"01110100", "01110110", "01110111", "01111001", "01111010", "01111011", "01111101", "01111101", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111011", "01111010", "01111000", 
"01110111", "01110101", "01110011", "01110010", "01110000", "01101110", "01101100", "01101010", "01101000", "01100110", "01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011101", "01011111", "01100000", 
"01100010", "01100011", "01100100", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", 
"01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01111000", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110010", 
"01110001", "01110001", "01110000", "01101111", "01101111", "01101110", "01101110", "01101101", "01101100", "01101011", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100100", "01100011", "01100010", "01100000", 
"01011111", "01011101", "01011100", "01011010", "01011100", "01011110", "01100000", "01100010", "01100100", "01100110", "01101000", "01101010", "01101100", "01101110", "01110000", "01110010", "01110011", "01110101", "01110111", "01111000", 
"01111010", "01111011", "01111100", "01111101", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111011", "01111001", "01111000", "01110110", "01110100", "01110011", "01110001", 
"01101111", "01101100", "01101010", "01101000", "01100110", "01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011101", "01011111", "01100001", "01100010", "01100100", "01100101", "01100110", "01100111", 
"01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", 
"01110101", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", 
"01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01111000", 
"01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", 
"01110000", "01101111", "01101111", "01101110", "01101101", "01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100101", "01100100", "01100010", "01100001", "01011111", "01011101", "01011100", 
"01011010", "01011100", "01011110", "01100000", "01100010", "01100100", "01100110", "01101000", "01101010", "01101100", "01101111", "01110001", "01110011", "01110100", "01110110", "01111000", "01111001", "01111011", "01111100", "01111101", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", "01111100", "01111011", "01111001", "01110111", "01110110", "01110100", "01110010", "01101111", "01101101", "01101011", "01101001", "01100111", 
"01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011110", "01011111", "01100001", "01100010", "01100100", "01100101", "01100110", "01101000", "01101001", "01101010", "01101011", "01101100", "01101100", 
"01101101", "01101110", "01101111", "01101111", "01110000", "01110001", "01110001", "01110010", "01110010", "01110011", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", 
"01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", 
"01110111", "01110111", "01110110", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110011", "01110010", "01110010", "01110001", "01110001", "01110000", "01101111", 
"01101111", "01101110", "01101101", "01101100", "01101100", "01101011", "01101010", "01101001", "01101000", "01100110", "01100101", "01100100", "01100010", "01100001", "01011111", "01011110", "01011100", "01011010", "01011100", "01011110", 
"01100000", "01100010", "01100100", "01100111", "01101001", "01101011", "01101101", "01101111", "01110010", "01110100", "01110110", "01110111", "01111001", "01111011", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111101", "01111100", "01111010", "01111000", "01110111", "01110101", "01110011", "01110001", "01101110", "01101100", "01101010", "01100111", "01100101", "01100011", "01100000", "01011110", "01011100", 
"01011010", "01011100", "01011110", "01100000", "01100001", "01100011", "01100100", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011", "01101100", "01101101", "01101110", "01101110", "01101111", "01110000", "01110000", 
"01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", 
"01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", 
"01110111", "01110110", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101110", 
"01101101", "01101100", "01101011", "01101010", "01101001", "01101000", "01100111", "01100110", "01100100", "01100011", "01100001", "01100000", "01011110", "01011100", "01011010", "01011100", "01011110", "01100000", "01100011", "01100101", 
"01100111", "01101010", "01101100", "01101110", "01110001", "01110011", "01110101", "01110111", "01111000", "01111010", "01111100", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111110", "01111110", "01111101", 
"01111011", "01111010", "01111000", "01110110", "01110100", "01110010", "01101111", "01101101", "01101010", "01101000", "01100110", "01100011", "01100001", "01011110", "01011100", "01011010", "01011100", "01011110", "01100000", "01100010", 
"01100011", "01100101", "01100110", "01100111", "01101001", "01101010", "01101011", "01101100", "01101101", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", 
"01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", 
"01110110", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101101", "01101100", 
"01101011", "01101010", "01101001", "01100111", "01100110", "01100101", "01100011", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011110", "01100001", "01100011", "01100110", "01101000", "01101010", "01101101", 
"01101111", "01110010", "01110100", "01110110", "01111000", "01111010", "01111011", "01111101", "01111110", "01111110", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111011", "01111001", "01110111", "01110101", 
"01110011", "01110000", "01101110", "01101011", "01101001", "01100110", "01100100", "01100001", "01011111", "01011100", "01011010", "01011100", "01011110", "01100000", "01100010", "01100100", "01100101", "01100111", "01101000", "01101001", 
"01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", "01110110", 
"01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", 
"01110110", "01110101", "01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101001", 
"01101000", "01100111", "01100101", "01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011111", "01100001", "01100100", "01100110", "01101001", "01101011", "01101110", "01110000", "01110011", "01110101", 
"01110111", "01111001", "01111011", "01111100", "01111101", "01111110", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111010", "01111000", "01110110", "01110100", "01110010", "01101111", "01101100", "01101010", 
"01100111", "01100100", "01100010", "01011111", "01011100", "01011010", "01011100", "01011110", "01100000", "01100010", "01100100", "01100110", "01100111", "01101000", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", 
"01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01110111", "01111000", "01111000", 
"01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", 
"01110101", "01110101", "01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101000", "01100111", "01100110", 
"01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011100", "01011111", "01100010", "01100100", "01100111", "01101010", "01101100", "01101111", "01110010", "01110100", "01110110", "01111000", "01111010", "01111100", 
"01111101", "01111110", "01111111", "01111111", "01111111", "01111110", "01111101", "01111100", "01111010", "01111000", "01110101", "01110011", "01110000", "01101101", "01101011", "01101000", "01100101", "01100010", "01011111", "01011100", 
"01011010", "01011100", "01011111", "01100001", "01100011", "01100100", "01100110", "01101000", "01101001", "01101010", "01101011", "01101101", "01101110", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", 
"01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110110", "01110101", "01110101", 
"01110100", "01110100", "01110011", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101110", "01101101", "01101011", "01101010", "01101001", "01101000", "01100110", "01100100", "01100011", "01100001", 
"01011111", "01011100", "01011010", "01011100", "01011111", "01100010", "01100101", "01101000", "01101011", "01101101", "01110000", "01110011", "01110101", "01111000", "01111010", "01111100", "01111101", "01111110", "01111111", "01111111", 
"01111111", "01111110", "01111101", "01111011", "01111001", "01110111", "01110100", "01110010", "01101111", "01101100", "01101001", "01100110", "01100011", "01100000", "01011101", "01011010", "01011100", "01011111", "01100001", "01100011", 
"01100101", "01100111", "01101000", "01101010", "01101011", "01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110101", "01110110", 
"01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110101", "01110100", 
"01110100", "01110011", "01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101011", "01101010", "01101000", "01100111", "01100101", "01100011", "01100001", "01011111", "01011100", "01011010", 
"01011101", "01100000", "01100011", "01100110", "01101001", "01101100", "01101111", "01110010", "01110100", "01110111", "01111001", "01111011", "01111101", "01111110", "01111111", "01111111", "01111111", "01111110", "01111101", "01111011", 
"01111000", "01110110", "01110011", "01110000", "01101101", "01101010", "01100110", "01100011", "01100000", "01011101", "01011010", "01011101", "01011111", "01100010", "01100100", "01100110", "01100111", "01101001", "01101010", "01101100", 
"01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", 
"01111010", "01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", 
"01110010", "01110010", "01110001", "01110000", "01101111", "01101110", "01101101", "01101100", "01101010", "01101001", "01100111", "01100110", "01100100", "01100010", "01011111", "01011101", "01011010", "01011101", "01100000", "01100011", 
"01100110", "01101010", "01101101", "01110000", "01110011", "01110110", "01111000", "01111011", "01111101", "01111110", "01111111", "01111111", "01111111", "01111110", "01111100", "01111010", "01111000", "01110101", "01110010", "01101110", 
"01101011", "01100111", "01100100", "01100000", "01011101", "01011010", "01011101", "01100000", "01100010", "01100100", "01100110", "01101000", "01101010", "01101011", "01101100", "01101110", "01101111", "01110000", "01110001", "01110010", 
"01110010", "01110011", "01110100", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111001", "01111010", "01111010", 
"01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111001", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110100", "01110011", "01110010", "01110010", 
"01110001", "01110000", "01101111", "01101110", "01101100", "01101011", "01101010", "01101000", "01100110", "01100100", "01100010", "01100000", "01011101", "01011010", "01011101", "01100000", "01100100", "01100111", "01101011", "01101110", 
"01110010", "01110101", "01111000", "01111010", "01111100", "01111110", "01111111", "01111111", "01111111", "01111110", "01111100", "01111001", "01110111", "01110011", "01110000", "01101100", "01101000", "01100101", "01100001", "01011101", 
"01011010", "01011101", "01100000", "01100011", "01100101", "01100111", "01101001", "01101010", "01101100", "01101101", "01101111", "01110000", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", 
"01110110", "01110111", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", 
"01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", 
"01111010", "01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01110000", 
"01101111", "01101101", "01101100", "01101010", "01101001", "01100111", "01100101", "01100011", "01100000", "01011101", "01011010", "01011101", "01100001", "01100101", "01101000", "01101100", "01110000", "01110011", "01110111", "01111001", 
"01111100", "01111110", "01111111", "01111111", "01111111", "01111101", "01111011", "01111000", "01110101", "01110010", "01101110", "01101010", "01100110", "01100010", "01011110", "01011010", "01011101", "01100000", "01100011", "01100110", 
"01101000", "01101010", "01101011", "01101101", "01101110", "01101111", "01110001", "01110010", "01110010", "01110011", "01110100", "01110101", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", 
"01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", 
"01111001", "01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110101", "01110100", "01110011", "01110010", "01110010", "01110001", "01101111", "01101110", "01101101", 
"01101011", "01101010", "01101000", "01100110", "01100011", "01100000", "01011101", "01011010", "01011110", "01100010", "01100110", "01101010", "01101110", "01110010", "01110101", "01111000", "01111011", "01111101", "01111111", "01111111", 
"01111110", "01111101", "01111011", "01110111", "01110100", "01101111", "01101011", "01100111", "01100010", "01011110", "01011010", "01011110", "01100001", "01100100", "01100110", "01101001", "01101011", "01101100", "01101110", "01101111", 
"01110001", "01110010", "01110011", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", 
"01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110011", "01110010", "01110001", "01101111", "01101110", "01101100", "01101011", "01101001", 
"01100110", "01100100", "01100001", "01011110", "01011010", "01011110", "01100010", "01100111", "01101011", "01101111", "01110100", "01110111", "01111011", "01111101", "01111110", "01111111", "01111110", "01111101", "01111010", "01110110", 
"01110010", "01101101", "01101000", "01100011", "01011110", "01011010", "01011110", "01100010", "01100101", "01100111", "01101010", "01101100", "01101101", "01101111", "01110000", "01110010", "01110011", "01110100", "01110100", "01110101", 
"01110110", "01110111", "01110111", "01111000", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", 
"01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111010", "01111001", 
"01111001", "01111000", "01111000", "01111000", "01110111", "01110111", "01110110", "01110101", "01110100", "01110100", "01110011", "01110010", "01110000", "01101111", "01101101", "01101100", "01101010", "01100111", "01100101", "01100010", 
"01011110", "01011010", "01011110", "01100011", "01101000", "01101101", "01110010", "01110110", "01111010", "01111101", "01111110", "01111111", "01111110", "01111100", "01111000", "01110100", "01101111", "01101010", "01100100", "01011111", 
"01011010", "01011110", "01100010", "01100110", "01101000", "01101011", "01101101", "01101111", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", 
"01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", 
"01111000", "01111000", "01110111", "01110111", "01110110", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101111", "01101101", "01101011", "01101000", "01100110", "01100010", "01011110", "01011010", "01011111", 
"01100100", "01101010", "01101111", "01110100", "01111000", "01111100", "01111110", "01111111", "01111110", "01111011", "01110111", "01110010", "01101100", "01100110", "01100000", "01011010", "01011111", "01100011", "01100111", "01101010", 
"01101100", "01101110", "01110000", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111010", "01111011", "01111011", "01111011", 
"01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111010", "01111001", "01111001", "01111000", 
"01111000", "01110111", "01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101110", "01101100", "01101010", "01100111", "01100011", "01011111", "01011010", "01100000", "01100110", "01101100", "01110010", 
"01110111", "01111011", "01111110", "01111111", "01111110", "01111010", "01110101", "01101110", "01100111", "01100000", "01011010", "01100000", "01100100", "01101000", "01101011", "01101110", "01110000", "01110010", "01110011", "01110100", 
"01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111001", "01111010", "01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111001", "01111000", "01111000", 
"01110111", "01110110", "01110101", "01110100", "01110011", "01110010", "01110000", "01101110", "01101011", "01101000", "01100100", "01100000", "01011010", "01100000", "01100111", "01101110", "01110101", "01111010", "01111110", "01111111", 
"01111101", "01111000", "01110010", "01101010", "01100010", "01011010", "01100000", "01100110", "01101010", "01101101", "01101111", "01110010", "01110011", "01110101", "01110110", "01110111", "01111000", "01111000", "01111001", "01111010", 
"01111010", "01111011", "01111011", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", 
"01110110", "01110101", "01110011", "01110010", "01101111", "01101101", "01101010", "01100110", "01100000", "01011010", "01100010", "01101010", "01110010", "01111000", "01111101", "01111111", "01111101", "01110110", "01101101", "01100011", 
"01011010", "01100010", "01100111", "01101100", "01101111", "01110010", "01110100", "01110101", "01110111", "01111000", "01111000", "01111001", "01111010", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111100", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", 
"01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111010", "01111001", "01111000", "01111000", "01110111", "01110101", 
"01110100", "01110010", "01101111", "01101100", "01100111", "01100010", "01011010", "01100011", "01101101", "01110110", "01111101", "01111111", "01111011", "01110010", "01100110", "01011010", "01100011", "01101010", "01101110", "01110010", 
"01110100", "01110110", "01110111", "01111000", "01111001", "01111010", "01111011", "01111011", "01111100", "01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111100", "01111011", "01111011", "01111010", "01111001", "01111000", "01110111", "01110110", "01110100", "01110010", 
"01101110", "01101010", "01100011", "01011010", "01100110", "01110010", "01111011", "01111111", "01111000", "01101010", "01011010", "01100110", "01101101", "01110010", "01110101", "01110111", "01111000", "01111010", "01111011", "01111011", 
"01111100", "01111100", "01111101", "01111101", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111101", "01111101", "01111100", "01111100", "01111011", "01111011", "01111010", "01111000", "01110111", "01110101", "01110010", "01101101", "01100110", 
"01011010", "01101010", "01111000", "01111111", "01110010", "01011010", "01101010", "01110010", "01110110", "01111000", "01111010", "01111011", "01111100", "01111101", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", 
"01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111101", "01111100", "01111011", "01111010", "01111000", "01110110", "01110010", "01101010", "01011010", "01110010", "01111111", 
"01011010", "01110010", "01111000", "01111011", "01111101", "01111101", "01111110", "01111110", "01111110", "01111110", "01111110", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", "01111111", 
"01111111", "01111111", "01111111", "01111111", "01111110", "01111110", "01111110", "01111110", "01111110", "01111101", "01111101", "01111011", "01111000", "01110010", "01011010" );
constant mem_im:Tmem:=  (
"00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "10100110", "00111001", "00101000", "00011111", 
"00011001", "00010101", "00010010", "00010000", "00001110", "00001101", "00001011", "00001011", "00001010", "00001001", "00001000", "00001000", "00000111", "00000111", "00000111", "00000110", "00000110", "00000110", "00000110", "00000101", 
"00000101", "00000101", "00000101", "00000101", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", 
"00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", 
"00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", 
"00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", 
"00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", 
"00000001", "00000001", "00000001", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", 
"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", 
"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", 
"11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", 
"11111110", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111100", "11111100", "11111100", "11111100", "11111100", 
"11111100", "11111100", "11111100", "11111011", "11111011", "11111011", "11111011", "11111011", "11111010", "11111010", "11111010", "11111010", "11111001", "11111001", "11111001", "11111000", "11111000", "11110111", "11110110", "11110101", 
"11110101", "11110011", "11110010", "11110000", "11101110", "11101011", "11100111", "11100001", "11011000", "11000111", "10100110", "00000000", "11000111", "10100110", "01000110", "00111001", "00101111", "00101000", "00100011", "00011111", 
"00011100", "00011001", "00010111", "00010101", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001101", "00001100", "00001011", "00001011", "00001011", "00001010", "00001010", "00001001", "00001001", 
"00001001", "00001000", "00001000", "00001000", "00001000", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000101", "00000101", 
"00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", 
"00000100", "00000100", "00000100", "00000100", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", 
"00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", 
"00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "11111110", 
"11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", 
"11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", 
"11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111100", "11111100", "11111100", "11111100", "11111100", 
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", 
"11111011", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111000", "11111000", "11111000", "11111000", "11110111", "11110111", 
"11110111", "11110110", "11110110", "11110101", "11110101", "11110101", "11110100", "11110011", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101011", "11101001", "11100111", "11100100", "11100001", 
"11011101", "11011000", "11010001", "11000111", "10111010", "10100110", "00111001", "00000000", "11011000", "10111010", "10100110", "01001100", "01000001", "00111001", "00110010", "00101101", "00101000", "00100100", "00100001", "00011111", 
"00011101", "00011011", "00011001", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00010000", "00001111", "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001100", 
"00001011", "00001011", "00001011", "00001011", "00001010", "00001010", "00001010", "00001001", "00001001", "00001001", "00001001", "00001001", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00000111", "00000111", 
"00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000101", "00000101", "00000101", 
"00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", 
"00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000011", "00000011", "00000011", "00000011", 
"00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "11111101", "11111101", "11111101", "11111101", "11111101", 
"11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111100", "11111100", "11111100", "11111100", "11111100", 
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111011", 
"11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", 
"11111010", "11111010", "11111010", "11111010", "11111010", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11110111", 
"11110111", "11110111", "11110111", "11110111", "11110110", "11110110", "11110110", "11110101", "11110101", "11110101", "11110101", "11110100", "11110100", "11110011", "11110011", "11110010", "11110010", "11110001", "11110001", "11110000", 
"11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11100111", "11100101", "11100011", "11100001", "11011111", "11011100", "11011000", "11010011", "11001110", "11000111", "10111111", "10110100", 
"10100110", "01000110", "00101000", "00000000", "11100001", "11000111", "10110100", "10100110", "01001111", "01000110", "00111111", "00111001", "00110100", "00101111", "00101011", "00101000", "00100101", "00100011", "00100001", "00011111", 
"00011101", "00011100", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010011", "00010010", "00010001", "00010001", "00010000", "00010000", "00001111", "00001111", "00001110", "00001110", 
"00001110", "00001101", "00001101", "00001101", "00001100", "00001100", "00001100", "00001011", "00001011", "00001011", "00001011", "00001011", "00001010", "00001010", "00001010", "00001010", "00001010", "00001001", "00001001", "00001001", 
"00001001", "00001001", "00001001", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", 
"00000111", "00000111", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000101", "00000101", "00000101", "00000101", 
"00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000100", "00000100", "00000100", "00000100", 
"00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", 
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", 
"11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", 
"11111010", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", 
"11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110110", "11110110", "11110110", "11110110", "11110110", "11110101", "11110101", "11110101", "11110101", "11110101", "11110100", "11110100", "11110100", "11110011", 
"11110011", "11110011", "11110010", "11110010", "11110010", "11110001", "11110001", "11110000", "11110000", "11101111", "11101111", "11101110", "11101101", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", 
"11100110", "11100100", "11100011", "11100001", "11011111", "11011101", "11011011", "11011000", "11010101", "11010001", "11001100", "11000111", "11000001", "10111010", "10110001", "10100110", "01001100", "00111001", "00011111", "00000000", 
"11100111", "11010001", "10111111", "10110001", "10100110", "01010001", "01001010", "01000011", "00111110", "00111001", "00110101", "00110001", "00101110", "00101011", "00101000", "00100110", "00100100", "00100010", "00100000", "00011111", 
"00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010110", "00010101", "00010100", "00010100", "00010011", "00010010", "00010010", "00010001", "00010001", "00010001", "00010000", "00010000", 
"00001111", "00001111", "00001111", "00001110", "00001110", "00001110", "00001101", "00001101", "00001101", "00001101", "00001100", "00001100", "00001100", "00001100", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", 
"00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", 
"00001000", "00001000", "00001000", "00001000", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000110", "00000110", "00000110", 
"00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000101", "00000101", "00000101", "00000101", "00000101", 
"00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", 
"11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111001", "11111001", 
"11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", 
"11111000", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110101", "11110101", "11110101", "11110101", "11110101", 
"11110101", "11110100", "11110100", "11110100", "11110100", "11110011", "11110011", "11110011", "11110011", "11110010", "11110010", "11110010", "11110001", "11110001", "11110001", "11110000", "11110000", "11101111", "11101111", "11101111", 
"11101110", "11101110", "11101101", "11101100", "11101100", "11101011", "11101010", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100001", "11100000", "11011110", "11011100", "11011010", 
"11011000", "11010101", "11010010", "11001111", "11001011", "11000111", "11000010", "10111101", "10110110", "10101111", "10100110", "01001111", "01000001", "00101111", "00011001", "00000000", "11101011", "11011000", "11000111", "10111010", 
"10101111", "10100110", "01010011", "01001100", "01000110", "01000001", "00111101", "00111001", "00110101", "00110010", "00101111", "00101101", "00101010", "00101000", "00100110", "00100100", "00100011", "00100001", "00100000", "00011111", 
"00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010111", "00010110", "00010101", "00010101", "00010100", "00010100", "00010011", "00010011", "00010010", "00010010", "00010010", "00010001", 
"00010001", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001111", "00001110", "00001110", "00001110", "00001110", "00001101", "00001101", "00001101", "00001101", "00001100", "00001100", "00001100", "00001100", 
"00001100", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001001", "00001001", "00001001", "00001001", "00001001", 
"00001001", "00001001", "00001001", "00001001", "00001001", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00000111", "00000111", "00000111", 
"00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", 
"00000110", "00000110", "00000110", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", 
"11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", 
"11111000", "11111000", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110101", 
"11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110100", "11110100", "11110100", "11110100", "11110100", "11110011", "11110011", "11110011", "11110011", "11110010", "11110010", "11110010", "11110010", "11110001", 
"11110001", "11110001", "11110001", "11110000", "11110000", "11110000", "11101111", "11101111", "11101110", "11101110", "11101110", "11101101", "11101101", "11101100", "11101100", "11101011", "11101011", "11101010", "11101001", "11101001", 
"11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011101", "11011100", "11011010", "11011000", "11010110", "11010011", "11010001", "11001110", "11001011", "11000111", 
"11000011", "10111111", "10111010", "10110100", "10101101", "10100110", "01010001", "01000110", "00111001", "00101000", "00010101", "00000000", "11101110", "11011101", "11001110", "11000001", "10110110", "10101101", "10100110", "01010100", 
"01001110", "01001001", "01000100", "01000000", "00111100", "00111001", "00110110", "00110011", "00110000", "00101110", "00101100", "00101010", "00101000", "00100111", "00100101", "00100100", "00100010", "00100001", "00100000", "00011111", 
"00011110", "00011101", "00011100", "00011011", "00011010", "00011010", "00011001", "00011000", "00011000", "00010111", "00010110", "00010110", "00010101", "00010101", "00010100", "00010100", "00010100", "00010011", "00010011", "00010010", 
"00010010", "00010010", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001111", "00001110", "00001110", "00001110", "00001110", "00001110", "00001101", "00001101", "00001101", 
"00001101", "00001101", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001010", "00001010", "00001010", "00001010", 
"00001010", "00001010", "00001010", "00001010", "00001010", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001000", "00001000", "00001000", "00001000", 
"00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "11111001", 
"11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", 
"11111000", "11111000", "11111000", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", 
"11110110", "11110110", "11110110", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110011", "11110011", "11110011", 
"11110011", "11110011", "11110010", "11110010", "11110010", "11110010", "11110010", "11110001", "11110001", "11110001", "11110001", "11110000", "11110000", "11110000", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", 
"11101101", "11101101", "11101100", "11101100", "11101100", "11101011", "11101011", "11101010", "11101010", "11101001", "11101000", "11101000", "11100111", "11100110", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", 
"11100000", "11011111", "11011110", "11011100", "11011011", "11011001", "11011000", "11010110", "11010100", "11010010", "11010000", "11001101", "11001010", "11000111", "11000100", "11000000", "10111100", "10110111", "10110010", "10101100", 
"10100110", "01010011", "01001010", "00111111", "00110010", "00100011", "00010010", "00000000", "11110000", "11100001", "11010011", "11000111", "10111101", "10110100", "10101100", "10100110", "01010100", "01001111", "01001011", "01000110", 
"01000011", "00111111", "00111100", "00111001", "00110110", "00110100", "00110001", "00101111", "00101101", "00101011", "00101010", "00101000", "00100111", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", 
"00011110", "00011101", "00011100", "00011100", "00011011", "00011010", "00011010", "00011001", "00011000", "00011000", "00010111", "00010111", "00010110", "00010110", "00010101", "00010101", "00010100", "00010100", "00010100", "00010011", 
"00010011", "00010011", "00010010", "00010010", "00010010", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001111", "00001110", "00001110", "00001110", 
"00001110", "00001110", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001011", "00001011", "00001011", "00001011", "00001011", 
"00001011", "00001011", "00001011", "00001011", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", 
"00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "11111000", "11111000", "11111000", "11111000", "11111000", 
"11111000", "11111000", "11111000", "11111000", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110110", "11110110", "11110110", 
"11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110100", "11110100", "11110100", "11110100", 
"11110100", "11110100", "11110100", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110010", "11110010", "11110010", "11110010", "11110010", "11110001", "11110001", "11110001", "11110001", "11110000", "11110000", 
"11110000", "11110000", "11101111", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", "11101101", "11101101", "11101101", "11101100", "11101100", "11101100", "11101011", "11101011", "11101010", "11101010", "11101001", 
"11101001", "11101000", "11101000", "11100111", "11100110", "11100110", "11100101", "11100100", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011001", "11011000", 
"11010110", "11010101", "11010011", "11010001", "11001111", "11001100", "11001010", "11000111", "11000100", "11000001", "10111101", "10111010", "10110101", "10110001", "10101100", "10100110", "01010100", "01001100", "01000011", "00111001", 
"00101101", "00011111", "00010000", "00000000", "11110010", "11100100", "11011000", "11001100", "11000010", "10111010", "10110010", "10101100", "10100110", "01010101", "01010000", "01001100", "01001000", "01000101", "01000001", "00111110", 
"00111011", "00111001", "00110110", "00110100", "00110010", "00110000", "00101110", "00101101", "00101011", "00101010", "00101000", "00100111", "00100110", "00100100", "00100011", "00100010", "00100001", "00100000", "00100000", "00011111", 
"00011110", "00011101", "00011101", "00011100", "00011011", "00011011", "00011010", "00011001", "00011001", "00011000", "00011000", "00010111", "00010111", "00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010100", 
"00010100", "00010011", "00010011", "00010011", "00010011", "00010010", "00010010", "00010010", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", 
"00001111", "00001111", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", 
"00001100", "00001100", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", 
"00001010", "00001010", "00001010", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", 
"11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", 
"11110101", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110010", "11110010", "11110010", "11110010", "11110010", 
"11110010", "11110001", "11110001", "11110001", "11110001", "11110001", "11110000", "11110000", "11110000", "11110000", "11110000", "11101111", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", "11101101", "11101101", 
"11101101", "11101101", "11101100", "11101100", "11101011", "11101011", "11101011", "11101010", "11101010", "11101010", "11101001", "11101001", "11101000", "11101000", "11100111", "11100111", "11100110", "11100101", "11100101", "11100100", 
"11100011", "11100011", "11100010", "11100001", "11100000", "11100000", "11011111", "11011110", "11011101", "11011100", "11011010", "11011001", "11011000", "11010110", "11010101", "11010011", "11010010", "11010000", "11001110", "11001100", 
"11001010", "11000111", "11000101", "11000010", "10111111", "10111011", "10111000", "10110100", "10110000", "10101011", "10100110", "01010100", "01001110", "01000110", "00111110", "00110100", "00101000", "00011100", "00001110", "00000000", 
"11110011", "11100111", "11011100", "11010001", "11000111", "10111111", "10110111", "10110001", "10101011", "10100110", "01010101", "01010001", "01001101", "01001010", "01000110", "01000011", "01000000", "00111110", "00111011", "00111001", 
"00110111", "00110101", "00110011", "00110001", "00101111", "00101110", "00101100", "00101011", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00100000", "00011111", 
"00011110", "00011101", "00011101", "00011100", "00011100", "00011011", "00011010", "00011010", "00011001", "00011001", "00011000", "00011000", "00011000", "00010111", "00010111", "00010110", "00010110", "00010110", "00010101", "00010101", 
"00010101", "00010100", "00010100", "00010100", "00010011", "00010011", "00010011", "00010010", "00010010", "00010010", "00010010", "00010001", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", 
"00010000", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", 
"00001101", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", 
"00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110101", "11110101", "11110101", "11110101", "11110101", 
"11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", 
"11110011", "11110011", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110000", "11110000", "11110000", "11110000", "11110000", "11101111", 
"11101111", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", "11101110", "11101101", "11101101", "11101101", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101010", "11101010", "11101010", 
"11101001", "11101001", "11101000", "11101000", "11101000", "11100111", "11100111", "11100110", "11100110", "11100101", "11100100", "11100100", "11100011", "11100011", "11100010", "11100001", "11100000", "11100000", "11011111", "11011110", 
"11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010101", "11010100", "11010010", "11010001", "11001111", "11001101", "11001011", "11001001", "11000111", "11000101", "11000010", "11000000", "10111101", 
"10111010", "10110110", "10110011", "10101111", "10101011", "10100110", "01010101", "01001111", "01001001", "01000001", "00111001", "00101111", "00100100", "00011001", "00001101", "00000000", "11110101", "11101001", "11011111", "11010101", 
"11001011", "11000011", "10111100", "10110101", "10110000", "10101011", "10100110", "01010110", "01010010", "01001110", "01001011", "01001000", "01000101", "01000010", "01000000", "00111101", "00111011", "00111001", "00110111", "00110101", 
"00110011", "00110001", "00110000", "00101110", "00101101", "00101100", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100010", "00100001", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011101", "00011100", "00011100", "00011011", "00011011", "00011010", "00011010", "00011001", "00011001", "00011000", "00011000", "00011000", "00010111", "00010111", "00010111", "00010110", "00010110", "00010110", 
"00010101", "00010101", "00010101", "00010100", "00010100", "00010100", "00010011", "00010011", "00010011", "00010011", "00010010", "00010010", "00010010", "00010010", "00010010", "00010001", "00010001", "00010001", "00010001", "00010000", 
"00010000", "00010000", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001101", "00001101", 
"00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001011", "00001011", "00001011", "00001011", 
"00001011", "00001011", "00001011", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", 
"11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110001", "11110001", "11110001", "11110001", 
"11110001", "11110001", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11101111", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", "11101110", "11101110", "11101101", "11101101", "11101101", 
"11101101", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", "11100111", "11100111", "11100110", "11100110", 
"11100101", "11100101", "11100100", "11100100", "11100011", "11100010", "11100010", "11100001", "11100001", "11100000", "11011111", "11011110", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", 
"11010110", "11010100", "11010011", "11010010", "11010000", "11001111", "11001101", "11001011", "11001001", "11000111", "11000101", "11000011", "11000000", "10111110", "10111011", "10111000", "10110101", "10110010", "10101110", "10101010", 
"10100110", "01010101", "01010000", "01001011", "01000100", "00111101", "00110101", "00101011", "00100001", "00010111", "00001011", "00000000", "11110101", "11101011", "11100001", "11011000", "11001111", "11000111", "11000000", "10111010", 
"10110100", "10101111", "10101010", "10100110", "01010110", "01010011", "01001111", "01001100", "01001001", "01000110", "01000100", "01000001", "00111111", "00111101", "00111011", "00111001", "00110111", "00110101", "00110100", "00110010", 
"00110001", "00101111", "00101110", "00101101", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100100", "00100011", "00100010", "00100001", "00100001", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011101", "00011101", "00011100", "00011100", "00011011", "00011011", "00011010", "00011010", "00011001", "00011001", "00011001", "00011000", "00011000", "00010111", "00010111", "00010111", "00010110", "00010110", 
"00010110", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", "00010100", "00010100", "00010011", "00010011", "00010011", "00010011", "00010010", "00010010", "00010010", "00010010", "00010010", "00010001", "00010001", 
"00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001110", "00001110", "00001110", "00001110", 
"00001110", "00001110", "00001110", "00001110", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "11110100", 
"11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110010", "11110010", "11110010", "11110010", "11110010", 
"11110010", "11110010", "11110010", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11101111", "11101111", "11101111", "11101111", 
"11101111", "11101110", "11101110", "11101110", "11101110", "11101110", "11101101", "11101101", "11101101", "11101101", "11101100", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101010", "11101010", 
"11101010", "11101001", "11101001", "11101001", "11101000", "11101000", "11100111", "11100111", "11100111", "11100110", "11100110", "11100101", "11100101", "11100100", "11100100", "11100011", "11100011", "11100010", "11100010", "11100001", 
"11100001", "11100000", "11011111", "11011111", "11011110", "11011101", "11011100", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010011", "11010010", "11010001", "11001111", "11001110", 
"11001100", "11001011", "11001001", "11000111", "11000101", "11000011", "11000001", "10111111", "10111100", "10111010", "10110111", "10110100", "10110001", "10101101", "10101010", "10100110", "01010110", "01010001", "01001100", "01000110", 
"01000000", "00111001", "00110001", "00101000", "00011111", "00010101", "00001011", "00000000", "11110110", "11101101", "11100011", "11011011", "11010010", "11001011", "11000100", "10111101", "10111000", "10110011", "10101110", "10101010", 
"10100110", "01010110", "01010011", "01010000", "01001101", "01001010", "01001000", "01000101", "01000011", "01000001", "00111110", "00111100", "00111011", "00111001", "00110111", "00110101", "00110100", "00110010", "00110001", "00110000", 
"00101111", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100110", "00100101", "00100100", "00100011", "00100011", "00100010", "00100001", "00100001", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011101", "00011101", "00011100", "00011100", "00011011", "00011011", "00011010", "00011010", "00011010", "00011001", "00011001", "00011001", "00011000", "00011000", "00011000", "00010111", "00010111", "00010111", 
"00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", "00010100", "00010100", "00010011", "00010011", "00010011", "00010011", "00010011", "00010010", "00010010", "00010010", "00010010", 
"00010010", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", 
"00001111", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "11110011", "11110011", "11110011", "11110011", "11110011", 
"11110011", "11110011", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110000", "11110000", 
"11110000", "11110000", "11110000", "11110000", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", "11101110", "11101110", "11101101", "11101101", "11101101", "11101101", "11101101", 
"11101100", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", 
"11100110", "11100110", "11100110", "11100101", "11100101", "11100100", "11100100", "11100011", "11100011", "11100010", "11100010", "11100001", "11100001", "11100000", "11011111", "11011111", "11011110", "11011101", "11011101", "11011100", 
"11011011", "11011010", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010001", "11010000", "11001111", "11001110", "11001100", "11001011", "11001001", "11000111", "11000101", "11000100", 
"11000010", "10111111", "10111101", "10111011", "10111000", "10110110", "10110011", "10110000", "10101101", "10101010", "10100110", "01010110", "01010010", "01001101", "01001000", "01000011", "00111100", "00110101", "00101110", "00100101", 
"00011101", "00010011", "00001010", "00000000", "11110111", "11101110", "11100101", "11011101", "11010101", "11001110", "11000111", "11000001", "10111011", "10110110", "10110010", "10101101", "10101010", "10100110", "01010111", "01010100", 
"01010001", "01001110", "01001011", "01001001", "01000110", "01000100", "01000010", "01000000", "00111110", "00111100", "00111010", "00111001", "00110111", "00110110", "00110100", "00110011", "00110010", "00110000", "00101111", "00101110", 
"00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100111", "00100110", "00100101", "00100100", "00100100", "00100011", "00100010", "00100010", "00100001", "00100000", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011101", "00011101", "00011100", "00011100", "00011100", "00011011", "00011011", "00011010", "00011010", "00011010", "00011001", "00011001", "00011001", "00011000", "00011000", "00011000", "00010111", "00010111", 
"00010111", "00010110", "00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", "00010100", "00010100", "00010100", "00010011", "00010011", "00010011", "00010011", "00010011", "00010010", 
"00010010", "00010010", "00010010", "00010010", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00001111", "00001111", "00001111", 
"00001111", "00001111", "00001111", "00001111", "00001111", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110001", "11110001", 
"11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11101110", 
"11101110", "11101110", "11101110", "11101110", "11101101", "11101101", "11101101", "11101101", "11101101", "11101100", "11101100", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101010", "11101010", 
"11101010", "11101010", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", "11100110", "11100110", "11100110", "11100101", "11100101", "11100100", "11100100", "11100100", "11100011", 
"11100011", "11100010", "11100010", "11100001", "11100001", "11100000", "11100000", "11011111", "11011110", "11011110", "11011101", "11011100", "11011100", "11011011", "11011010", "11011001", "11011001", "11011000", "11010111", "11010110", 
"11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001110", "11001101", "11001100", "11001010", "11001001", "11000111", "11000110", "11000100", "11000010", "11000000", "10111110", "10111100", "10111010", "10110111", 
"10110101", "10110010", "10101111", "10101100", "10101001", "10100110", "01010110", "01010011", "01001110", "01001010", "01000101", "00111111", "00111001", "00110010", "00101011", "00100011", "00011011", "00010010", "00001001", "00000000", 
"11111000", "11101111", "11100111", "11011111", "11011000", "11010001", "11001010", "11000100", "10111111", "10111010", "10110101", "10110001", "10101101", "10101001", "10100110", "01010111", "01010100", "01010001", "01001111", "01001100", 
"01001010", "01001000", "01000101", "01000011", "01000001", "00111111", "00111110", "00111100", "00111010", "00111001", "00110111", "00110110", "00110101", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", 
"00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100111", "00100110", "00100101", "00100100", "00100100", "00100011", "00100011", "00100010", "00100001", "00100001", "00100000", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011101", "00011101", "00011101", "00011100", "00011100", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011001", "00011001", "00011001", "00011000", "00011000", "00011000", "00010111", 
"00010111", "00010111", "00010111", "00010110", "00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", "00010100", "00010100", "00010100", "00010011", "00010011", "00010011", "00010011", 
"00010011", "00010010", "00010010", "00010010", "00010010", "00010010", "00010010", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", 
"00010000", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", 
"11110000", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", "11101110", "11101110", "11101110", "11101101", "11101101", "11101101", "11101101", "11101101", "11101100", 
"11101100", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101010", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", "11100111", 
"11100111", "11100111", "11100110", "11100110", "11100110", "11100101", "11100101", "11100101", "11100100", "11100100", "11100011", "11100011", "11100011", "11100010", "11100010", "11100001", "11100001", "11100000", "11100000", "11011111", 
"11011111", "11011110", "11011101", "11011101", "11011100", "11011100", "11011011", "11011010", "11011001", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", 
"11001110", "11001101", "11001011", "11001010", "11001001", "11000111", "11000110", "11000100", "11000010", "11000001", "10111111", "10111101", "10111011", "10111000", "10110110", "10110100", "10110001", "10101111", "10101100", "10101001", 
"10100110", "01010111", "01010011", "01001111", "01001011", "01000110", "01000001", "00111100", "00110110", "00101111", "00101000", "00100001", "00011001", "00010001", "00001000", "00000000", "11111000", "11110000", "11101001", "11100001", 
"11011010", "11010011", "11001101", "11000111", "11000010", "10111101", "10111000", "10110100", "10110000", "10101100", "10101001", "10100110", "01010111", "01010100", "01010010", "01001111", "01001101", "01001011", "01001001", "01000110", 
"01000100", "01000011", "01000001", "00111111", "00111101", "00111100", "00111010", "00111001", "00110111", "00110110", "00110101", "00110100", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", 
"00101011", "00101010", "00101001", "00101000", "00100111", "00100111", "00100110", "00100101", "00100101", "00100100", "00100011", "00100011", "00100010", "00100010", "00100001", "00100001", "00100000", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011011", "00011011", "00011010", "00011010", "00011010", "00011010", "00011001", "00011001", "00011001", "00011000", "00011000", "00011000", 
"00010111", "00010111", "00010111", "00010111", "00010110", "00010110", "00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", "00010100", "00010100", "00010100", "00010011", "00010011", 
"00010011", "00010011", "00010011", "00010011", "00010010", "00010010", "00010010", "00010010", "00010010", "00010010", "00010010", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010000", "00010000", 
"00010000", "00010000", "00010000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", "11101110", 
"11101110", "11101110", "11101110", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101100", "11101100", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101010", "11101010", 
"11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", "11100110", "11100110", "11100110", "11100110", "11100101", "11100101", "11100100", 
"11100100", "11100100", "11100011", "11100011", "11100011", "11100010", "11100010", "11100001", "11100001", "11100000", "11100000", "11011111", "11011111", "11011110", "11011110", "11011101", "11011101", "11011100", "11011011", "11011011", 
"11011010", "11011001", "11011001", "11011000", "11010111", "11010110", "11010101", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001100", "11001011", "11001010", "11001001", "11000111", 
"11000110", "11000100", "11000011", "11000001", "10111111", "10111101", "10111100", "10111010", "10110111", "10110101", "10110011", "10110001", "10101110", "10101100", "10101001", "10100110", "01010111", "01010100", "01010000", "01001100", 
"01001000", "01000011", "00111110", "00111001", "00110011", "00101101", "00100110", "00011111", "00010111", "00010000", "00001000", "00000000", "11111001", "11110001", "11101010", "11100011", "11011100", "11010110", "11010000", "11001010", 
"11000101", "11000000", "10111011", "10110111", "10110011", "10101111", "10101100", "10101001", "10100110", "01010111", "01010101", "01010010", "01010000", "01001110", "01001011", "01001001", "01000111", "01000110", "01000100", "01000010", 
"01000000", "00111111", "00111101", "00111100", "00111010", "00111001", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", 
"00101010", "00101001", "00101000", "00100111", "00100111", "00100110", "00100110", "00100101", "00100100", "00100100", "00100011", "00100011", "00100010", "00100010", "00100001", "00100001", "00100000", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011110", "00011101", "00011101", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011001", "00011001", "00011001", "00011001", "00011000", "00011000", 
"00011000", "00011000", "00010111", "00010111", "00010111", "00010111", "00010110", "00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", "00010100", "00010100", "00010100", 
"00010100", "00010011", "00010011", "00010011", "00010011", "00010011", "00010011", "00010010", "00010010", "00010010", "00010010", "00010010", "00010010", "00010010", "00010001", "00010001", "00010001", "00010001", "00010001", "11101111", 
"11101111", "11101111", "11101111", "11101111", "11101111", "11101110", "11101110", "11101110", "11101110", "11101110", "11101110", "11101110", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101100", "11101100", 
"11101100", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101011", "11101010", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", 
"11101000", "11100111", "11100111", "11100111", "11100111", "11100110", "11100110", "11100110", "11100101", "11100101", "11100101", "11100100", "11100100", "11100100", "11100011", "11100011", "11100010", "11100010", "11100010", "11100001", 
"11100001", "11100000", "11100000", "11011111", "11011111", "11011110", "11011110", "11011101", "11011101", "11011100", "11011100", "11011011", "11011010", "11011010", "11011001", "11011001", "11011000", "11010111", "11010110", "11010110", 
"11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11000111", "11000110", "11000100", "11000011", "11000001", "11000000", "10111110", 
"10111100", "10111010", "10111001", "10110111", "10110101", "10110010", "10110000", "10101110", "10101011", "10101001", "10100110", "01010111", "01010100", "01010001", "01001101", "01001001", "01000101", "01000000", "00111011", "00110110", 
"00110000", "00101010", "00100100", "00011101", "00010110", "00001111", "00000111", "00000000", "11111001", "11110010", "11101011", "11100100", "11011110", "11011000", "11010010", "11001100", "11000111", "11000010", "10111110", "10111010", 
"10110110", "10110010", "10101111", "10101100", "10101001", "10100110", "01010111", "01010101", "01010011", "01010000", "01001110", "01001100", "01001010", "01001000", "01000110", "01000101", "01000011", "01000001", "01000000", "00111110", 
"00111101", "00111011", "00111010", "00111001", "00111000", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101101", "00101100", "00101011", "00101010", "00101010", 
"00101001", "00101000", "00101000", "00100111", "00100110", "00100110", "00100101", "00100100", "00100100", "00100011", "00100011", "00100010", "00100010", "00100001", "00100001", "00100000", "00100000", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011001", "00011001", "00011001", "00011001", "00011000", 
"00011000", "00011000", "00011000", "00010111", "00010111", "00010111", "00010111", "00010110", "00010110", "00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010101", "00010101", "00010101", "00010100", "00010100", 
"00010100", "00010100", "00010100", "00010011", "00010011", "00010011", "00010011", "00010011", "00010011", "00010011", "00010010", "00010010", "00010010", "00010010", "00010010", "11101110", "11101110", "11101110", "11101110", "11101110", 
"11101110", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101100", "11101100", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101011", "11101011", "11101010", 
"11101010", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", "11100111", "11100110", "11100110", "11100110", "11100101", 
"11100101", "11100101", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100001", "11100001", "11100000", "11100000", "11100000", "11011111", "11011111", "11011110", "11011110", 
"11011101", "11011101", "11011100", "11011100", "11011011", "11011010", "11011010", "11011001", "11011000", "11011000", "11010111", "11010110", "11010110", "11010101", "11010100", "11010011", "11010011", "11010010", "11010001", "11010000", 
"11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001000", "11000111", "11000110", "11000101", "11000011", "11000010", "11000000", "10111111", "10111101", "10111011", "10111010", "10111000", "10110110", "10110100", 
"10110010", "10110000", "10101101", "10101011", "10101001", "10100110", "01010111", "01010100", "01010001", "01001110", "01001010", "01000110", "01000010", "00111110", "00111001", "00110100", "00101110", "00101000", "00100010", "00011100", 
"00010101", "00001110", "00000111", "00000000", "11111001", "11110011", "11101100", "11100110", "11100000", "11011010", "11010100", "11001111", "11001010", "11000101", "11000000", "10111100", "10111000", "10110101", "10110001", "10101110", 
"10101011", "10101001", "10100110", "01010111", "01010101", "01010011", "01010001", "01001111", "01001101", "01001011", "01001001", "01000111", "01000110", "01000100", "01000010", "01000001", "00111111", "00111110", "00111101", "00111011", 
"00111010", "00111001", "00111000", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00110000", "00101111", "00101110", "00101101", "00101100", "00101100", "00101011", "00101010", "00101001", "00101001", 
"00101000", "00101000", "00100111", "00100110", "00100110", "00100101", "00100101", "00100100", "00100100", "00100011", "00100011", "00100010", "00100010", "00100001", "00100001", "00100000", "00100000", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011001", "00011001", "00011001", "00011001", 
"00011000", "00011000", "00011000", "00011000", "00010111", "00010111", "00010111", "00010111", "00010111", "00010110", "00010110", "00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010101", "00010101", "00010101", 
"00010100", "00010100", "00010100", "00010100", "00010100", "00010100", "00010011", "00010011", "00010011", "00010011", "00010011", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101100", "11101100", "11101100", 
"11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101011", "11101011", "11101010", "11101010", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101001", "11101001", "11101000", 
"11101000", "11101000", "11101000", "11100111", "11100111", "11100111", "11100111", "11100110", "11100110", "11100110", "11100101", "11100101", "11100101", "11100101", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", 
"11100010", "11100010", "11100010", "11100001", "11100001", "11100000", "11100000", "11100000", "11011111", "11011111", "11011110", "11011110", "11011101", "11011101", "11011100", "11011100", "11011011", "11011011", "11011010", "11011010", 
"11011001", "11011000", "11011000", "11010111", "11010111", "11010110", "11010101", "11010100", "11010100", "11010011", "11010010", "11010001", "11010000", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", 
"11001000", "11000111", "11000110", "11000101", "11000011", "11000010", "11000001", "10111111", "10111110", "10111100", "10111010", "10111001", "10110111", "10110101", "10110011", "10110001", "10101111", "10101101", "10101011", "10101001", 
"10100110", "01010111", "01010101", "01010010", "01001111", "01001011", "01001000", "01000100", "01000000", "00111011", "00110110", "00110001", "00101100", "00100110", "00100000", "00011010", "00010100", "00001101", "00000111", "00000000", 
"11111010", "11110011", "11101101", "11100111", "11100001", "11011100", "11010110", "11010001", "11001100", "11000111", "11000011", "10111111", "10111011", "10110111", "10110100", "10110001", "10101110", "10101011", "10101001", "10100110", 
"01011000", "01010101", "01010011", "01010001", "01001111", "01001101", "01001100", "01001010", "01001000", "01000110", "01000101", "01000011", "01000010", "01000000", "00111111", "00111110", "00111100", "00111011", "00111010", "00111001", 
"00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101110", "00101101", "00101100", "00101011", "00101011", "00101010", "00101001", "00101001", "00101000", 
"00101000", "00100111", "00100110", "00100110", "00100101", "00100101", "00100100", "00100100", "00100011", "00100011", "00100010", "00100010", "00100010", "00100001", "00100001", "00100000", "00100000", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011010", "00011001", "00011001", "00011001", 
"00011001", "00011000", "00011000", "00011000", "00011000", "00011000", "00010111", "00010111", "00010111", "00010111", "00010111", "00010110", "00010110", "00010110", "00010110", "00010110", "00010101", "00010101", "00010101", "00010101", 
"00010101", "00010101", "00010100", "00010100", "00010100", "00010100", "00010100", "11101100", "11101100", "11101100", "11101100", "11101100", "11101100", "11101011", "11101011", "11101011", "11101011", "11101011", "11101011", "11101010", 
"11101010", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", "11100111", "11100110", "11100110", 
"11100110", "11100110", "11100101", "11100101", "11100101", "11100100", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100001", "11100001", "11100000", "11100000", "11100000", 
"11011111", "11011111", "11011110", "11011110", "11011110", "11011101", "11011101", "11011100", "11011100", "11011011", "11011011", "11011010", "11011010", "11011001", "11011000", "11011000", "11010111", "11010111", "11010110", "11010101", 
"11010101", "11010100", "11010011", "11010010", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000010", 
"11000001", "11000000", "10111110", "10111101", "10111011", "10111010", "10111000", "10110110", "10110100", "10110011", "10110001", "10101111", "10101101", "10101011", "10101000", "10100110", "01010111", "01010101", "01010010", "01001111", 
"01001100", "01001001", "01000101", "01000001", "00111101", "00111001", "00110100", "00101111", "00101010", "00100100", "00011111", "00011001", "00010011", "00001101", "00000110", "00000000", "11111010", "11110100", "11101110", "11101000", 
"11100011", "11011101", "11011000", "11010011", "11001110", "11001001", "11000101", "11000001", "10111101", "10111010", "10110110", "10110011", "10110000", "10101101", "10101011", "10101000", "10100110", "01011000", "01010110", "01010100", 
"01010010", "01010000", "01001110", "01001100", "01001010", "01001001", "01000111", "01000110", "01000100", "01000011", "01000001", "01000000", "00111111", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", 
"00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00110000", "00101111", "00101110", "00101101", "00101101", "00101100", "00101011", "00101011", "00101010", "00101001", "00101001", "00101000", "00101000", 
"00100111", "00100111", "00100110", "00100101", "00100101", "00100100", "00100100", "00100100", "00100011", "00100011", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00011111", "00011111", 
"00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011010", "00011001", "00011001", 
"00011001", "00011001", "00011000", "00011000", "00011000", "00011000", "00011000", "00010111", "00010111", "00010111", "00010111", "00010111", "00010110", "00010110", "00010110", "00010110", "00010110", "00010110", "00010101", "00010101", 
"00010101", "00010101", "00010101", "11101011", "11101011", "11101011", "11101011", "11101011", "11101011", "11101010", "11101010", "11101010", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101001", "11101001", 
"11101000", "11101000", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", "11100111", "11100110", "11100110", "11100110", "11100110", "11100101", "11100101", "11100101", "11100101", "11100100", "11100100", "11100100", 
"11100011", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100001", "11100001", "11100000", "11100000", "11100000", "11011111", "11011111", "11011111", "11011110", "11011110", "11011101", "11011101", "11011100", 
"11011100", "11011100", "11011011", "11011011", "11011010", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010110", "11010101", "11010101", "11010100", "11010011", "11010011", "11010010", "11010001", "11010000", 
"11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000001", "11000000", "10111111", "10111101", "10111100", "10111010", 
"10111001", "10110111", "10110110", "10110100", "10110010", "10110000", "10101110", "10101100", "10101010", "10101000", "10100110", "01011000", "01010101", "01010011", "01010000", "01001101", "01001010", "01000110", "01000011", "00111111", 
"00111011", "00110111", "00110010", "00101101", "00101000", "00100011", "00011101", "00011000", "00010010", "00001100", "00000110", "00000000", "11111010", "11110101", "11101111", "11101001", "11100100", "11011111", "11011001", "11010101", 
"11010000", "11001011", "11000111", "11000011", "10111111", "10111100", "10111000", "10110101", "10110010", "10110000", "10101101", "10101011", "10101000", "10100110", "01011000", "01010110", "01010100", "01010010", "01010000", "01001110", 
"01001101", "01001011", "01001010", "01001000", "01000110", "01000101", "01000100", "01000010", "01000001", "01000000", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", 
"00110100", "00110011", "00110010", "00110001", "00110001", "00110000", "00101111", "00101110", "00101110", "00101101", "00101100", "00101100", "00101011", "00101010", "00101010", "00101001", "00101001", "00101000", "00101000", "00100111", 
"00100111", "00100110", "00100110", "00100101", "00100101", "00100100", "00100100", "00100011", "00100011", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011110", "00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011010", "00011001", 
"00011001", "00011001", "00011001", "00011000", "00011000", "00011000", "00011000", "00011000", "00010111", "00010111", "00010111", "00010111", "00010111", "00010111", "00010110", "00010110", "00010110", "00010110", "00010110", "11101010", 
"11101010", "11101010", "11101010", "11101010", "11101010", "11101001", "11101001", "11101001", "11101001", "11101001", "11101001", "11101000", "11101000", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", "11100111", 
"11100110", "11100110", "11100110", "11100110", "11100101", "11100101", "11100101", "11100101", "11100100", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100010", "11100001", 
"11100001", "11100001", "11100000", "11100000", "11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011101", "11011101", "11011100", "11011100", "11011011", "11011011", "11011010", "11011010", "11011001", "11011001", 
"11011000", "11011000", "11010111", "11010111", "11010110", "11010110", "11010101", "11010100", "11010100", "11010011", "11010010", "11010010", "11010001", "11010000", "11001111", "11001111", "11001110", "11001101", "11001100", "11001011", 
"11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000000", "10111111", "10111110", "10111100", "10111011", "10111010", "10111000", "10110110", "10110101", "10110011", "10110010", 
"10110000", "10101110", "10101100", "10101010", "10101000", "10100110", "01011000", "01010101", "01010011", "01010000", "01001110", "01001011", "01001000", "01000100", "01000001", "00111101", "00111001", "00110101", "00110000", "00101011", 
"00100111", "00100001", "00011100", "00010111", "00010001", "00001011", "00000110", "00000000", "11111010", "11110101", "11110000", "11101010", "11100101", "11100000", "11011011", "11010110", "11010010", "11001101", "11001001", "11000101", 
"11000010", "10111110", "10111011", "10110111", "10110101", "10110010", "10101111", "10101101", "10101010", "10101000", "10100110", "01011000", "01010110", "01010100", "01010010", "01010001", "01001111", "01001101", "01001100", "01001010", 
"01001001", "01000111", "01000110", "01000100", "01000011", "01000010", "01000001", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", 
"00110011", "00110010", "00110001", "00110000", "00110000", "00101111", "00101110", "00101101", "00101101", "00101100", "00101100", "00101011", "00101010", "00101010", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", 
"00100110", "00100110", "00100101", "00100101", "00100100", "00100100", "00100100", "00100011", "00100011", "00100010", "00100010", "00100010", "00100001", "00100001", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011110", "00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011010", "00011010", 
"00011001", "00011001", "00011001", "00011001", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00010111", "00010111", "00010111", "00010111", "00010111", "11101010", "11101001", "11101001", "11101001", "11101001", 
"11101001", "11101000", "11101000", "11101000", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", "11100111", "11100110", "11100110", "11100110", "11100110", "11100110", "11100101", "11100101", "11100101", "11100101", 
"11100100", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100010", "11100001", "11100001", "11100001", "11100000", "11100000", "11100000", "11011111", "11011111", "11011110", 
"11011110", "11011110", "11011101", "11011101", "11011100", "11011100", "11011100", "11011011", "11011011", "11011010", "11011010", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010110", "11010110", "11010101", 
"11010100", "11010100", "11010011", "11010011", "11010010", "11010001", "11010000", "11010000", "11001111", "11001110", "11001101", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", 
"11000100", "11000011", "11000010", "11000001", "10111111", "10111110", "10111101", "10111100", "10111010", "10111001", "10110111", "10110110", "10110100", "10110011", "10110001", "10101111", "10101110", "10101100", "10101010", "10101000", 
"10100110", "01011000", "01010110", "01010011", "01010001", "01001110", "01001011", "01001001", "01000101", "01000010", "00111110", "00111011", "00110111", "00110011", "00101110", "00101010", "00100101", "00100000", "00011011", "00010110", 
"00010000", "00001011", "00000110", "00000000", "11111011", "11110101", "11110000", "11101011", "11100110", "11100001", "11011100", "11011000", "11010011", "11001111", "11001011", "11000111", "11000100", "11000000", "10111101", "10111010", 
"10110111", "10110100", "10110001", "10101111", "10101100", "10101010", "10101000", "10100110", "01011000", "01010110", "01010100", "01010011", "01010001", "01001111", "01001110", "01001100", "01001011", "01001001", "01001000", "01000110", 
"01000101", "01000100", "01000011", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110100", "00110011", "00110010", 
"00110001", "00110001", "00110000", "00101111", "00101110", "00101110", "00101101", "00101101", "00101100", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100110", 
"00100110", "00100101", "00100101", "00100100", "00100100", "00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011111", "00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", "00011010", 
"00011010", "00011001", "00011001", "00011001", "00011001", "00011001", "00011000", "00011000", "00011000", "00011000", "00011000", "11101001", "11101000", "11101000", "11101000", "11101000", "11101000", "11100111", "11100111", "11100111", 
"11100111", "11100111", "11100110", "11100110", "11100110", "11100110", "11100110", "11100101", "11100101", "11100101", "11100101", "11100100", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", "11100011", "11100010", 
"11100010", "11100010", "11100001", "11100001", "11100001", "11100001", "11100000", "11100000", "11100000", "11011111", "11011111", "11011111", "11011110", "11011110", "11011101", "11011101", "11011101", "11011100", "11011100", "11011100", 
"11011011", "11011011", "11011010", "11011010", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", "11010100", "11010011", "11010011", "11010010", "11010010", "11010001", 
"11010000", "11001111", "11001111", "11001110", "11001101", "11001100", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", 
"10111101", "10111100", "10111011", "10111010", "10111000", "10110111", "10110101", "10110100", "10110010", "10110001", "10101111", "10101101", "10101100", "10101010", "10101000", "10100110", "01011000", "01010110", "01010100", "01010001", 
"01001111", "01001100", "01001001", "01000110", "01000011", "01000000", "00111100", "00111001", "00110101", "00110001", "00101101", "00101000", "00100100", "00011111", "00011010", "00010101", "00010000", "00001011", "00000101", "00000000", 
"11111011", "11110110", "11110001", "11101100", "11100111", "11100010", "11011110", "11011001", "11010101", "11010001", "11001101", "11001001", "11000101", "11000010", "10111111", "10111100", "10111001", "10110110", "10110011", "10110001", 
"10101110", "10101100", "10101010", "10101000", "10100110", "01011000", "01010110", "01010101", "01010011", "01010001", "01010000", "01001110", "01001101", "01001011", "01001010", "01001000", "01000111", "01000110", "01000101", "01000011", 
"01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110101", "00110100", "00110011", "00110010", "00110010", "00110001", 
"00110000", "00101111", "00101111", "00101110", "00101110", "00101101", "00101100", "00101100", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100110", "00100110", 
"00100101", "00100101", "00100101", "00100100", "00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011111", "00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", 
"00011010", "00011001", "00011001", "00011001", "00011001", "00011001", "00011001", "11101000", "11100111", "11100111", "11100111", "11100111", "11100111", "11100111", "11100110", "11100110", "11100110", "11100110", "11100101", "11100101", 
"11100101", "11100101", "11100101", "11100100", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100001", "11100001", "11100001", "11100001", "11100000", "11100000", 
"11100000", "11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011101", "11011101", "11011101", "11011100", "11011100", "11011011", "11011011", "11011011", "11011010", "11011010", "11011001", "11011001", "11011000", 
"11011000", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", "11010100", "11010100", "11010011", "11010010", "11010010", "11010001", "11010001", "11010000", "11001111", "11001110", "11001110", "11001101", "11001100", 
"11001011", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111011", "10111010", "10111001", "10111000", 
"10110110", "10110101", "10110011", "10110010", "10110000", "10101111", "10101101", "10101011", "10101010", "10101000", "10100110", "01011000", "01010110", "01010100", "01010010", "01001111", "01001101", "01001010", "01000111", "01000100", 
"01000001", "00111110", "00111011", "00110111", "00110011", "00101111", "00101011", "00100111", "00100010", "00011110", "00011001", "00010100", "00001111", "00001010", "00000101", "00000000", "11111011", "11110110", "11110001", "11101101", 
"11101000", "11100011", "11011111", "11011011", "11010110", "11010010", "11001111", "11001011", "11000111", "11000100", "11000001", "10111101", "10111010", "10111000", "10110101", "10110011", "10110000", "10101110", "10101100", "10101010", 
"10101000", "10100110", "01011000", "01010110", "01010101", "01010011", "01010010", "01010000", "01001111", "01001101", "01001100", "01001010", "01001001", "01001000", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", 
"01000000", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110101", "00110100", "00110011", "00110010", "00110010", "00110001", "00110000", "00110000", 
"00101111", "00101111", "00101110", "00101101", "00101101", "00101100", "00101100", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100110", "00100110", "00100110", 
"00100101", "00100101", "00100100", "00100100", "00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011111", "00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011011", "00011010", "00011010", "00011010", 
"00011010", "00011010", "00011001", "11100111", "11100111", "11100110", "11100110", "11100110", "11100110", "11100110", "11100101", "11100101", "11100101", "11100101", "11100100", "11100100", "11100100", "11100100", "11100100", "11100011", 
"11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100001", "11100001", "11100001", "11100001", "11100000", "11100000", "11100000", "11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011101", 
"11011101", "11011101", "11011100", "11011100", "11011100", "11011011", "11011011", "11011010", "11011010", "11011010", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", 
"11010100", "11010100", "11010011", "11010011", "11010010", "11010001", "11010001", "11010000", "11010000", "11001111", "11001110", "11001110", "11001101", "11001100", "11001011", "11001011", "11001010", "11001001", "11001000", "11000111", 
"11000110", "11000101", "11000100", "11000100", "11000011", "11000010", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111000", "10110111", "10110110", "10110100", "10110011", "10110001", "10110000", 
"10101110", "10101101", "10101011", "10101010", "10101000", "10100110", "01011000", "01010110", "01010100", "01010010", "01010000", "01001101", "01001011", "01001000", "01000110", "01000011", "00111111", "00111100", "00111001", "00110101", 
"00110001", "00101110", "00101010", "00100101", "00100001", "00011101", "00011000", "00010011", "00001111", "00001010", "00000101", "00000000", "11111011", "11110111", "11110010", "11101101", "11101001", "11100100", "11100000", "11011100", 
"11011000", "11010100", "11010000", "11001100", "11001001", "11000110", "11000010", "10111111", "10111100", "10111010", "10110111", "10110100", "10110010", "10110000", "10101110", "10101100", "10101010", "10101000", "10100110", "01011000", 
"01010111", "01010101", "01010011", "01010010", "01010000", "01001111", "01001110", "01001100", "01001011", "01001010", "01001000", "01000111", "01000110", "01000101", "01000100", "01000010", "01000001", "01000000", "00111111", "00111110", 
"00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110110", "00110101", "00110100", "00110011", "00110011", "00110010", "00110001", "00110001", "00110000", "00101111", "00101111", 
"00101110", "00101110", "00101101", "00101101", "00101100", "00101100", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", 
"00100101", "00100100", "00100100", "00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011111", "00011110", "00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011100", "00011011", "00011011", "00011011", "00011011", "00011011", "00011010", "11100110", 
"11100110", "11100101", "11100101", "11100101", "11100101", "11100101", "11100100", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100010", "11100001", "11100001", 
"11100001", "11100001", "11100000", "11100000", "11100000", "11100000", "11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011101", "11011101", "11011101", "11011100", "11011100", "11011100", "11011011", "11011011", 
"11011010", "11011010", "11011010", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", "11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010001", 
"11010001", "11010000", "11001111", "11001111", "11001110", "11001101", "11001101", "11001100", "11001011", "11001010", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000010", 
"11000001", "11000000", "10111111", "10111110", "10111100", "10111011", "10111010", "10111001", "10111000", "10110110", "10110101", "10110100", "10110010", "10110001", "10110000", "10101110", "10101101", "10101011", "10101001", "10101000", 
"10100110", "01011000", "01010110", "01010100", "01010010", "01010000", "01001110", "01001100", "01001001", "01000110", "01000100", "01000001", "00111110", "00111010", "00110111", "00110100", "00110000", "00101100", "00101000", "00100100", 
"00100000", "00011100", "00010111", "00010011", "00001110", "00001001", "00000101", "00000000", "11111011", "11110111", "11110010", "11101110", "11101010", "11100101", "11100001", "11011101", "11011001", "11010101", "11010010", "11001110", 
"11001011", "11000111", "11000100", "11000001", "10111110", "10111011", "10111001", "10110110", "10110100", "10110010", "10101111", "10101101", "10101011", "10101010", "10101000", "10100110", "01011000", "01010111", "01010101", "01010100", 
"01010010", "01010001", "01001111", "01001110", "01001101", "01001011", "01001010", "01001001", "01001000", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", 
"00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110110", "00110110", "00110101", "00110100", "00110100", "00110011", "00110010", "00110010", "00110001", "00110000", "00110000", "00101111", "00101111", "00101110", 
"00101101", "00101101", "00101100", "00101100", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100101", "00100101", 
"00100101", "00100100", "00100100", "00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011111", "00011110", "00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011101", "00011100", "00011100", "00011100", "00011100", "00011100", "00011011", "11100101", "11100101", "11100100", "11100100", "11100100", 
"11100100", "11100100", "11100011", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100010", "11100001", "11100001", "11100001", "11100001", "11100000", "11100000", "11100000", "11100000", "11011111", "11011111", 
"11011111", "11011110", "11011110", "11011110", "11011101", "11011101", "11011101", "11011100", "11011100", "11011100", "11011011", "11011011", "11011011", "11011010", "11011010", "11011001", "11011001", "11011001", "11011000", "11011000", 
"11010111", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", "11010100", "11010100", "11010011", "11010011", "11010010", "11010001", "11010001", "11010000", "11010000", "11001111", "11001110", "11001110", "11001101", 
"11001100", "11001100", "11001011", "11001010", "11001010", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", 
"10111011", "10111010", "10111000", "10110111", "10110110", "10110101", "10110011", "10110010", "10110001", "10101111", "10101110", "10101100", "10101011", "10101001", "10101000", "10100110", "01011000", "01010110", "01010101", "01010011", 
"01010001", "01001110", "01001100", "01001010", "01000111", "01000101", "01000010", "00111111", "00111100", "00111001", "00110101", "00110010", "00101110", "00101011", "00100111", "00100011", "00011111", "00011011", "00010110", "00010010", 
"00001110", "00001001", "00000101", "00000000", "11111100", "11110111", "11110011", "11101111", "11101010", "11100110", "11100010", "11011110", "11011010", "11010111", "11010011", "11001111", "11001100", "11001001", "11000110", "11000011", 
"11000000", "10111101", "10111010", "10111000", "10110110", "10110011", "10110001", "10101111", "10101101", "10101011", "10101001", "10101000", "10100110", "01011000", "01010111", "01010101", "01010100", "01010010", "01010001", "01010000", 
"01001110", "01001101", "01001100", "01001011", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", 
"00111010", "00111001", "00111000", "00110111", "00110111", "00110110", "00110101", "00110100", "00110100", "00110011", "00110010", "00110010", "00110001", "00110001", "00110000", "00101111", "00101111", "00101110", "00101110", "00101101", 
"00101101", "00101100", "00101100", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100101", "00100101", "00100101", 
"00100100", "00100100", "00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011111", "00011110", "00011110", "00011110", "00011110", "00011101", "00011101", "00011101", "00011101", "00011100", "00011100", "11100100", "11100100", "11100100", "11100011", "11100011", "11100011", "11100011", "11100010", "11100010", 
"11100010", "11100010", "11100001", "11100001", "11100001", "11100001", "11100000", "11100000", "11100000", "11100000", "11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011110", "11011101", "11011101", "11011101", 
"11011100", "11011100", "11011100", "11011011", "11011011", "11011011", "11011010", "11011010", "11011001", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", 
"11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010001", "11010001", "11010000", "11001111", "11001111", "11001110", "11001110", "11001101", "11001100", "11001100", "11001011", "11001010", "11001001", "11001001", 
"11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110101", 
"10110100", "10110011", "10110010", "10110000", "10101111", "10101110", "10101100", "10101011", "10101001", "10101000", "10100110", "01011000", "01010111", "01010101", "01010011", "01010001", "01001111", "01001101", "01001010", "01001000", 
"01000110", "01000011", "01000000", "00111101", "00111010", "00110111", "00110100", "00110001", "00101101", "00101001", "00100110", "00100010", "00011110", "00011010", "00010110", "00010001", "00001101", "00001001", "00000100", "00000000", 
"11111100", "11111000", "11110011", "11101111", "11101011", "11100111", "11100011", "11011111", "11011100", "11011000", "11010100", "11010001", "11001110", "11001010", "11000111", "11000100", "11000001", "10111111", "10111100", "10111010", 
"10110111", "10110101", "10110011", "10110001", "10101111", "10101101", "10101011", "10101001", "10101000", "10100110", "01011000", "01010111", "01010101", "01010100", "01010011", "01010001", "01010000", "01001111", "01001101", "01001100", 
"01001011", "01001010", "01001001", "01001000", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111010", "00111001", 
"00111000", "00110111", "00110111", "00110110", "00110101", "00110101", "00110100", "00110011", "00110011", "00110010", "00110001", "00110001", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101101", "00101101", 
"00101100", "00101100", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", "00100101", "00100100", 
"00100100", "00100100", "00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011111", "00011110", "00011110", "00011110", "00011110", "00011101", "00011101", "11100011", "11100011", "11100011", "11100010", "11100010", "11100010", "11100010", "11100001", "11100001", "11100001", "11100001", "11100000", "11100000", 
"11100000", "11100000", "11011111", "11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011101", "11011101", "11011101", "11011100", "11011100", "11011100", "11011100", "11011011", "11011011", "11011010", "11011010", 
"11011010", "11011001", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", "11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010001", 
"11010001", "11010000", "11010000", "11001111", "11001111", "11001110", "11001101", "11001101", "11001100", "11001011", "11001011", "11001010", "11001001", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", 
"11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110001", "10110000", "10101111", 
"10101101", "10101100", "10101011", "10101001", "10101000", "10100110", "01011000", "01010111", "01010101", "01010011", "01010001", "01001111", "01001101", "01001011", "01001001", "01000110", "01000100", "01000001", "00111111", "00111100", 
"00111001", "00110110", "00110010", "00101111", "00101100", "00101000", "00100100", "00100001", "00011101", "00011001", "00010101", "00010001", "00001101", "00001000", "00000100", "00000000", "11111100", "11111000", "11110100", "11110000", 
"11101100", "11101000", "11100100", "11100000", "11011101", "11011001", "11010110", "11010010", "11001111", "11001100", "11001001", "11000110", "11000011", "11000000", "10111110", "10111011", "10111001", "10110110", "10110100", "10110010", 
"10110000", "10101110", "10101101", "10101011", "10101001", "10101000", "10100110", "01011000", "01010111", "01010110", "01010100", "01010011", "01010010", "01010000", "01001111", "01001110", "01001101", "01001011", "01001010", "01001001", 
"01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", 
"00110111", "00110110", "00110101", "00110101", "00110100", "00110011", "00110011", "00110010", "00110010", "00110001", "00110001", "00110000", "00101111", "00101111", "00101110", "00101110", "00101101", "00101101", "00101100", "00101100", 
"00101100", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", "00100101", "00100101", "00100100", 
"00100100", "00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", 
"00011111", "00011110", "00011110", "11100010", "11100010", "11100010", "11100001", "11100001", "11100001", "11100001", "11100000", "11100000", "11100000", "11100000", "11011111", "11011111", "11011111", "11011111", "11011110", "11011110", 
"11011110", "11011110", "11011101", "11011101", "11011101", "11011100", "11011100", "11011100", "11011011", "11011011", "11011011", "11011010", "11011010", "11011010", "11011001", "11011001", "11011001", "11011000", "11011000", "11010111", 
"11010111", "11010111", "11010110", "11010110", "11010101", "11010101", "11010100", "11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010001", "11010001", "11010000", "11001111", "11001111", "11001110", "11001110", 
"11001101", "11001101", "11001100", "11001011", "11001011", "11001010", "11001001", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "10111111", 
"10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110011", "10110010", "10110001", "10110000", "10101110", "10101101", "10101100", "10101010", "10101001", "10101000", 
"10100110", "01011000", "01010111", "01010101", "01010011", "01010010", "01010000", "01001110", "01001100", "01001010", "01000111", "01000101", "01000010", "01000000", "00111101", "00111010", "00110111", "00110100", "00110001", "00101110", 
"00101010", "00100111", "00100011", "00100000", "00011100", "00011000", "00010100", "00010000", "00001100", "00001000", "00000100", "00000000", "11111100", "11111000", "11110100", "11110000", "11101100", "11101001", "11100101", "11100001", 
"11011110", "11011010", "11010111", "11010011", "11010000", "11001101", "11001010", "11000111", "11000100", "11000010", "10111111", "10111101", "10111010", "10111000", "10110110", "10110100", "10110010", "10110000", "10101110", "10101100", 
"10101011", "10101001", "10101000", "10100110", "01011000", "01010111", "01010110", "01010100", "01010011", "01010010", "01010001", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01000111", "01000110", 
"01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110111", "00110110", 
"00110101", "00110101", "00110100", "00110100", "00110011", "00110010", "00110010", "00110001", "00110001", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101101", "00101101", "00101100", "00101100", "00101011", 
"00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", "00100101", "00100101", "00100100", "00100100", 
"00100100", "00100011", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "00100000", "00011111", "00011111", "00011111", "11100001", 
"11100001", "11100001", "11100001", "11100000", "11100000", "11100000", "11100000", "11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011110", "11011101", "11011101", "11011101", "11011101", "11011100", "11011100", 
"11011100", "11011011", "11011011", "11011011", "11011010", "11011010", "11011010", "11011001", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", "11010101", 
"11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010001", "11010001", "11010000", "11010000", "11001111", "11001111", "11001110", "11001110", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", 
"11001001", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111010", 
"10111001", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10101111", "10101110", "10101101", "10101100", "10101010", "10101001", "10101000", "10100110", "01011000", "01010111", "01010101", "01010100", 
"01010010", "01010000", "01001110", "01001100", "01001010", "01001000", "01000110", "01000011", "01000001", "00111110", "00111100", "00111001", "00110110", "00110011", "00110000", "00101101", "00101001", "00100110", "00100010", "00011111", 
"00011011", "00010111", "00010100", "00010000", "00001100", "00001000", "00000100", "00000000", "11111100", "11111000", "11110101", "11110001", "11101101", "11101001", "11100110", "11100010", "11011111", "11011011", "11011000", "11010101", 
"11010001", "11001110", "11001011", "11001001", "11000110", "11000011", "11000001", "10111110", "10111100", "10111010", "10110111", "10110101", "10110011", "10110001", "10110000", "10101110", "10101100", "10101011", "10101001", "10101000", 
"10100110", "01011000", "01010111", "01010110", "01010101", "01010011", "01010010", "01010001", "01010000", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", 
"01000011", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111001", "00111001", "00111000", "00110111", "00110111", "00110110", "00110110", "00110101", 
"00110100", "00110100", "00110011", "00110011", "00110010", "00110001", "00110001", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101101", "00101101", "00101101", "00101100", "00101100", "00101011", "00101011", 
"00101010", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", "00100101", "00100101", "00100100", "00100100", "00100100", 
"00100100", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "00100001", "00100000", "00100000", "00100000", "11100000", "11100000", "11100000", "11100000", "11011111", 
"11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011110", "11011101", "11011101", "11011101", "11011100", "11011100", "11011100", "11011100", "11011011", "11011011", "11011011", "11011010", "11011010", "11011010", 
"11011001", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010110", "11010101", "11010101", "11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", 
"11010001", "11010001", "11010000", "11010000", "11001111", "11001111", "11001110", "11001101", "11001101", "11001100", "11001100", "11001011", "11001010", "11001010", "11001001", "11001001", "11001000", "11000111", "11000111", "11000110", 
"11000101", "11000100", "11000100", "11000011", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", 
"10110011", "10110010", "10110000", "10101111", "10101110", "10101101", "10101011", "10101010", "10101001", "10101000", "10100110", "01011000", "01010111", "01010101", "01010100", "01010010", "01010000", "01001111", "01001101", "01001011", 
"01001001", "01000110", "01000100", "01000010", "00111111", "00111101", "00111010", "00110111", "00110101", "00110010", "00101111", "00101011", "00101000", "00100101", "00100001", "00011110", "00011010", "00010111", "00010011", "00001111", 
"00001011", "00001000", "00000100", "00000000", "11111100", "11111001", "11110101", "11110001", "11101110", "11101010", "11100110", "11100011", "11100000", "11011100", "11011001", "11010110", "11010011", "11010000", "11001101", "11001010", 
"11000111", "11000101", "11000010", "11000000", "10111101", "10111011", "10111001", "10110111", "10110101", "10110011", "10110001", "10101111", "10101110", "10101100", "10101010", "10101001", "10101000", "10100110", "01011000", "01010111", 
"01010110", "01010101", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000010", 
"01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111001", "00111001", "00111000", "00110111", "00110111", "00110110", "00110110", "00110101", "00110100", "00110100", 
"00110011", "00110011", "00110010", "00110010", "00110001", "00110001", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101101", "00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101010", 
"00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100110", "00100101", "00100101", "00100101", "00100100", "00100100", "00100100", 
"00100011", "00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100010", "00100001", "00100001", "00100001", "11011111", "11011111", "11011111", "11011111", "11011110", "11011110", "11011110", "11011110", "11011101", 
"11011101", "11011101", "11011101", "11011100", "11011100", "11011100", "11011011", "11011011", "11011011", "11011010", "11011010", "11011010", "11011010", "11011001", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", 
"11010111", "11010110", "11010110", "11010110", "11010101", "11010101", "11010100", "11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010001", "11010001", "11010000", "11010000", "11001111", "11001111", "11001110", 
"11001110", "11001101", "11001101", "11001100", "11001100", "11001011", "11001010", "11001010", "11001001", "11001001", "11001000", "11000111", "11000111", "11000110", "11000101", "11000100", "11000100", "11000011", "11000010", "11000001", 
"11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", 
"10101101", "10101011", "10101010", "10101001", "10101000", "10100110", "01011000", "01010111", "01010110", "01010100", "01010010", "01010001", "01001111", "01001101", "01001011", "01001001", "01000111", "01000101", "01000011", "01000000", 
"00111110", "00111011", "00111001", "00110110", "00110011", "00110000", "00101101", "00101010", "00100111", "00100100", "00100000", "00011101", "00011010", "00010110", "00010010", "00001111", "00001011", "00000111", "00000100", "00000000", 
"11111100", "11111001", "11110101", "11110010", "11101110", "11101011", "11100111", "11100100", "11100000", "11011101", "11011010", "11010111", "11010100", "11010001", "11001110", "11001011", "11001001", "11000110", "11000011", "11000001", 
"10111111", "10111100", "10111010", "10111000", "10110110", "10110100", "10110010", "10110001", "10101111", "10101101", "10101100", "10101010", "10101001", "10101000", "10100110", "01011001", "01010111", "01010110", "01010101", "01010100", 
"01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", 
"00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110110", "00110110", "00110101", "00110101", "00110100", "00110011", "00110011", 
"00110010", "00110010", "00110001", "00110001", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101110", "00101101", "00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101010", "00101010", 
"00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00100111", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", "00100101", "00100101", "00100100", "00100100", "00100100", "00100100", 
"00100011", "00100011", "00100011", "00100010", "00100010", "00100010", "00100010", "11011111", "11011110", "11011110", "11011110", "11011110", "11011101", "11011101", "11011101", "11011100", "11011100", "11011100", "11011100", "11011011", 
"11011011", "11011011", "11011010", "11011010", "11011010", "11011001", "11011001", "11011001", "11011001", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010110", "11010101", "11010101", "11010100", 
"11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010010", "11010001", "11010001", "11010000", "11010000", "11001111", "11001111", "11001110", "11001110", "11001101", "11001101", "11001100", "11001011", "11001011", 
"11001010", "11001010", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "10111111", "10111110", "10111110", "10111101", 
"10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101100", "10101011", "10101010", "10101001", "10100111", 
"10100110", "01011000", "01010111", "01010110", "01010100", "01010011", "01010001", "01001111", "01001110", "01001100", "01001010", "01001000", "01000110", "01000100", "01000001", "00111111", "00111101", "00111010", "00110111", "00110101", 
"00110010", "00101111", "00101100", "00101001", "00100110", "00100011", "00100000", "00011100", "00011001", "00010101", "00010010", "00001110", "00001011", "00000111", "00000100", "00000000", "11111100", "11111001", "11110101", "11110010", 
"11101111", "11101011", "11101000", "11100100", "11100001", "11011110", "11011011", "11011000", "11010101", "11010010", "11001111", "11001100", "11001010", "11000111", "11000101", "11000010", "11000000", "10111110", "10111100", "10111010", 
"10111000", "10110110", "10110100", "10110010", "10110000", "10101111", "10101101", "10101100", "10101010", "10101001", "10100111", "10100110", "01011001", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010000", 
"01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111110", 
"00111110", "00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110010", 
"00110010", "00110001", "00110001", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101101", "00101101", "00101101", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "00101010", "00101010", 
"00101001", "00101001", "00101000", "00101000", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", "00100101", "00100101", "00100100", "00100100", "00100100", "00100100", "00100011", 
"00100011", "00100011", "00100011", "11011110", "11011101", "11011101", "11011101", "11011101", "11011100", "11011100", "11011100", "11011100", "11011011", "11011011", "11011011", "11011010", "11011010", "11011010", "11011001", "11011001", 
"11011001", "11011000", "11011000", "11011000", "11011000", "11010111", "11010111", "11010110", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", 
"11010001", "11010001", "11010000", "11010000", "11001111", "11001111", "11001110", "11001110", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001001", "11001000", "11001000", "11000111", 
"11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", 
"10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10100111", "10100110", "01011001", "01010111", "01010110", "01010100", 
"01010011", "01010001", "01010000", "01001110", "01001100", "01001010", "01001000", "01000110", "01000100", "01000010", "01000000", "00111110", "00111011", "00111001", "00110110", "00110100", "00110001", "00101110", "00101011", "00101000", 
"00100101", "00100010", "00011111", "00011100", "00011000", "00010101", "00010001", "00001110", "00001011", "00000111", "00000100", "00000000", "11111101", "11111001", "11110110", "11110010", "11101111", "11101100", "11101000", "11100101", 
"11100010", "11011111", "11011100", "11011001", "11010110", "11010011", "11010000", "11001110", "11001011", "11001000", "11000110", "11000100", "11000001", "10111111", "10111101", "10111011", "10111001", "10110111", "10110101", "10110011", 
"10110010", "10110000", "10101110", "10101101", "10101011", "10101010", "10101001", "10100111", "10100110", "01011001", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", 
"01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111101", "00111101", 
"00111100", "00111011", "00111011", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", "00110001", 
"00110001", "00110000", "00110000", "00101111", "00101111", "00101111", "00101110", "00101110", "00101101", "00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "00101010", "00101010", "00101001", 
"00101001", "00101000", "00101000", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", "00100101", "00100101", "00100101", "00100100", "00100100", "00100100", "00100100", "11011101", 
"11011100", "11011100", "11011100", "11011100", "11011011", "11011011", "11011011", "11011011", "11011010", "11011010", "11011010", "11011001", "11011001", "11011001", "11011000", "11011000", "11011000", "11011000", "11010111", "11010111", 
"11010110", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", "11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010001", "11010001", "11010001", "11010000", "11010000", "11001111", "11001111", 
"11001110", "11001110", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", 
"11000011", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", 
"10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10100111", "10100110", "01011001", "01010111", "01010110", "01010101", "01010011", "01010010", "01010000", "01001110", "01001101", 
"01001011", "01001001", "01000111", "01000101", "01000011", "01000001", "00111111", "00111100", "00111010", "00111000", "00110101", "00110010", "00110000", "00101101", "00101010", "00100111", "00100100", "00100001", "00011110", "00011011", 
"00011000", "00010100", "00010001", "00001110", "00001010", "00000111", "00000011", "00000000", "11111101", "11111001", "11110110", "11110011", "11101111", "11101100", "11101001", "11100110", "11100011", "11100000", "11011101", "11011010", 
"11010111", "11010100", "11010001", "11001111", "11001100", "11001010", "11000111", "11000101", "11000011", "11000000", "10111110", "10111100", "10111010", "10111000", "10110110", "10110101", "10110011", "10110001", "10110000", "10101110", 
"10101101", "10101011", "10101010", "10101001", "10100111", "10100110", "01011001", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", 
"01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", 
"00111011", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", "00110001", "00110001", "00110000", 
"00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101110", "00101101", "00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "00101010", "00101001", "00101001", "00101001", 
"00101000", "00101000", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100101", "00100101", "00100101", "00100101", "00100100", "11011100", "11011100", "11011011", "11011011", "11011011", 
"11011011", "11011010", "11011010", "11011010", "11011001", "11011001", "11011001", "11011000", "11011000", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", 
"11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010010", "11010001", "11010001", "11010000", "11010000", "11010000", "11001111", "11001111", "11001110", "11001110", "11001101", "11001101", "11001100", "11001100", 
"11001011", "11001011", "11001010", "11001010", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", 
"10111110", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", 
"10101100", "10101011", "10101010", "10101001", "10100111", "10100110", "01011001", "01010111", "01010110", "01010101", "01010011", "01010010", "01010000", "01001111", "01001101", "01001011", "01001010", "01001000", "01000110", "01000100", 
"01000010", "01000000", "00111101", "00111011", "00111001", "00110110", "00110100", "00110001", "00101111", "00101100", "00101001", "00100110", "00100011", "00100000", "00011101", "00011010", "00010111", "00010100", "00010001", "00001101", 
"00001010", "00000111", "00000011", "00000000", "11111101", "11111001", "11110110", "11110011", "11110000", "11101101", "11101010", "11100110", "11100011", "11100000", "11011110", "11011011", "11011000", "11010101", "11010010", "11010000", 
"11001101", "11001011", "11001000", "11000110", "11000100", "11000010", "10111111", "10111101", "10111011", "10111010", "10111000", "10110110", "10110100", "10110011", "10110001", "10101111", "10101110", "10101101", "10101011", "10101010", 
"10101001", "10100111", "10100110", "01011001", "01011000", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001001", 
"01001000", "01000111", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111100", "00111011", "00111011", "00111010", 
"00111001", "00111001", "00111000", "00111000", "00110111", "00110111", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", "00110010", "00110001", "00110001", "00110000", "00110000", 
"00101111", "00101111", "00101111", "00101110", "00101110", "00101101", "00101101", "00101101", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", 
"00101000", "00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "00100110", "00100110", "00100101", "11011011", "11011011", "11011010", "11011010", "11011010", "11011010", "11011001", "11011001", "11011001", 
"11011000", "11011000", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", 
"11010001", "11010001", "11010001", "11010000", "11010000", "11001111", "11001111", "11001110", "11001110", "11001110", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", "11001001", "11001001", "11001000", 
"11001000", "11000111", "11000111", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111100", "10111100", "10111011", 
"10111010", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101000", "10100111", 
"10100110", "01011001", "01010111", "01010110", "01010101", "01010011", "01010010", "01010001", "01001111", "01001101", "01001100", "01001010", "01001000", "01000110", "01000101", "01000011", "01000001", "00111110", "00111100", "00111010", 
"00111000", "00110101", "00110011", "00110000", "00101110", "00101011", "00101000", "00100101", "00100010", "00100000", "00011101", "00011010", "00010110", "00010011", "00010000", "00001101", "00001010", "00000111", "00000011", "00000000", 
"11111101", "11111010", "11110111", "11110011", "11110000", "11101101", "11101010", "11100111", "11100100", "11100001", "11011110", "11011100", "11011001", "11010110", "11010011", "11010001", "11001110", "11001100", "11001010", "11000111", 
"11000101", "11000011", "11000001", "10111111", "10111101", "10111011", "10111001", "10110111", "10110101", "10110100", "10110010", "10110001", "10101111", "10101110", "10101100", "10101011", "10101010", "10101001", "10100111", "10100110", 
"01011001", "01011000", "01010111", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", 
"01000110", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111100", "00111011", "00111011", "00111010", "00111001", "00111001", 
"00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", "00110001", "00110001", "00110000", "00110000", "00110000", "00101111", 
"00101111", "00101110", "00101110", "00101110", "00101101", "00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", 
"00101000", "00101000", "00100111", "00100111", "00100111", "00100110", "00100110", "11011010", "11011010", "11011010", "11011001", "11011001", "11011001", "11011000", "11011000", "11011000", "11011000", "11010111", "11010111", "11010111", 
"11010110", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", "11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010010", "11010001", "11010001", "11010000", "11010000", "11010000", "11001111", 
"11001111", "11001110", "11001110", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000101", "11000101", 
"11000100", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110110", 
"10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101001", "10101000", "10100111", "10100110", "01011001", "01010111", "01010110", "01010101", 
"01010100", "01010010", "01010001", "01001111", "01001110", "01001100", "01001011", "01001001", "01000111", "01000101", "01000011", "01000001", "00111111", "00111101", "00111011", "00111001", "00110110", "00110100", "00110010", "00101111", 
"00101101", "00101010", "00100111", "00100100", "00100010", "00011111", "00011100", "00011001", "00010110", "00010011", "00010000", "00001101", "00001001", "00000110", "00000011", "00000000", "11111101", "11111010", "11110111", "11110100", 
"11110001", "11101110", "11101011", "11101000", "11100101", "11100010", "11011111", "11011100", "11011010", "11010111", "11010100", "11010010", "11001111", "11001101", "11001011", "11001000", "11000110", "11000100", "11000010", "11000000", 
"10111110", "10111100", "10111010", "10111000", "10110111", "10110101", "10110011", "10110010", "10110000", "10101111", "10101110", "10101100", "10101011", "10101010", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", 
"01010110", "01010101", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000101", "01000101", 
"01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111100", "00111011", "00111011", "00111010", "00111001", "00111001", "00111000", "00111000", 
"00110111", "00110111", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", "00110001", "00110001", "00110001", "00110000", "00110000", "00101111", "00101111", "00101111", 
"00101110", "00101110", "00101101", "00101101", "00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00101000", 
"00101000", "00100111", "00100111", "11011001", "11011001", "11011001", "11011000", "11011000", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", 
"11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", "11010001", "11010001", "11010001", "11010000", "11010000", "11001111", "11001111", "11001111", "11001110", "11001110", "11001101", "11001101", "11001100", 
"11001100", "11001011", "11001011", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000010", "11000010", "11000001", 
"11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", 
"10110000", "10101111", "10101111", "10101110", "10101101", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010110", "01010101", "01010100", "01010010", "01010001", "01010000", "01001110", 
"01001101", "01001011", "01001001", "01001000", "01000110", "01000100", "01000010", "01000000", "00111110", "00111100", "00111010", "00111000", "00110101", "00110011", "00110001", "00101110", "00101100", "00101001", "00100110", "00100100", 
"00100001", "00011110", "00011011", "00011000", "00010101", "00010010", "00001111", "00001100", "00001001", "00000110", "00000011", "00000000", "11111101", "11111010", "11110111", "11110100", "11110001", "11101110", "11101011", "11101000", 
"11100101", "11100011", "11100000", "11011101", "11011010", "11011000", "11010101", "11010011", "11010000", "11001110", "11001100", "11001001", "11000111", "11000101", "11000011", "11000001", "10111111", "10111101", "10111011", "10111010", 
"10111000", "10110110", "10110101", "10110011", "10110010", "10110000", "10101111", "10101101", "10101100", "10101011", "10101010", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", 
"01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000011", 
"01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110111", 
"00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", "00110010", "00110001", "00110001", "00110000", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", 
"00101110", "00101101", "00101101", "00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "00101010", "00101010", "00101001", "00101001", "00101001", "00101000", "00101000", "00101000", "11011000", 
"11011000", "11011000", "11011000", "11010111", "11010111", "11010111", "11010110", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", "11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", 
"11010010", "11010001", "11010001", "11010000", "11010000", "11010000", "11001111", "11001111", "11001110", "11001110", "11001110", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001001", 
"11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", 
"10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", 
"10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010110", "01010101", "01010100", "01010011", "01010001", "01010000", "01001110", "01001101", "01001011", "01001010", "01001000", "01000110", 
"01000101", "01000011", "01000001", "00111111", "00111101", "00111011", "00111001", "00110111", "00110100", "00110010", "00110000", "00101101", "00101011", "00101000", "00100110", "00100011", "00100000", "00011101", "00011011", "00011000", 
"00010101", "00010010", "00001111", "00001100", "00001001", "00000110", "00000011", "00000000", "11111101", "11111010", "11110111", "11110100", "11110001", "11101110", "11101100", "11101001", "11100110", "11100011", "11100001", "11011110", 
"11011011", "11011001", "11010110", "11010100", "11010001", "11001111", "11001101", "11001010", "11001000", "11000110", "11000100", "11000010", "11000000", "10111110", "10111100", "10111011", "10111001", "10110111", "10110110", "10110100", 
"10110011", "10110001", "10110000", "10101110", "10101101", "10101100", "10101011", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", 
"01010000", "01001111", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", 
"01000000", "01000000", "00111111", "00111111", "00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", 
"00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110011", "00110010", "00110010", "00110001", "00110001", "00110001", "00110000", "00110000", "00101111", "00101111", "00101111", "00101110", "00101110", "00101110", 
"00101101", "00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101011", "00101011", "00101010", "00101010", "00101010", "00101001", "00101001", "00101001", "11011000", "11010111", "11010111", "11010111", "11010110", 
"11010110", "11010110", "11010101", "11010101", "11010101", "11010101", "11010100", "11010100", "11010100", "11010011", "11010011", "11010010", "11010010", "11010010", "11010001", "11010001", "11010001", "11010000", "11010000", "11001111", 
"11001111", "11001111", "11001110", "11001110", "11001101", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", 
"11000110", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", 
"10111000", "10111000", "10110111", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", 
"10100110", "01011001", "01011000", "01010111", "01010101", "01010100", "01010011", "01010010", "01010000", "01001111", "01001101", "01001100", "01001010", "01001001", "01000111", "01000101", "01000100", "01000010", "01000000", "00111110", 
"00111100", "00111010", "00111000", "00110110", "00110011", "00110001", "00101111", "00101100", "00101010", "00100111", "00100101", "00100010", "00011111", "00011101", "00011010", "00010111", "00010100", "00010010", "00001111", "00001100", 
"00001001", "00000110", "00000011", "00000000", "11111101", "11111010", "11110111", "11110101", "11110010", "11101111", "11101100", "11101001", "11100111", "11100100", "11100001", "11011111", "11011100", "11011001", "11010111", "11010101", 
"11010010", "11010000", "11001110", "11001011", "11001001", "11000111", "11000101", "11000011", "11000001", "10111111", "10111110", "10111100", "10111010", "10111000", "10110111", "10110101", "10110100", "10110010", "10110001", "10110000", 
"10101110", "10101101", "10101100", "10101011", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", 
"01001110", "01001101", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", 
"00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111011", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110101", "00110101", 
"00110100", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", "00110001", "00110001", "00110001", "00110000", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101110", "00101101", "00101101", 
"00101101", "00101100", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "00101010", "00101010", "00101010", "11010111", "11010110", "11010110", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", 
"11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", "11010010", "11010001", "11010001", "11010000", "11010000", "11010000", "11001111", "11001111", "11001111", "11001110", "11001110", "11001101", "11001101", 
"11001100", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000101", "11000100", "11000011", "11000011", 
"11000010", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", 
"10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010101", 
"01010100", "01010011", "01010010", "01010000", "01001111", "01001110", "01001100", "01001011", "01001001", "01001000", "01000110", "01000100", "01000010", "01000001", "00111111", "00111101", "00111011", "00111001", "00110111", "00110101", 
"00110010", "00110000", "00101110", "00101011", "00101001", "00100111", "00100100", "00100001", "00011111", "00011100", "00011001", "00010111", "00010100", "00010001", "00001110", "00001011", "00001001", "00000110", "00000011", "00000000", 
"11111101", "11111010", "11111000", "11110101", "11110010", "11101111", "11101100", "11101010", "11100111", "11100100", "11100010", "11011111", "11011101", "11011010", "11011000", "11010101", "11010011", "11010001", "11001111", "11001100", 
"11001010", "11001000", "11000110", "11000100", "11000010", "11000000", "10111111", "10111101", "10111011", "10111010", "10111000", "10110110", "10110101", "10110011", "10110010", "10110001", "10101111", "10101110", "10101101", "10101100", 
"10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001101", "01001100", 
"01001011", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", 
"00111110", "00111101", "00111101", "00111100", "00111011", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110101", "00110101", "00110101", "00110100", 
"00110100", "00110011", "00110011", "00110010", "00110010", "00110010", "00110001", "00110001", "00110000", "00110000", "00110000", "00101111", "00101111", "00101111", "00101110", "00101110", "00101110", "00101101", "00101101", "00101101", 
"00101100", "00101100", "00101100", "00101011", "00101011", "00101011", "00101010", "11010110", "11010110", "11010101", "11010101", "11010101", "11010100", "11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", 
"11010010", "11010001", "11010001", "11010001", "11010000", "11010000", "11010000", "11001111", "11001111", "11001110", "11001110", "11001110", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001011", "11001010", 
"11001010", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000101", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "10111111", 
"10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", 
"10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010100", "01010011", "01010010", "01010001", "01001111", 
"01001110", "01001101", "01001011", "01001010", "01001000", "01000110", "01000101", "01000011", "01000001", "01000000", "00111110", "00111100", "00111010", "00111000", "00110110", "00110100", "00110001", "00101111", "00101101", "00101011", 
"00101000", "00100110", "00100011", "00100001", "00011110", "00011100", "00011001", "00010110", "00010100", "00010001", "00001110", "00001011", "00001000", "00000110", "00000011", "00000000", "11111101", "11111010", "11111000", "11110101", 
"11110010", "11110000", "11101101", "11101010", "11101000", "11100101", "11100010", "11100000", "11011101", "11011011", "11011001", "11010110", "11010100", "11010010", "11010000", "11001101", "11001011", "11001001", "11000111", "11000101", 
"11000011", "11000010", "11000000", "10111110", "10111100", "10111011", "10111001", "10110111", "10110110", "10110101", "10110011", "10110010", "10110000", "10101111", "10101110", "10101101", "10101011", "10101010", "10101001", "10101000", 
"10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", 
"01001001", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", "00111110", "00111101", 
"00111100", "00111100", "00111011", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", 
"00110011", "00110011", "00110010", "00110010", "00110001", "00110001", "00110001", "00110000", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101110", "00101101", "00101101", "00101101", "00101100", "00101100", 
"00101100", "00101100", "00101011", "11010101", "11010101", "11010100", "11010100", "11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", "11010010", "11010001", "11010001", "11010000", "11010000", "11010000", 
"11001111", "11001111", "11001111", "11001110", "11001110", "11001101", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11000111", 
"11000111", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", 
"10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", 
"10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010011", "01010010", "01010001", "01010000", "01001110", "01001101", "01001011", "01001010", "01001001", 
"01000111", "01000101", "01000100", "01000010", "01000000", "00111110", "00111101", "00111011", "00111001", "00110111", "00110101", "00110011", "00110000", "00101110", "00101100", "00101010", "00100111", "00100101", "00100011", "00100000", 
"00011110", "00011011", "00011000", "00010110", "00010011", "00010000", "00001110", "00001011", "00001000", "00000110", "00000011", "00000000", "11111101", "11111011", "11111000", "11110101", "11110011", "11110000", "11101101", "11101011", 
"11101000", "11100110", "11100011", "11100001", "11011110", "11011100", "11011001", "11010111", "11010101", "11010011", "11010000", "11001110", "11001100", "11001010", "11001000", "11000110", "11000100", "11000011", "11000001", "10111111", 
"10111101", "10111100", "10111010", "10111001", "10110111", "10110110", "10110100", "10110011", "10110001", "10110000", "10101111", "10101110", "10101101", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", 
"01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001110", "01001101", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", 
"01000111", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", "00111101", "00111101", "00111100", "00111100", 
"00111011", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110011", 
"00110010", "00110010", "00110010", "00110001", "00110001", "00110000", "00110000", "00110000", "00101111", "00101111", "00101111", "00101110", "00101110", "00101110", "00101101", "00101101", "00101101", "00101100", "00101100", "11010100", 
"11010100", "11010100", "11010011", "11010011", "11010011", "11010010", "11010010", "11010010", "11010001", "11010001", "11010001", "11010000", "11010000", "11010000", "11001111", "11001111", "11001110", "11001110", "11001110", "11001101", 
"11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000101", "11000100", 
"11000100", "11000011", "11000011", "11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", 
"10110111", "10110110", "10110110", "10110101", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", 
"10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010011", "01010010", "01010001", "01010000", "01001111", "01001101", "01001100", "01001010", "01001001", "01000111", "01000110", "01000100", "01000011", "01000001", 
"00111111", "00111101", "00111100", "00111010", "00111000", "00110110", "00110100", "00110010", "00110000", "00101101", "00101011", "00101001", "00100111", "00100100", "00100010", "00011111", "00011101", "00011010", "00011000", "00010101", 
"00010011", "00010000", "00001101", "00001011", "00001000", "00000101", "00000011", "00000000", "11111101", "11111011", "11111000", "11110101", "11110011", "11110000", "11101110", "11101011", "11101001", "11100110", "11100100", "11100001", 
"11011111", "11011100", "11011010", "11011000", "11010110", "11010011", "11010001", "11001111", "11001101", "11001011", "11001001", "11000111", "11000101", "11000100", "11000010", "11000000", "10111110", "10111101", "10111011", "10111010", 
"10111000", "10110111", "10110101", "10110100", "10110010", "10110001", "10110000", "10101111", "10101110", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", 
"01010101", "01010100", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000110", 
"01000110", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000001", "01000001", "01000000", "01000000", "00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", 
"00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00110111", "00110111", "00110111", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", 
"00110010", "00110001", "00110001", "00110001", "00110000", "00110000", "00110000", "00101111", "00101111", "00101110", "00101110", "00101110", "00101110", "00101101", "00101101", "11010011", "11010011", "11010011", "11010010", "11010010", 
"11010010", "11010010", "11010001", "11010001", "11010000", "11010000", "11010000", "11001111", "11001111", "11001111", "11001110", "11001110", "11001110", "11001101", "11001101", "11001100", "11001100", "11001100", "11001011", "11001011", 
"11001010", "11001010", "11001001", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", 
"11000000", "11000000", "10111111", "10111111", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", 
"10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", 
"01010101", "01010100", "01010010", "01010001", "01010000", "01001111", "01001110", "01001100", "01001011", "01001001", "01001000", "01000110", "01000101", "01000011", "01000010", "01000000", "00111110", "00111100", "00111011", "00111001", 
"00110111", "00110101", "00110011", "00110001", "00101111", "00101101", "00101010", "00101000", "00100110", "00100100", "00100001", "00011111", "00011100", "00011010", "00010111", "00010101", "00010010", "00010000", "00001101", "00001011", 
"00001000", "00000101", "00000011", "00000000", "11111101", "11111011", "11111000", "11110110", "11110011", "11110001", "11101110", "11101100", "11101001", "11100111", "11100100", "11100010", "11011111", "11011101", "11011011", "11011001", 
"11010110", "11010100", "11010010", "11010000", "11001110", "11001100", "11001010", "11001000", "11000110", "11000100", "11000011", "11000001", "10111111", "10111110", "10111100", "10111011", "10111001", "10111000", "10110110", "10110101", 
"10110011", "10110010", "10110001", "10110000", "10101111", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010100", 
"01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01000111", "01000111", "01000110", "01000101", "01000101", 
"01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111010", "00111010", 
"00111001", "00111001", "00111000", "00111000", "00110111", "00110111", "00110111", "00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110100", "00110011", "00110011", "00110011", "00110010", "00110010", "00110001", 
"00110001", "00110001", "00110000", "00110000", "00110000", "00101111", "00101111", "00101111", "00101110", "00101110", "00101110", "11010011", "11010010", "11010010", "11010010", "11010001", "11010001", "11010001", "11010000", "11010000", 
"11010000", "11001111", "11001111", "11001111", "11001110", "11001110", "11001101", "11001101", "11001101", "11001100", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001001", "11001001", "11001001", "11001000", 
"11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "10111111", "10111111", "10111110", "10111110", 
"10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110001", "10110000", "10110000", 
"10101111", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010001", "01010000", 
"01001111", "01001110", "01001101", "01001011", "01001010", "01001000", "01000111", "01000101", "01000100", "01000010", "01000001", "00111111", "00111101", "00111100", "00111010", "00111000", "00110110", "00110100", "00110010", "00110000", 
"00101110", "00101100", "00101010", "00100111", "00100101", "00100011", "00100001", "00011110", "00011100", "00011001", "00010111", "00010100", "00010010", "00001111", "00001101", "00001010", "00001000", "00000101", "00000011", "00000000", 
"11111101", "11111011", "11111000", "11110110", "11110011", "11110001", "11101110", "11101100", "11101010", "11100111", "11100101", "11100010", "11100000", "11011110", "11011100", "11011001", "11010111", "11010101", "11010011", "11010001", 
"11001111", "11001101", "11001011", "11001001", "11000111", "11000101", "11000100", "11000010", "11000000", "10111111", "10111101", "10111100", "10111010", "10111001", "10110111", "10110110", "10110100", "10110011", "10110010", "10110001", 
"10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010010", "01010001", 
"01010001", "01010000", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000011", 
"01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111010", "00111010", "00111001", "00111001", 
"00111000", "00111000", "00110111", "00110111", "00110111", "00110110", "00110110", "00110101", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110011", "00110010", "00110010", "00110010", "00110001", "00110001", 
"00110001", "00110000", "00110000", "00101111", "00101111", "00101111", "00101111", "11010010", "11010001", "11010001", "11010001", "11010001", "11010000", "11010000", "11001111", "11001111", "11001111", "11001110", "11001110", "11001110", 
"11001101", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001011", "11001010", "11001010", "11001001", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", 
"11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", 
"10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", "10101011", 
"10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01001111", "01001110", "01001101", "01001100", "01001010", 
"01001001", "01000111", "01000110", "01000100", "01000011", "01000001", "01000000", "00111110", "00111100", "00111011", "00111001", "00110111", "00110101", "00110011", "00110001", "00101111", "00101101", "00101011", "00101001", "00100111", 
"00100100", "00100010", "00100000", "00011110", "00011011", "00011001", "00010110", "00010100", "00010010", "00001111", "00001101", "00001010", "00001000", "00000101", "00000011", "00000000", "11111110", "11111011", "11111001", "11110110", 
"11110100", "11110001", "11101111", "11101100", "11101010", "11101000", "11100101", "11100011", "11100001", "11011110", "11011100", "11011010", "11011000", "11010110", "11010100", "11010010", "11010000", "11001110", "11001100", "11001010", 
"11001000", "11000110", "11000101", "11000011", "11000001", "11000000", "10111110", "10111101", "10111011", "10111010", "10111000", "10110111", "10110101", "10110100", "10110011", "10110010", "10110000", "10101111", "10101110", "10101101", 
"10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", 
"01001110", "01001110", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000010", 
"01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", 
"00110111", "00110111", "00110111", "00110110", "00110110", "00110101", "00110101", "00110101", "00110100", "00110100", "00110011", "00110011", "00110011", "00110010", "00110010", "00110010", "00110001", "00110001", "00110001", "00110000", 
"00110000", "00110000", "00101111", "11010001", "11010001", "11010000", "11010000", "11010000", "11001111", "11001111", "11001111", "11001110", "11001110", "11001110", "11001101", "11001101", "11001101", "11001100", "11001100", "11001011", 
"11001011", "11001011", "11001010", "11001010", "11001001", "11001001", "11001001", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", 
"11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", 
"10110110", "10110101", "10110101", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10100111", 
"10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001110", "01001101", "01001100", "01001011", "01001001", "01001000", "01000110", "01000101", "01000011", 
"01000010", "01000000", "00111111", "00111101", "00111011", "00111010", "00111000", "00110110", "00110100", "00110010", "00110000", "00101110", "00101100", "00101010", "00101000", "00100110", "00100100", "00100010", "00011111", "00011101", 
"00011011", "00011000", "00010110", "00010100", "00010001", "00001111", "00001100", "00001010", "00000111", "00000101", "00000010", "00000000", "11111110", "11111011", "11111001", "11110110", "11110100", "11110001", "11101111", "11101101", 
"11101010", "11101000", "11100110", "11100011", "11100001", "11011111", "11011101", "11011011", "11011001", "11010110", "11010100", "11010010", "11010000", "11001111", "11001101", "11001011", "11001001", "11000111", "11000101", "11000100", 
"11000010", "11000001", "10111111", "10111101", "10111100", "10111010", "10111001", "10111000", "10110110", "10110101", "10110100", "10110011", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", 
"10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", 
"01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", 
"01000000", "01000000", "00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111100", "00111011", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00111000", "00110111", 
"00110111", "00110110", "00110110", "00110101", "00110101", "00110101", "00110100", "00110100", "00110100", "00110011", "00110011", "00110010", "00110010", "00110010", "00110001", "00110001", "00110001", "00110000", "00110000", "11010000", 
"11010000", "11010000", "11001111", "11001111", "11001111", "11001110", "11001110", "11001110", "11001101", "11001101", "11001100", "11001100", "11001100", "11001011", "11001011", "11001011", "11001010", "11001010", "11001001", "11001001", 
"11001000", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000000", "11000000", "10111111", 
"10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", 
"10110010", "10110001", "10110001", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", 
"01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001101", "01001100", "01001011", "01001010", "01001000", "01000111", "01000110", "01000100", "01000011", "01000001", "00111111", "00111110", "00111100", 
"00111011", "00111001", "00110111", "00110101", "00110011", "00110001", "00110000", "00101110", "00101100", "00101010", "00100111", "00100101", "00100011", "00100001", "00011111", "00011101", "00011010", "00011000", "00010110", "00010011", 
"00010001", "00001111", "00001100", "00001010", "00000111", "00000101", "00000010", "00000000", "11111110", "11111011", "11111001", "11110110", "11110100", "11110010", "11101111", "11101101", "11101011", "11101000", "11100110", "11100100", 
"11100010", "11100000", "11011101", "11011011", "11011001", "11010111", "11010101", "11010011", "11010001", "11001111", "11001101", "11001100", "11001010", "11001000", "11000110", "11000101", "11000011", "11000001", "11000000", "10111110", 
"10111101", "10111011", "10111010", "10111001", "10110111", "10110110", "10110101", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", 
"10100110", "01011001", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", 
"01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", 
"00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00111000", "00110111", "00110111", "00110110", 
"00110110", "00110110", "00110101", "00110101", "00110100", "00110100", "00110100", "00110011", "00110011", "00110011", "00110010", "00110010", "00110010", "00110001", "00110001", "11001111", "11001111", "11001111", "11001110", "11001110", 
"11001110", "11001101", "11001101", "11001101", "11001100", "11001100", "11001100", "11001011", "11001011", "11001010", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11001000", "11000111", "11000111", "11000110", 
"11000110", "11000101", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", 
"10111100", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110000", "10110000", "10101111", 
"10101110", "10101101", "10101101", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", 
"01010000", "01001111", "01001110", "01001101", "01001011", "01001010", "01001001", "01000111", "01000110", "01000101", "01000011", "01000010", "01000000", "00111111", "00111101", "00111011", "00111010", "00111000", "00110110", "00110100", 
"00110011", "00110001", "00101111", "00101101", "00101011", "00101001", "00100111", "00100101", "00100011", "00100000", "00011110", "00011100", "00011010", "00011000", "00010101", "00010011", "00010001", "00001110", "00001100", "00001010", 
"00000111", "00000101", "00000010", "00000000", "11111110", "11111011", "11111001", "11110111", "11110100", "11110010", "11110000", "11101101", "11101011", "11101001", "11100111", "11100100", "11100010", "11100000", "11011110", "11011100", 
"11011010", "11011000", "11010110", "11010100", "11010010", "11010000", "11001110", "11001100", "11001011", "11001001", "11000111", "11000110", "11000100", "11000010", "11000001", "10111111", "10111110", "10111100", "10111011", "10111010", 
"10111000", "10110111", "10110110", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", 
"01010111", "01010111", "01010110", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", 
"01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", 
"00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111011", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110110", 
"00110101", "00110101", "00110100", "00110100", "00110100", "00110011", "00110011", "00110011", "00110010", "00110010", "00110010", "11001111", "11001110", "11001110", "11001110", "11001101", "11001101", "11001101", "11001100", "11001100", 
"11001100", "11001011", "11001011", "11001010", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000101", "11000101", "11000101", "11000100", "11000100", 
"11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", 
"10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", 
"10101010", "10101001", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", 
"01001010", "01001001", "01001000", "01000110", "01000101", "01000100", "01000010", "01000001", "00111111", "00111110", "00111100", "00111010", "00111001", "00110111", "00110101", "00110100", "00110010", "00110000", "00101110", "00101100", 
"00101010", "00101000", "00100110", "00100100", "00100010", "00100000", "00011110", "00011100", "00011001", "00010111", "00010101", "00010011", "00010000", "00001110", "00001100", "00001001", "00000111", "00000101", "00000010", "00000000", 
"11111110", "11111011", "11111001", "11110111", "11110101", "11110010", "11110000", "11101110", "11101011", "11101001", "11100111", "11100101", "11100011", "11100001", "11011111", "11011101", "11011010", "11011000", "11010111", "11010101", 
"11010011", "11010001", "11001111", "11001101", "11001011", "11001010", "11001000", "11000110", "11000101", "11000011", "11000010", "11000000", "10111111", "10111101", "10111100", "10111010", "10111001", "10111000", "10110111", "10110101", 
"10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010111", "01010110", 
"01010101", "01010100", "01010100", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", 
"01000111", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111101", 
"00111101", "00111100", "00111100", "00111011", "00111011", "00111010", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110110", "00110101", "00110101", 
"00110101", "00110100", "00110100", "00110011", "00110011", "00110011", "00110010", "11001110", "11001110", "11001101", "11001101", "11001101", "11001100", "11001100", "11001011", "11001011", "11001011", "11001010", "11001010", "11001010", 
"11001001", "11001001", "11001000", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", 
"11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110110", 
"10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", 
"10100110", "01011001", "01011000", "01010111", "01010110", "01010101", "01010100", "01010100", "01010011", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001001", "01001000", "01000111", "01000110", 
"01000100", "01000011", "01000001", "01000000", "00111110", "00111101", "00111011", "00111010", "00111000", "00110110", "00110101", "00110011", "00110001", "00101111", "00101101", "00101011", "00101001", "00101000", "00100110", "00100011", 
"00100001", "00011111", "00011101", "00011011", "00011001", "00010111", "00010101", "00010010", "00010000", "00001110", "00001011", "00001001", "00000111", "00000101", "00000010", "00000000", "11111110", "11111011", "11111001", "11110111", 
"11110101", "11110010", "11110000", "11101110", "11101100", "11101010", "11101000", "11100101", "11100011", "11100001", "11011111", "11011101", "11011011", "11011001", "11010111", "11010101", "11010011", "11010010", "11010000", "11001110", 
"11001100", "11001011", "11001001", "11000111", "11000110", "11000100", "11000010", "11000001", "11000000", "10111110", "10111101", "10111011", "10111010", "10111001", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", 
"10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010100", "01010100", 
"01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000110", 
"01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111100", 
"00111100", "00111011", "00111011", "00111010", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110110", "00110101", "00110101", "00110101", "00110100", 
"00110100", "00110100", "00110011", "11001101", "11001101", "11001100", "11001100", "11001100", "11001011", "11001011", "11001011", "11001010", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11001000", "11000111", 
"11000111", "11000110", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", 
"10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", 
"10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", 
"01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01000111", "01000110", "01000101", "01000011", "01000010", "01000000", "00111111", 
"00111110", "00111100", "00111010", "00111001", "00110111", "00110101", "00110100", "00110010", "00110000", "00101110", "00101101", "00101011", "00101001", "00100111", "00100101", "00100011", "00100001", "00011111", "00011101", "00011011", 
"00011000", "00010110", "00010100", "00010010", "00010000", "00001110", "00001011", "00001001", "00000111", "00000101", "00000010", "00000000", "11111110", "11111100", "11111001", "11110111", "11110101", "11110011", "11110001", "11101110", 
"11101100", "11101010", "11101000", "11100110", "11100100", "11100010", "11100000", "11011110", "11011100", "11011010", "11011000", "11010110", "11010100", "11010010", "11010000", "11001111", "11001101", "11001011", "11001010", "11001000", 
"11000110", "11000101", "11000011", "11000010", "11000000", "10111111", "10111110", "10111100", "10111011", "10111010", "10111000", "10110111", "10110110", "10110101", "10110100", "10110010", "10110001", "10110000", "10101111", "10101110", 
"10101101", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", 
"01010001", "01010000", "01010000", "01001111", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", 
"01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111101", "00111100", "00111100", "00111011", 
"00111011", "00111010", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00111000", "00110111", "00110111", "00110110", "00110110", "00110110", "00110101", "00110101", "00110101", "00110100", "00110100", "11001100", 
"11001100", "11001100", "11001011", "11001011", "11001011", "11001010", "11001010", "11001010", "11001001", "11001001", "11001000", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000110", "11000101", "11000101", 
"11000100", "11000100", "11000011", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", 
"10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", 
"10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010011", "01010010", 
"01010001", "01010000", "01001111", "01001110", "01001100", "01001011", "01001010", "01001001", "01001000", "01000110", "01000101", "01000100", "01000010", "01000001", "01000000", "00111110", "00111101", "00111011", "00111010", "00111000", 
"00110110", "00110101", "00110011", "00110001", "00110000", "00101110", "00101100", "00101010", "00101000", "00100110", "00100100", "00100010", "00100000", "00011110", "00011100", "00011010", "00011000", "00010110", "00010100", "00010010", 
"00001111", "00001101", "00001011", "00001001", "00000111", "00000100", "00000010", "00000000", "11111110", "11111100", "11111001", "11110111", "11110101", "11110011", "11110001", "11101111", "11101101", "11101010", "11101000", "11100110", 
"11100100", "11100010", "11100000", "11011110", "11011100", "11011010", "11011000", "11010111", "11010101", "11010011", "11010001", "11001111", "11001110", "11001100", "11001010", "11001001", "11000111", "11000110", "11000100", "11000011", 
"11000001", "11000000", "10111110", "10111101", "10111100", "10111010", "10111001", "10111000", "10110111", "10110110", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", 
"10101010", "10101001", "10101001", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", 
"01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", 
"01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111010", 
"00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00111000", "00110111", "00110111", "00110111", "00110110", "00110110", "00110101", "00110101", "00110101", "11001100", "11001011", "11001011", "11001011", "11001010", 
"11001010", "11001001", "11001001", "11001001", "11001000", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000011", "11000010", 
"11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", 
"10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101011", "10101011", 
"10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", 
"01001100", "01001010", "01001001", "01001000", "01000111", "01000110", "01000100", "01000011", "01000010", "01000000", "00111111", "00111101", "00111100", "00111010", "00111001", "00110111", "00110110", "00110100", "00110010", "00110001", 
"00101111", "00101101", "00101011", "00101001", "00101000", "00100110", "00100100", "00100010", "00100000", "00011110", "00011100", "00011010", "00011000", "00010110", "00010011", "00010001", "00001111", "00001101", "00001011", "00001001", 
"00000111", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11110111", "11110101", "11110011", "11110001", "11101111", "11101101", "11101011", "11101001", "11100111", "11100101", "11100011", "11100001", "11011111", 
"11011101", "11011011", "11011001", "11010111", "11010101", "11010100", "11010010", "11010000", "11001110", "11001101", "11001011", "11001010", "11001000", "11000110", "11000101", "11000011", "11000010", "11000001", "10111111", "10111110", 
"10111101", "10111011", "10111010", "10111001", "10111000", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101001", 
"10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", 
"01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000010", 
"01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111100", "00111011", "00111011", "00111010", "00111010", "00111010", 
"00111001", "00111001", "00111000", "00111000", "00111000", "00110111", "00110111", "00110111", "00110110", "00110110", "00110110", "11001011", "11001010", "11001010", "11001010", "11001001", "11001001", "11001001", "11001000", "11001000", 
"11001000", "11000111", "11000111", "11000110", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "10111111", 
"10111111", "10111110", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110101", 
"10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101000", "10101000", "10100111", 
"10100110", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001000", "01000111", 
"01000110", "01000101", "01000011", "01000010", "01000001", "00111111", "00111110", "00111101", "00111011", "00111010", "00111000", "00110110", "00110101", "00110011", "00110010", "00110000", "00101110", "00101100", "00101011", "00101001", 
"00100111", "00100101", "00100011", "00100001", "00011111", "00011101", "00011011", "00011001", "00010111", "00010101", "00010011", "00010001", "00001111", "00001101", "00001011", "00001001", "00000110", "00000100", "00000010", "00000000", 
"11111110", "11111100", "11111010", "11111000", "11110101", "11110011", "11110001", "11101111", "11101101", "11101011", "11101001", "11100111", "11100101", "11100011", "11100001", "11011111", "11011101", "11011100", "11011010", "11011000", 
"11010110", "11010100", "11010011", "11010001", "11001111", "11001110", "11001100", "11001010", "11001001", "11000111", "11000110", "11000100", "11000011", "11000001", "11000000", "10111111", "10111101", "10111100", "10111011", "10111010", 
"10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100110", 
"01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", 
"01001100", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", 
"01000001", "01000000", "01000000", "00111111", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111100", "00111011", "00111011", "00111010", "00111010", "00111010", "00111001", "00111001", 
"00111000", "00111000", "00111000", "00110111", "00110111", "00110111", "00110110", "11001010", "11001010", "11001001", "11001001", "11001001", "11001000", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000110", 
"11000101", "11000101", "11000100", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", 
"10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110001", 
"10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01010111", "01010111", 
"01010110", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000110", "01000101", "01000100", "01000011", "01000001", 
"01000000", "00111111", "00111101", "00111100", "00111010", "00111001", "00110111", "00110110", "00110100", "00110010", "00110001", "00101111", "00101101", "00101100", "00101010", "00101000", "00100110", "00100100", "00100011", "00100001", 
"00011111", "00011101", "00011011", "00011001", "00010111", "00010101", "00010011", "00010001", "00001111", "00001101", "00001011", "00001000", "00000110", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11111000", 
"11110110", "11110100", "11110010", "11101111", "11101101", "11101011", "11101001", "11100111", "11100110", "11100100", "11100010", "11100000", "11011110", "11011100", "11011010", "11011000", "11010111", "11010101", "11010011", "11010010", 
"11010000", "11001110", "11001101", "11001011", "11001001", "11001000", "11000110", "11000101", "11000100", "11000010", "11000001", "10111111", "10111110", "10111101", "10111100", "10111010", "10111001", "10111000", "10110111", "10110110", 
"10110101", "10110100", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", 
"01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001011", 
"01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", 
"01000000", "00111111", "00111111", "00111110", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111100", "00111011", "00111011", "00111010", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", 
"00111000", "00110111", "00110111", "11001001", "11001001", "11001001", "11001000", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000110", "11000101", "11000101", "11000100", "11000100", "11000100", "11000011", 
"11000011", "11000010", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", 
"10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", 
"10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010010", 
"01010001", "01010001", "01010000", "01001111", "01001110", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000100", "01000011", "01000010", "01000001", "00111111", "00111110", "00111100", "00111011", 
"00111010", "00111000", "00110111", "00110101", "00110011", "00110010", "00110000", "00101110", "00101101", "00101011", "00101001", "00101000", "00100110", "00100100", "00100010", "00100000", "00011110", "00011100", "00011010", "00011001", 
"00010111", "00010101", "00010011", "00010001", "00001110", "00001100", "00001010", "00001000", "00000110", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11111000", "11110110", "11110100", "11110010", "11110000", 
"11101110", "11101100", "11101010", "11101000", "11100110", "11100100", "11100010", "11100000", "11011110", "11011101", "11011011", "11011001", "11010111", "11010110", "11010100", "11010010", "11010001", "11001111", "11001101", "11001100", 
"11001010", "11001001", "11000111", "11000110", "11000100", "11000011", "11000010", "11000000", "10111111", "10111110", "10111100", "10111011", "10111010", "10111001", "10111000", "10110110", "10110101", "10110100", "10110011", "10110010", 
"10110001", "10110000", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", 
"01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", 
"01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000001", "01000000", "01000000", "00111111", 
"00111111", "00111110", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111011", "00111010", "00111010", "00111010", "00111001", "00111001", "00111000", "00111000", "00111000", "11001001", 
"11001000", "11001000", "11001000", "11000111", "11000111", "11000110", "11000110", "11000110", "11000101", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000010", "11000001", "11000001", 
"11000000", "11000000", "10111111", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110111", 
"10110110", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", 
"10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", 
"01001101", "01001100", "01001011", "01001010", "01001000", "01000111", "01000110", "01000101", "01000100", "01000010", "01000001", "01000000", "00111110", "00111101", "00111100", "00111010", "00111001", "00110111", "00110110", "00110100", 
"00110011", "00110001", "00101111", "00101110", "00101100", "00101010", "00101001", "00100111", "00100101", "00100011", "00100010", "00100000", "00011110", "00011100", "00011010", "00011000", "00010110", "00010100", "00010010", "00010000", 
"00001110", "00001100", "00001010", "00001000", "00000110", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11111000", "11110110", "11110100", "11110010", "11110000", "11101110", "11101100", "11101010", "11101000", 
"11100110", "11100100", "11100011", "11100001", "11011111", "11011101", "11011011", "11011010", "11011000", "11010110", "11010100", "11010011", "11010001", "11010000", "11001110", "11001100", "11001011", "11001001", "11001000", "11000110", 
"11000101", "11000100", "11000010", "11000001", "11000000", "10111110", "10111101", "10111100", "10111011", "10111010", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", 
"10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", 
"01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", 
"01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "01000000", "00111111", "00111111", "00111110", 
"00111110", "00111101", "00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111011", "00111010", "00111010", "00111010", "00111001", "00111001", "00111000", "11001000", "11001000", "11000111", "11000111", "11000110", 
"11000110", "11000110", "11000101", "11000101", "11000101", "11000100", "11000100", "11000011", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "11000000", "10111111", "10111111", "10111110", 
"10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", 
"10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", 
"10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", 
"01001000", "01000110", "01000101", "01000100", "01000011", "01000010", "01000000", "00111111", "00111110", "00111100", "00111011", "00111010", "00111000", "00110111", "00110101", "00110100", "00110010", "00110000", "00101111", "00101101", 
"00101100", "00101010", "00101000", "00100110", "00100101", "00100011", "00100001", "00011111", "00011101", "00011100", "00011010", "00011000", "00010110", "00010100", "00010010", "00010000", "00001110", "00001100", "00001010", "00001000", 
"00000110", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11111000", "11110110", "11110100", "11110010", "11110000", "11101110", "11101100", "11101010", "11101001", "11100111", "11100101", "11100011", "11100001", 
"11011111", "11011110", "11011100", "11011010", "11011000", "11010111", "11010101", "11010011", "11010010", "11010000", "11001111", "11001101", "11001100", "11001010", "11001001", "11000111", "11000110", "11000100", "11000011", "11000010", 
"11000000", "10111111", "10111110", "10111101", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", 
"10101100", "10101011", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", 
"01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", 
"01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111111", "00111110", "00111110", "00111101", 
"00111101", "00111101", "00111100", "00111100", "00111011", "00111011", "00111011", "00111010", "00111010", "00111010", "00111001", "11000111", "11000111", "11000110", "11000110", "11000110", "11000101", "11000101", "11000101", "11000100", 
"11000100", "11000011", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111101", "10111100", "10111100", 
"10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110001", 
"10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", 
"01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000011", 
"01000010", "01000001", "01000000", "00111110", "00111101", "00111100", "00111010", "00111001", "00110111", "00110110", "00110100", "00110011", "00110001", "00110000", "00101110", "00101101", "00101011", "00101001", "00101000", "00100110", 
"00100100", "00100010", "00100001", "00011111", "00011101", "00011011", "00011001", "00010111", "00010110", "00010100", "00010010", "00010000", "00001110", "00001100", "00001010", "00001000", "00000110", "00000100", "00000010", "00000000", 
"11111110", "11111100", "11111010", "11111000", "11110110", "11110100", "11110010", "11110000", "11101111", "11101101", "11101011", "11101001", "11100111", "11100101", "11100011", "11100010", "11100000", "11011110", "11011100", "11011011", 
"11011001", "11010111", "11010110", "11010100", "11010010", "11010001", "11001111", "11001110", "11001100", "11001011", "11001001", "11001000", "11000111", "11000101", "11000100", "11000010", "11000001", "11000000", "10111111", "10111101", 
"10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101011", "10101010", 
"10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", 
"01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", 
"01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111110", "00111101", "00111101", "00111100", 
"00111100", "00111100", "00111011", "00111011", "00111011", "00111010", "00111010", "11000110", "11000110", "11000110", "11000101", "11000101", "11000101", "11000100", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", 
"11000010", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", 
"10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", 
"10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", 
"01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000001", "01000000", "00111111", "00111110", 
"00111100", "00111011", "00111001", "00111000", "00110111", "00110101", "00110100", "00110010", "00110001", "00101111", "00101110", "00101100", "00101010", "00101001", "00100111", "00100101", "00100100", "00100010", "00100000", "00011110", 
"00011101", "00011011", "00011001", "00010111", "00010101", "00010011", "00010001", "00010000", "00001110", "00001100", "00001010", "00001000", "00000110", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11111000", 
"11110110", "11110101", "11110011", "11110001", "11101111", "11101101", "11101011", "11101001", "11100111", "11100110", "11100100", "11100010", "11100000", "11011111", "11011101", "11011011", "11011001", "11011000", "11010110", "11010101", 
"11010011", "11010001", "11010000", "11001110", "11001101", "11001011", "11001010", "11001001", "11000111", "11000110", "11000101", "11000011", "11000010", "11000001", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", 
"10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101000", "10101000", 
"10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001110", 
"01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000101", "01000100", 
"01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111100", 
"00111011", "00111011", "00111011", "11000110", "11000101", "11000101", "11000101", "11000100", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "11000000", 
"10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", 
"10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", 
"10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", 
"01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "00111111", "00111110", "00111101", "00111011", "00111010", "00111001", "00110111", 
"00110110", "00110101", "00110011", "00110010", "00110000", "00101111", "00101101", "00101011", "00101010", "00101000", "00100111", "00100101", "00100011", "00100001", "00100000", "00011110", "00011100", "00011010", "00011001", "00010111", 
"00010101", "00010011", "00010001", "00001111", "00001101", "00001011", "00001010", "00001000", "00000110", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11111000", "11110111", "11110101", "11110011", "11110001", 
"11101111", "11101101", "11101011", "11101010", "11101000", "11100110", "11100100", "11100011", "11100001", "11011111", "11011101", "11011100", "11011010", "11011000", "11010111", "11010101", "11010100", "11010010", "11010001", "11001111", 
"11001110", "11001100", "11001011", "11001001", "11001000", "11000111", "11000101", "11000100", "11000011", "11000001", "11000000", "10111111", "10111110", "10111101", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", 
"10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", 
"01011000", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", 
"01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", 
"01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "01000000", "00111111", "00111111", "00111110", "00111110", "00111110", "00111101", "00111101", "00111100", "00111100", "00111100", "00111011", "11000101", 
"11000101", "11000100", "11000100", "11000100", "11000011", "11000011", "11000010", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", 
"10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", 
"10110011", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", 
"10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", 
"01001001", "01001000", "01000111", "01000110", "01000101", "01000011", "01000010", "01000001", "01000000", "00111111", "00111101", "00111100", "00111011", "00111001", "00111000", "00110111", "00110101", "00110100", "00110010", "00110001", 
"00101111", "00101110", "00101100", "00101011", "00101001", "00101000", "00100110", "00100100", "00100011", "00100001", "00011111", "00011101", "00011100", "00011010", "00011000", "00010110", "00010101", "00010011", "00010001", "00001111", 
"00001101", "00001011", "00001001", "00001000", "00000110", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11111001", "11110111", "11110101", "11110011", "11110001", "11101111", "11101110", "11101100", "11101010", 
"11101000", "11100110", "11100101", "11100011", "11100001", "11100000", "11011110", "11011100", "11011011", "11011001", "11010111", "11010110", "11010100", "11010011", "11010001", "11010000", "11001110", "11001101", "11001011", "11001010", 
"11001001", "11000111", "11000110", "11000101", "11000011", "11000010", "11000001", "11000000", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", 
"10110010", "10110001", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", 
"01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", 
"01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", 
"01000001", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111101", "00111100", "00111100", "11000100", "11000100", "11000100", "11000011", "11000011", 
"11000011", "11000010", "11000010", "11000001", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", 
"10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", 
"10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", 
"01010110", "01010110", "01010101", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", 
"01000100", "01000011", "01000010", "01000000", "00111111", "00111110", "00111101", "00111011", "00111010", "00111001", "00110111", "00110110", "00110101", "00110011", "00110010", "00110000", "00101111", "00101101", "00101100", "00101010", 
"00101001", "00100111", "00100101", "00100100", "00100010", "00100000", "00011111", "00011101", "00011011", "00011010", "00011000", "00010110", "00010100", "00010010", "00010001", "00001111", "00001101", "00001011", "00001001", "00000111", 
"00000110", "00000100", "00000010", "00000000", "11111110", "11111100", "11111010", "11111001", "11110111", "11110101", "11110011", "11110001", "11110000", "11101110", "11101100", "11101010", "11101000", "11100111", "11100101", "11100011", 
"11100010", "11100000", "11011110", "11011101", "11011011", "11011001", "11011000", "11010110", "11010101", "11010011", "11010010", "11010000", "11001111", "11001101", "11001100", "11001011", "11001001", "11001000", "11000111", "11000101", 
"11000100", "11000011", "11000010", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", 
"10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", 
"01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", 
"01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", 
"01000001", "01000000", "01000000", "00111111", "00111111", "00111111", "00111110", "00111110", "00111101", "00111101", "00111101", "11000100", "11000011", "11000011", "11000011", "11000010", "11000010", "11000001", "11000001", "11000001", 
"11000000", "11000000", "10111111", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", 
"10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", 
"10101100", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010011", 
"01010011", "01010010", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", 
"00111110", "00111101", "00111100", "00111011", "00111001", "00111000", "00110111", "00110101", "00110100", "00110011", "00110001", "00110000", "00101110", "00101101", "00101011", "00101010", "00101000", "00100111", "00100101", "00100011", 
"00100010", "00100000", "00011110", "00011101", "00011011", "00011001", "00011000", "00010110", "00010100", "00010010", "00010000", "00001111", "00001101", "00001011", "00001001", "00000111", "00000110", "00000100", "00000010", "00000000", 
"11111110", "11111100", "11111011", "11111001", "11110111", "11110101", "11110011", "11110010", "11110000", "11101110", "11101100", "11101011", "11101001", "11100111", "11100101", "11100100", "11100010", "11100000", "11011111", "11011101", 
"11011100", "11011010", "11011000", "11010111", "11010101", "11010100", "11010010", "11010001", "11001111", "11001110", "11001101", "11001011", "11001010", "11001001", "11000111", "11000110", "11000101", "11000011", "11000010", "11000001", 
"11000000", "10111111", "10111110", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10101111", "10101110", "10101101", 
"10101101", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010100", 
"01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", 
"01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", 
"01000000", "00111111", "00111111", "00111110", "00111110", "00111110", "00111101", "11000011", "11000011", "11000010", "11000010", "11000010", "11000001", "11000001", "11000000", "11000000", "11000000", "10111111", "10111111", "10111110", 
"10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", 
"10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", 
"10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010000", "01001111", 
"01001110", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111011", "00111010", 
"00111001", "00110111", "00110110", "00110101", "00110011", "00110010", "00110001", "00101111", "00101110", "00101100", "00101011", "00101001", "00101000", "00100110", "00100100", "00100011", "00100001", "00100000", "00011110", "00011100", 
"00011011", "00011001", "00010111", "00010101", "00010100", "00010010", "00010000", "00001110", "00001101", "00001011", "00001001", "00000111", "00000101", "00000100", "00000010", "00000000", "11111110", "11111100", "11111011", "11111001", 
"11110111", "11110101", "11110100", "11110010", "11110000", "11101110", "11101101", "11101011", "11101001", "11100111", "11100110", "11100100", "11100010", "11100001", "11011111", "11011110", "11011100", "11011010", "11011001", "11010111", 
"11010110", "11010100", "11010011", "11010001", "11010000", "11001111", "11001101", "11001100", "11001010", "11001001", "11001000", "11000111", "11000101", "11000100", "11000011", "11000010", "11000000", "10111111", "10111110", "10111101", 
"10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101101", "10101100", "10101100", "10101011", 
"10101010", "10101010", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", 
"01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", 
"01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", 
"00111111", "00111110", "00111110", "11000010", "11000010", "11000010", "11000001", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", 
"10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", 
"10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", 
"01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111110", "00111101", "00111100", "00111011", "00111001", "00111000", "00110111", "00110110", "00110100", 
"00110011", "00110001", "00110000", "00101111", "00101101", "00101100", "00101010", "00101001", "00100111", "00100110", "00100100", "00100010", "00100001", "00011111", "00011110", "00011100", "00011010", "00011001", "00010111", "00010101", 
"00010011", "00010010", "00010000", "00001110", "00001100", "00001011", "00001001", "00000111", "00000101", "00000100", "00000010", "00000000", "11111110", "11111100", "11111011", "11111001", "11110111", "11110101", "11110100", "11110010", 
"11110000", "11101111", "11101101", "11101011", "11101001", "11101000", "11100110", "11100100", "11100011", "11100001", "11100000", "11011110", "11011100", "11011011", "11011001", "11011000", "11010110", "11010101", "11010011", "11010010", 
"11010001", "11001111", "11001110", "11001100", "11001011", "11001010", "11001000", "11000111", "11000110", "11000101", "11000100", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", 
"10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101001", 
"10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010000", 
"01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", 
"01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000001", "01000000", "01000000", "00111111", "00111111", "00111111", "11000010", 
"11000001", "11000001", "11000001", "11000000", "11000000", "10111111", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111010", 
"10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", 
"10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", 
"01010111", "01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", 
"01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111100", "00111011", "00111010", "00111001", "00111000", "00110110", "00110101", "00110100", "00110010", "00110001", "00101111", "00101110", 
"00101101", "00101011", "00101010", "00101000", "00100111", "00100101", "00100100", "00100010", "00100000", "00011111", "00011101", "00011100", "00011010", "00011000", "00010111", "00010101", "00010011", "00010001", "00010000", "00001110", 
"00001100", "00001011", "00001001", "00000111", "00000101", "00000100", "00000010", "00000000", "11111110", "11111101", "11111011", "11111001", "11110111", "11110110", "11110100", "11110010", "11110000", "11101111", "11101101", "11101011", 
"11101010", "11101000", "11100110", "11100101", "11100011", "11100010", "11100000", "11011110", "11011101", "11011011", "11011010", "11011000", "11010111", "11010101", "11010100", "11010011", "11010001", "11010000", "11001110", "11001101", 
"11001100", "11001010", "11001001", "11001000", "11000111", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", 
"10110101", "10110100", "10110100", "10110011", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", 
"01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", 
"01000101", "01000100", "01000100", "01000100", "01000011", "01000011", "01000010", "01000010", "01000010", "01000001", "01000001", "01000000", "01000000", "01000000", "00111111", "11000001", "11000001", "11000000", "11000000", "11000000", 
"10111111", "10111111", "10111110", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10111000", "10110111", 
"10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", 
"10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010100", "01010100", 
"01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", 
"01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111001", "00111000", "00110111", "00110110", "00110100", "00110011", "00110010", "00110000", "00101111", "00101101", "00101100", "00101011", "00101001", "00101000", 
"00100110", "00100101", "00100011", "00100010", "00100000", "00011110", "00011101", "00011011", "00011010", "00011000", "00010110", "00010101", "00010011", "00010001", "00010000", "00001110", "00001100", "00001010", "00001001", "00000111", 
"00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111001", "11110111", "11110110", "11110100", "11110010", "11110001", "11101111", "11101101", "11101100", "11101010", "11101000", "11100111", "11100101", 
"11100100", "11100010", "11100000", "11011111", "11011101", "11011100", "11011010", "11011001", "11010111", "11010110", "11010100", "11010011", "11010010", "11010000", "11001111", "11001110", "11001100", "11001011", "11001010", "11001000", 
"11000111", "11000110", "11000101", "11000100", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", 
"10110011", "10110010", "10110001", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", 
"01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", 
"01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000110", "01000101", "01000101", "01000100", 
"01000100", "01000011", "01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000001", "01000000", "01000000", "11000000", "11000000", "11000000", "10111111", "10111111", "10111111", "10111110", "10111110", "10111101", 
"10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", 
"10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101010", 
"10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", 
"01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111100", 
"00111011", "00111010", "00111001", "00111000", "00110110", "00110101", "00110100", "00110010", "00110001", "00110000", "00101110", "00101101", "00101100", "00101010", "00101001", "00100111", "00100110", "00100100", "00100011", "00100001", 
"00100000", "00011110", "00011100", "00011011", "00011001", "00011000", "00010110", "00010100", "00010011", "00010001", "00001111", "00001110", "00001100", "00001010", "00001001", "00000111", "00000101", "00000011", "00000010", "00000000", 
"11111110", "11111101", "11111011", "11111001", "11111000", "11110110", "11110100", "11110011", "11110001", "11101111", "11101110", "11101100", "11101010", "11101001", "11100111", "11100110", "11100100", "11100010", "11100001", "11011111", 
"11011110", "11011100", "11011011", "11011001", "11011000", "11010110", "11010101", "11010100", "11010010", "11010001", "11001111", "11001110", "11001101", "11001100", "11001010", "11001001", "11001000", "11000111", "11000101", "11000100", 
"11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110001", 
"10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", 
"01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", 
"01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000101", "01000100", "01000100", "01000011", 
"01000011", "01000011", "01000010", "01000010", "01000001", "01000001", "01000001", "11000000", "10111111", "10111111", "10111111", "10111110", "10111110", "10111101", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", 
"10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", 
"10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001100", 
"01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111001", "00111000", "00110111", 
"00110110", "00110100", "00110011", "00110010", "00110001", "00101111", "00101110", "00101100", "00101011", "00101010", "00101000", "00100111", "00100101", "00100100", "00100010", "00100001", "00011111", "00011110", "00011100", "00011010", 
"00011001", "00010111", "00010110", "00010100", "00010010", "00010001", "00001111", "00001101", "00001100", "00001010", "00001000", "00000111", "00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111001", 
"11111000", "11110110", "11110100", "11110011", "11110001", "11101111", "11101110", "11101100", "11101011", "11101001", "11100111", "11100110", "11100100", "11100011", "11100001", "11100000", "11011110", "11011101", "11011011", "11011010", 
"11011000", "11010111", "11010101", "11010100", "11010011", "11010001", "11010000", "11001111", "11001101", "11001100", "11001011", "11001010", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000001", "11000000", 
"10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101110", 
"10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", 
"01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", 
"01001010", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000100", "01000011", "01000011", "01000010", 
"01000010", "01000010", "01000001", "10111111", "10111111", "10111110", "10111110", "10111110", "10111101", "10111101", "10111100", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111010", "10111001", "10111001", 
"10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", 
"10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", 
"01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", 
"01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110110", "00110101", "00110100", "00110011", "00110001", 
"00110000", "00101111", "00101101", "00101100", "00101011", "00101001", "00101000", "00100110", "00100101", "00100011", "00100010", "00100000", "00011111", "00011101", "00011100", "00011010", "00011001", "00010111", "00010101", "00010100", 
"00010010", "00010001", "00001111", "00001101", "00001100", "00001010", "00001000", "00000111", "00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111001", "11111000", "11110110", "11110101", "11110011", 
"11110001", "11110000", "11101110", "11101100", "11101011", "11101001", "11101000", "11100110", "11100101", "11100011", "11100010", "11100000", "11011111", "11011101", "11011100", "11011010", "11011001", "11010111", "11010110", "11010101", 
"11010011", "11010010", "11010001", "11001111", "11001110", "11001101", "11001011", "11001010", "11001001", "11001000", "11000111", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", 
"10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101101", "10101101", "10101100", 
"10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", 
"01010011", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", 
"01001001", "01001001", "01001000", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "01000011", "01000010", "01000010", "10111111", 
"10111110", "10111110", "10111101", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10111000", "10110111", "10110111", "10110110", 
"10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", 
"10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", 
"01010011", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", 
"01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111001", "00111000", "00110111", "00110110", "00110101", "00110011", "00110010", "00110001", "00101111", "00101110", "00101101", "00101011", 
"00101010", "00101001", "00100111", "00100110", "00100100", "00100011", "00100001", "00100000", "00011110", "00011101", "00011011", "00011010", "00011000", "00010111", "00010101", "00010100", "00010010", "00010000", "00001111", "00001101", 
"00001011", "00001010", "00001000", "00000111", "00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111001", "11111000", "11110110", "11110101", "11110011", "11110001", "11110000", "11101110", "11101101", 
"11101011", "11101010", "11101000", "11100110", "11100101", "11100011", "11100010", "11100000", "11011111", "11011110", "11011100", "11011011", "11011001", "11011000", "11010110", "11010101", "11010100", "11010010", "11010001", "11010000", 
"11001111", "11001101", "11001100", "11001011", "11001010", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", 
"10101001", "10101001", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", 
"01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001001", 
"01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000100", "01000011", "01000011", "01000010", "10111110", "10111110", "10111101", "10111101", "10111100", 
"10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", 
"10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", 
"10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", 
"01010000", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "00111111", "00111110", 
"00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110110", "00110101", "00110100", "00110011", "00110001", "00110000", "00101111", "00101110", "00101100", "00101011", "00101010", "00101000", "00100111", "00100101", 
"00100100", "00100010", "00100001", "00100000", "00011110", "00011101", "00011011", "00011010", "00011000", "00010110", "00010101", "00010011", "00010010", "00010000", "00001111", "00001101", "00001011", "00001010", "00001000", "00000111", 
"00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111010", "11111000", "11110110", "11110101", "11110011", "11110010", "11110000", "11101110", "11101101", "11101011", "11101010", "11101000", "11100111", 
"11100101", "11100100", "11100010", "11100001", "11011111", "11011110", "11011100", "11011011", "11011010", "11011000", "11010111", "11010110", "11010100", "11010011", "11010010", "11010000", "11001111", "11001110", "11001101", "11001011", 
"11001010", "11001001", "11001000", "11000111", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110111", 
"10110110", "10110101", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", 
"10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", 
"01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", 
"01000111", "01000111", "01000110", "01000110", "01000101", "01000101", "01000101", "01000100", "01000100", "01000011", "01000011", "10111101", "10111101", "10111101", "10111100", "10111100", "10111011", "10111011", "10111011", "10111010", 
"10111010", "10111001", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", 
"10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001110", "01001110", "01001101", 
"01001100", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111001", 
"00111000", "00110111", "00110110", "00110101", "00110011", "00110010", "00110001", "00110000", "00101110", "00101101", "00101100", "00101010", "00101001", "00101000", "00100110", "00100101", "00100100", "00100010", "00100001", "00011111", 
"00011110", "00011100", "00011011", "00011001", "00011000", "00010110", "00010101", "00010011", "00010010", "00010000", "00001110", "00001101", "00001011", "00001010", "00001000", "00000110", "00000101", "00000011", "00000010", "00000000", 
"11111110", "11111101", "11111011", "11111010", "11111000", "11110111", "11110101", "11110011", "11110010", "11110000", "11101111", "11101101", "11101100", "11101010", "11101001", "11100111", "11100110", "11100100", "11100011", "11100001", 
"11100000", "11011110", "11011101", "11011100", "11011010", "11011001", "11010111", "11010110", "11010101", "11010011", "11010010", "11010001", "11010000", "11001110", "11001101", "11001100", "11001011", "11001010", "11001000", "11000111", 
"11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110101", "10110100", 
"10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10100111", "10100111", "10100110", 
"01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", 
"01001111", "01001110", "01001110", "01001101", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", 
"01000110", "01000110", "01000101", "01000101", "01000100", "01000100", "01000100", "10111101", "10111100", "10111100", "10111100", "10111011", "10111011", "10111010", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", 
"10110111", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", 
"10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01010111", 
"01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", 
"01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110110", "00110101", "00110100", 
"00110011", "00110010", "00110000", "00101111", "00101110", "00101101", "00101011", "00101010", "00101001", "00100111", "00100110", "00100100", "00100011", "00100010", "00100000", "00011111", "00011101", "00011100", "00011010", "00011001", 
"00010111", "00010110", "00010100", "00010011", "00010001", "00010000", "00001110", "00001101", "00001011", "00001001", "00001000", "00000110", "00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111010", 
"11111000", "11110111", "11110101", "11110100", "11110010", "11110000", "11101111", "11101101", "11101100", "11101010", "11101001", "11100111", "11100110", "11100100", "11100011", "11100010", "11100000", "11011111", "11011101", "11011100", 
"11011011", "11011001", "11011000", "11010111", "11010101", "11010100", "11010011", "11010001", "11010000", "11001111", "11001110", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000100", "11000011", 
"11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110001", 
"10110001", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", 
"01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001111", "01001110", 
"01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000111", "01000110", "01000110", "01000101", 
"01000101", "01000101", "01000100", "10111100", "10111100", "10111011", "10111011", "10111011", "10111010", "10111010", "10111001", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110110", 
"10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", 
"10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", 
"01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", 
"01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110010", "00110001", "00110000", "00101111", 
"00101101", "00101100", "00101011", "00101001", "00101000", "00100111", "00100101", "00100100", "00100011", "00100001", "00100000", "00011110", "00011101", "00011100", "00011010", "00011001", "00010111", "00010110", "00010100", "00010011", 
"00010001", "00010000", "00001110", "00001100", "00001011", "00001001", "00001000", "00000110", "00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111010", "11111000", "11110111", "11110101", "11110100", 
"11110010", "11110001", "11101111", "11101110", "11101100", "11101011", "11101001", "11101000", "11100110", "11100101", "11100011", "11100010", "11100000", "11011111", "11011110", "11011100", "11011011", "11011010", "11011000", "11010111", 
"11010110", "11010100", "11010011", "11010010", "11010001", "11001111", "11001110", "11001101", "11001100", "11001011", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", 
"10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110000", "10110000", "10101111", 
"10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", 
"01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", 
"01001100", "01001100", "01001011", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "01000110", "01000101", "01000101", "10111011", 
"10111011", "10111011", "10111010", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110101", "10110100", "10110100", "10110011", 
"10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", 
"10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", 
"01010000", "01010000", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", 
"00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110101", "00110100", "00110011", "00110010", "00110001", "00101111", "00101110", "00101101", "00101100", "00101010", "00101001", 
"00101000", "00100110", "00100101", "00100100", "00100010", "00100001", "00100000", "00011110", "00011101", "00011011", "00011010", "00011000", "00010111", "00010101", "00010100", "00010010", "00010001", "00001111", "00001110", "00001100", 
"00001011", "00001001", "00001000", "00000110", "00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111010", "11111000", "11110111", "11110101", "11110100", "11110010", "11110001", "11101111", "11101110", 
"11101100", "11101011", "11101001", "11101000", "11100111", "11100101", "11100100", "11100010", "11100001", "11011111", "11011110", "11011101", "11011011", "11011010", "11011001", "11010111", "11010110", "11010101", "11010100", "11010010", 
"11010001", "11010000", "11001111", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111110", "10111101", 
"10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101101", "10101101", 
"10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", 
"01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001100", 
"01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000111", "01000110", "01000110", "01000101", "10111011", "10111011", "10111010", "10111010", "10111001", 
"10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", 
"10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", 
"01001101", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111011", 
"00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110001", "00110000", "00101111", "00101110", "00101100", "00101011", "00101010", "00101001", "00100111", "00100110", "00100101", "00100011", 
"00100010", "00100001", "00011111", "00011110", "00011100", "00011011", "00011001", "00011000", "00010111", "00010101", "00010100", "00010010", "00010001", "00001111", "00001110", "00001100", "00001011", "00001001", "00001000", "00000110", 
"00000101", "00000011", "00000010", "00000000", "11111110", "11111101", "11111011", "11111010", "11111000", "11110111", "11110101", "11110100", "11110010", "11110001", "11110000", "11101110", "11101101", "11101011", "11101010", "11101000", 
"11100111", "11100101", "11100100", "11100011", "11100001", "11100000", "11011110", "11011101", "11011100", "11011010", "11011001", "11011000", "11010111", "11010101", "11010100", "11010011", "11010010", "11010000", "11001111", "11001110", 
"11001101", "11001100", "11001011", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", 
"10101010", "10101010", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", 
"01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", 
"01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01001000", "01000111", "01000111", "01000110", "01000110", "10111010", "10111010", "10111010", "10111001", "10111001", "10111000", "10111000", "10111000", "10110111", 
"10110111", "10110110", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", 
"10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", 
"01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001110", "01001110", "01001101", "01001100", "01001011", "01001011", "01001010", 
"01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", 
"00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101110", "00101101", "00101100", "00101011", "00101001", "00101000", "00100111", "00100110", "00100100", "00100011", "00100010", "00100000", "00011111", "00011101", 
"00011100", "00011011", "00011001", "00011000", "00010110", "00010101", "00010011", "00010010", "00010000", "00001111", "00001110", "00001100", "00001011", "00001001", "00001000", "00000110", "00000101", "00000011", "00000010", "00000000", 
"11111111", "11111101", "11111100", "11111010", "11111001", "11110111", "11110110", "11110100", "11110011", "11110001", "11110000", "11101110", "11101101", "11101011", "11101010", "11101001", "11100111", "11100110", "11100100", "11100011", 
"11100010", "11100000", "11011111", "11011101", "11011100", "11011011", "11011010", "11011000", "11010111", "11010110", "11010100", "11010011", "11010010", "11010001", "11010000", "11001110", "11001101", "11001100", "11001011", "11001010", 
"11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", 
"10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", 
"10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", 
"01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001011", "01001010", "01001010", "01001001", 
"01001001", "01001001", "01001000", "01001000", "01000111", "01000111", "01000111", "10111010", "10111001", "10111001", "10111001", "10111000", "10111000", "10110111", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", 
"10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", 
"10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010110", "01010110", "01010101", "01010101", 
"01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", 
"01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", 
"00110000", "00101111", "00101110", "00101101", "00101100", "00101010", "00101001", "00101000", "00100110", "00100101", "00100100", "00100011", "00100001", "00100000", "00011110", "00011101", "00011100", "00011010", "00011001", "00010111", 
"00010110", "00010101", "00010011", "00010010", "00010000", "00001111", "00001101", "00001100", "00001010", "00001001", "00000111", "00000110", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111010", 
"11111001", "11110111", "11110110", "11110100", "11110011", "11110001", "11110000", "11101110", "11101101", "11101100", "11101010", "11101001", "11100111", "11100110", "11100101", "11100011", "11100010", "11100001", "11011111", "11011110", 
"11011101", "11011011", "11011010", "11011001", "11010111", "11010110", "11010101", "11010100", "11010011", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001010", "11001001", "11001000", "11000111", "11000110", 
"11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110100", 
"10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", 
"10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", 
"01010000", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001010", "01001001", "01001001", "01001000", 
"01001000", "01001000", "01000111", "10111001", "10111001", "10111000", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110100", "10110011", "10110011", 
"10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", 
"10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010010", 
"01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", 
"01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101101", "00101100", 
"00101011", "00101010", "00101001", "00100111", "00100110", "00100101", "00100011", "00100010", "00100001", "00011111", "00011110", "00011101", "00011011", "00011010", "00011001", "00010111", "00010110", "00010100", "00010011", "00010010", 
"00010000", "00001111", "00001101", "00001100", "00001010", "00001001", "00000111", "00000110", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111010", "11111001", "11110111", "11110110", "11110100", 
"11110011", "11110001", "11110000", "11101111", "11101101", "11101100", "11101010", "11101001", "11101000", "11100110", "11100101", "11100100", "11100010", "11100001", "11100000", "11011110", "11011101", "11011100", "11011010", "11011001", 
"11011000", "11010111", "11010101", "11010100", "11010011", "11010010", "11010001", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", 
"11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110011", "10110011", "10110010", 
"10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", 
"01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010001", "01010000", "01010000", 
"01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001001", "01001000", "01001000", "10111001", 
"10111000", "10111000", "10110111", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", 
"10110000", "10101111", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", 
"01001101", "01001101", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", 
"00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00101111", "00101110", "00101101", "00101100", "00101011", "00101001", "00101000", "00100111", 
"00100110", "00100100", "00100011", "00100010", "00100000", "00011111", "00011110", "00011100", "00011011", "00011010", "00011000", "00010111", "00010110", "00010100", "00010011", "00010001", "00010000", "00001111", "00001101", "00001100", 
"00001010", "00001001", "00000111", "00000110", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111010", "11111001", "11110111", "11110110", "11110101", "11110011", "11110010", "11110000", "11101111", 
"11101101", "11101100", "11101011", "11101001", "11101000", "11100111", "11100101", "11100100", "11100011", "11100001", "11100000", "11011111", "11011101", "11011100", "11011011", "11011001", "11011000", "11010111", "11010110", "11010101", 
"11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", 
"10111110", "10111110", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", 
"10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", 
"01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", 
"01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001010", "01001001", "01001001", "01001000", "10111000", "10111000", "10110111", "10110111", "10110110", 
"10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", 
"10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", 
"01010111", "01010111", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001100", "01001011", "01001011", 
"01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", 
"00111000", "00110111", "00110110", "00110101", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101011", "00101010", "00101001", "00101000", "00100111", "00100101", "00100100", "00100011", "00100001", 
"00100000", "00011111", "00011101", "00011100", "00011011", "00011001", "00011000", "00010111", "00010101", "00010100", "00010011", "00010001", "00010000", "00001110", "00001101", "00001011", "00001010", "00001001", "00000111", "00000110", 
"00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111010", "11111001", "11110111", "11110110", "11110101", "11110011", "11110010", "11110000", "11101111", "11101110", "11101100", "11101011", "11101010", 
"11101000", "11100111", "11100101", "11100100", "11100011", "11100010", "11100000", "11011111", "11011110", "11011100", "11011011", "11011010", "11011001", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010000", 
"11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", 
"10111100", "10111011", "10111010", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101110", 
"10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", 
"01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001111", "01001110", "01001110", "01001101", 
"01001101", "01001100", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001010", "01001001", "01001001", "10110111", "10110111", "10110111", "10110110", "10110110", "10110110", "10110101", "10110101", "10110100", 
"10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", 
"10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010101", "01010101", 
"01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", 
"01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", 
"00110011", "00110010", "00110001", "00110000", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00100111", "00100110", "00100101", "00100100", "00100010", "00100001", "00100000", "00011110", "00011101", "00011100", 
"00011011", "00011001", "00011000", "00010110", "00010101", "00010100", "00010010", "00010001", "00010000", "00001110", "00001101", "00001011", "00001010", "00001001", "00000111", "00000110", "00000100", "00000011", "00000001", "00000000", 
"11111111", "11111101", "11111100", "11111010", "11111001", "11111000", "11110110", "11110101", "11110011", "11110010", "11110001", "11101111", "11101110", "11101100", "11101011", "11101010", "11101000", "11100111", "11100110", "11100100", 
"11100011", "11100010", "11100001", "11011111", "11011110", "11011101", "11011100", "11011010", "11011001", "11011000", "11010111", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001100", 
"11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101100", 
"10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", 
"01010100", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001101", "01001100", 
"01001100", "01001011", "01001011", "01001011", "01001010", "01001010", "01001001", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110011", "10110010", 
"10110010", "10110001", "10110001", "10110000", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", 
"10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", 
"01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", 
"01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110010", "00110001", "00110000", "00101111", 
"00101110", "00101101", "00101100", "00101011", "00101001", "00101000", "00100111", "00100110", "00100100", "00100011", "00100010", "00100001", "00011111", "00011110", "00011101", "00011100", "00011010", "00011001", "00011000", "00010110", 
"00010101", "00010100", "00010010", "00010001", "00001111", "00001110", "00001101", "00001011", "00001010", "00001000", "00000111", "00000110", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111010", 
"11111001", "11111000", "11110110", "11110101", "11110100", "11110010", "11110001", "11101111", "11101110", "11101101", "11101011", "11101010", "11101001", "11100111", "11100110", "11100101", "11100011", "11100010", "11100001", "11100000", 
"11011110", "11011101", "11011100", "11011011", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", 
"11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", 
"10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", 
"10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", 
"01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001100", "01001011", 
"01001011", "01001010", "01001010", "10110110", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", 
"10101111", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", 
"01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000000", "00111111", 
"00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101100", "00101011", "00101010", 
"00101001", "00101000", "00100111", "00100101", "00100100", "00100011", "00100010", "00100000", "00011111", "00011110", "00011101", "00011011", "00011010", "00011001", "00010111", "00010110", "00010101", "00010011", "00010010", "00010001", 
"00001111", "00001110", "00001100", "00001011", "00001010", "00001000", "00000111", "00000110", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111010", "11111001", "11111000", "11110110", "11110101", 
"11110100", "11110010", "11110001", "11110000", "11101110", "11101101", "11101100", "11101010", "11101001", "11101000", "11100110", "11100101", "11100100", "11100010", "11100001", "11100000", "11011111", "11011101", "11011100", "11011011", 
"11011010", "11011001", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", 
"11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", 
"10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", 
"10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", 
"01010010", "01010001", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001100", "01001011", "01001011", "01001011", "10110110", 
"10110101", "10110101", "10110101", "10110100", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101111", "10101110", "10101110", 
"10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", 
"01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001100", "01001011", 
"01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111011", 
"00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00100111", "00100110", "00100101", 
"00100100", "00100011", "00100001", "00100000", "00011111", "00011110", "00011100", "00011011", "00011010", "00011000", "00010111", "00010110", "00010100", "00010011", "00010010", "00010000", "00001111", "00001110", "00001100", "00001011", 
"00001010", "00001000", "00000111", "00000110", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111011", "11111001", "11111000", "11110110", "11110101", "11110100", "11110010", "11110001", "11110000", 
"11101110", "11101101", "11101100", "11101010", "11101001", "11101000", "11100111", "11100101", "11100100", "11100011", "11100010", "11100000", "11011111", "11011110", "11011101", "11011011", "11011010", "11011001", "11011000", "11010111", 
"11010110", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", 
"11000001", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", 
"10110010", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010010", "01010001", 
"01010001", "01010000", "01010000", "01001111", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "10110101", "10110101", "10110101", "10110100", "10110100", 
"10110011", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", 
"10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", 
"01010101", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", 
"01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", 
"00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100011", "00100010", "00100001", "00100000", 
"00011110", "00011101", "00011100", "00011011", "00011001", "00011000", "00010111", "00010110", "00010100", "00010011", "00010010", "00010000", "00001111", "00001110", "00001100", "00001011", "00001010", "00001000", "00000111", "00000101", 
"00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111011", "11111001", "11111000", "11110111", "11110101", "11110100", "11110011", "11110001", "11110000", "11101111", "11101101", "11101100", "11101011", 
"11101001", "11101000", "11100111", "11100110", "11100100", "11100011", "11100010", "11100001", "11011111", "11011110", "11011101", "11011100", "11011011", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", 
"11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000000", "10111111", 
"10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", 
"10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", 
"01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", 
"01010000", "01001111", "01001111", "01001110", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001100", "10110101", "10110100", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110010", 
"10110001", "10110001", "10110000", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", 
"10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", "01010010", 
"01010010", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01000111", "01000111", "01000110", "01000101", "01000100", 
"01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", 
"00110001", "00110000", "00101111", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100101", "00100100", "00100011", "00100010", "00100001", "00011111", "00011110", "00011101", "00011100", "00011010", 
"00011001", "00011000", "00010111", "00010101", "00010100", "00010011", "00010001", "00010000", "00001111", "00001101", "00001100", "00001011", "00001001", "00001000", "00000111", "00000101", "00000100", "00000011", "00000001", "00000000", 
"11111111", "11111101", "11111100", "11111011", "11111001", "11111000", "11110111", "11110101", "11110100", "11110011", "11110001", "11110000", "11101111", "11101101", "11101100", "11101011", "11101010", "11101000", "11100111", "11100110", 
"11100101", "11100011", "11100010", "11100001", "11100000", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", 
"11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111101", "10111100", 
"10111011", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", 
"10101110", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", 
"01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01010000", "01001111", "01001111", 
"01001110", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "10110100", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10110000", 
"10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01001111", 
"01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000010", "01000001", "01000000", 
"01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", 
"00101100", "00101011", "00101010", "00101001", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100000", "00011111", "00011110", "00011101", "00011011", "00011010", "00011001", "00011000", "00010110", "00010101", 
"00010100", "00010011", "00010001", "00010000", "00001111", "00001101", "00001100", "00001011", "00001001", "00001000", "00000111", "00000101", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111011", 
"11111001", "11111000", "11110111", "11110101", "11110100", "11110011", "11110010", "11110000", "11101111", "11101110", "11101100", "11101011", "11101010", "11101001", "11100111", "11100110", "11100101", "11100100", "11100010", "11100001", 
"11100000", "11011111", "11011110", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", 
"11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101100", 
"10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", 
"01010110", "01010101", "01010101", "01010100", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001111", "01001110", "01001110", 
"01001101", "01001101", "01001101", "10110100", "10110011", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101111", "10101110", "10101110", "10101101", 
"10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", 
"01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", 
"01001100", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", 
"00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101010", "00101001", "00101000", 
"00100111", "00100110", "00100101", "00100100", "00100010", "00100001", "00100000", "00011111", "00011110", "00011100", "00011011", "00011010", "00011001", "00010111", "00010110", "00010101", "00010100", "00010010", "00010001", "00010000", 
"00001110", "00001101", "00001100", "00001011", "00001001", "00001000", "00000111", "00000101", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111011", "11111001", "11111000", "11110111", "11110110", 
"11110100", "11110011", "11110010", "11110000", "11101111", "11101110", "11101101", "11101011", "11101010", "11101001", "11101000", "11100110", "11100101", "11100100", "11100011", "11100001", "11100000", "11011111", "11011110", "11011101", 
"11011100", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", 
"11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", 
"10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", 
"10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", 
"01010100", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "10110011", 
"10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", 
"10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", 
"01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", 
"01001000", "01000111", "01000111", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", 
"00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100100", "00100011", 
"00100010", "00100001", "00100000", "00011111", "00011101", "00011100", "00011011", "00011010", "00011000", "00010111", "00010110", "00010101", "00010011", "00010010", "00010001", "00010000", "00001110", "00001101", "00001100", "00001010", 
"00001001", "00001000", "00000111", "00000101", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111011", "11111010", "11111000", "11110111", "11110110", "11110100", "11110011", "11110010", "11110001", 
"11101111", "11101110", "11101101", "11101100", "11101010", "11101001", "11101000", "11100111", "11100101", "11100100", "11100011", "11100010", "11100001", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", 
"11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", 
"11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110101", "10110101", 
"10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", 
"10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010100", 
"01010011", "01010011", "01010010", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001110", "10110011", "10110010", "10110010", "10110010", "10110001", 
"10110001", "10110000", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", 
"10101000", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", 
"01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000101", 
"01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", 
"00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00011111", "00011110", 
"00011101", "00011100", "00011011", "00011001", "00011000", "00010111", "00010110", "00010100", "00010011", "00010010", "00010001", "00001111", "00001110", "00001101", "00001100", "00001010", "00001001", "00001000", "00000110", "00000101", 
"00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111011", "11111010", "11111000", "11110111", "11110110", "11110101", "11110011", "11110010", "11110001", "11101111", "11101110", "11101101", "11101100", 
"11101011", "11101001", "11101000", "11100111", "11100110", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", 
"11010100", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", 
"11000001", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", 
"10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", 
"10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", 
"01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "10110010", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10110000", "10101111", 
"10101111", "10101110", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", 
"01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000011", "01000010", 
"01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", 
"00101111", "00101110", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011010", "00011001", 
"00011000", "00010111", "00010101", "00010100", "00010011", "00010010", "00010001", "00001111", "00001110", "00001101", "00001011", "00001010", "00001001", "00001000", "00000110", "00000101", "00000100", "00000011", "00000001", "00000000", 
"11111111", "11111101", "11111100", "11111011", "11111010", "11111000", "11110111", "11110110", "11110101", "11110011", "11110010", "11110001", "11110000", "11101110", "11101101", "11101100", "11101011", "11101010", "11101000", "11100111", 
"11100110", "11100101", "11100100", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", 
"11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "10111111", "10111111", 
"10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", 
"10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", 
"01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", 
"01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001111", "10110010", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", 
"10101101", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", 
"01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", 
"01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01000111", "01000111", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111110", 
"00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", 
"00101010", "00101001", "00101000", "00100111", "00100110", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011100", "00011011", "00011010", "00011001", "00011000", "00010110", "00010101", "00010100", 
"00010011", "00010010", "00010000", "00001111", "00001110", "00001101", "00001011", "00001010", "00001001", "00001000", "00000110", "00000101", "00000100", "00000011", "00000001", "00000000", "11111111", "11111101", "11111100", "11111011", 
"11111010", "11111000", "11110111", "11110110", "11110101", "11110011", "11110010", "11110001", "11110000", "11101111", "11101101", "11101100", "11101011", "11101010", "11101001", "11100111", "11100110", "11100101", "11100100", "11100011", 
"11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", 
"11001100", "11001011", "11001010", "11001001", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", 
"10111011", "10111011", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", 
"10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", 
"01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010001", "01010000", 
"01010000", "01001111", "01001111", "10110001", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", 
"10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", 
"01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", 
"01001001", "01001000", "01001000", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111010", 
"00111001", "00111000", "00110111", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00100111", "00100110", 
"00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011101", "00011100", "00011011", "00011010", "00011001", "00010111", "00010110", "00010101", "00010100", "00010011", "00010001", "00010000", "00001111", 
"00001110", "00001101", "00001011", "00001010", "00001001", "00001000", "00000110", "00000101", "00000100", "00000011", "00000001", "00000000", "11111111", "11111110", "11111100", "11111011", "11111010", "11111001", "11110111", "11110110", 
"11110101", "11110100", "11110010", "11110001", "11110000", "11101111", "11101110", "11101100", "11101011", "11101010", "11101001", "11101000", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011110", 
"11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", 
"11001001", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", 
"10101101", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", 
"01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010001", "01010000", "01010000", "01010000", "10110001", 
"10110000", "10110000", "10110000", "10101111", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", 
"10101000", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010011", "01010011", 
"01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000110", 
"01000110", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", 
"00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", 
"00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011000", "00010111", "00010110", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", "00001110", "00001100", "00001011", "00001010", 
"00001001", "00000111", "00000110", "00000101", "00000100", "00000010", "00000001", "00000000", "11111111", "11111110", "11111100", "11111011", "11111010", "11111001", "11110111", "11110110", "11110101", "11110100", "11110011", "11110001", 
"11110000", "11101111", "11101110", "11101101", "11101011", "11101010", "11101001", "11101000", "11100111", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011100", "11011011", "11011010", 
"11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001001", "11001000", "11000111", 
"11000110", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", 
"10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101100", "10101100", "10101011", 
"10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", 
"01010110", "01010101", "01010101", "01010100", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "10110000", "10110000", "10110000", "10101111", "10101111", 
"10101110", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", 
"01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", 
"01000010", "01000001", "01000001", "01000000", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00110111", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", 
"00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", 
"00011100", "00011011", "00011001", "00011000", "00010111", "00010110", "00010101", "00010011", "00010010", "00010001", "00010000", "00001111", "00001101", "00001100", "00001011", "00001010", "00001001", "00000111", "00000110", "00000101", 
"00000100", "00000010", "00000001", "00000000", "11111111", "11111110", "11111100", "11111011", "11111010", "11111001", "11110111", "11110110", "11110101", "11110100", "11110011", "11110001", "11110000", "11101111", "11101110", "11101101", 
"11101100", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11010111", "11010110", 
"11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", 
"11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", 
"10110100", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", 
"10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", 
"01010100", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010010", "01010001", "01010001", "01010000", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101110", "10101101", "10101101", 
"10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", 
"01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001101", 
"01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000000", "00111111", 
"00111111", "00111110", "00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110001", "00110000", "00101111", "00101110", 
"00101101", "00101100", "00101011", "00101010", "00101001", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011011", "00011010", "00011001", "00011000", 
"00010111", "00010110", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001101", "00001100", "00001011", "00001010", "00001001", "00000111", "00000110", "00000101", "00000100", "00000010", "00000001", "00000000", 
"11111111", "11111110", "11111100", "11111011", "11111010", "11111001", "11111000", "11110110", "11110101", "11110100", "11110011", "11110010", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101001", "11101000", 
"11100111", "11100110", "11100101", "11100100", "11100011", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", 
"11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001001", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", 
"11000000", "10111111", "10111111", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", 
"10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", 
"10101000", "10101000", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010100", 
"01010011", "01010011", "01010010", "01010010", "01010010", "01010001", "01010001", "10101111", "10101111", "10101111", "10101110", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", 
"10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", 
"01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001010", 
"01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111110", "00111101", "00111101", "00111100", 
"00111011", "00111010", "00111001", "00111000", "00110111", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", 
"00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010101", "00010100", "00010011", 
"00010010", "00010001", "00010000", "00001110", "00001101", "00001100", "00001011", "00001010", "00001000", "00000111", "00000110", "00000101", "00000100", "00000010", "00000001", "00000000", "11111111", "11111110", "11111100", "11111011", 
"11111010", "11111001", "11111000", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101000", "11100111", "11100110", "11100101", "11100100", 
"11100011", "11100010", "11100001", "11100000", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", 
"11001110", "11001101", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111110", 
"10111110", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", 
"10110001", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", 
"10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010100", "01010011", "01010011", "01010011", 
"01010010", "01010010", "01010001", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", 
"10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", 
"01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01000111", 
"01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", 
"00110111", "00110110", "00110101", "00110100", "00110011", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", 
"00100100", "00100011", "00100010", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00001111", "00001110", 
"00001101", "00001100", "00001011", "00001010", "00001000", "00000111", "00000110", "00000101", "00000100", "00000010", "00000001", "00000000", "11111111", "11111110", "11111100", "11111011", "11111010", "11111001", "11111000", "11110111", 
"11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", 
"11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010110", "11010101", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", 
"11001011", "11001010", "11001001", "11001000", "11001000", "11000111", "11000110", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", 
"10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110000", "10110000", "10101111", 
"10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", 
"01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "10101111", 
"10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", 
"01010000", "01010000", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", 
"01000011", "01000011", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", "00111010", "00111001", "00111000", "00111000", "00110111", "00110110", "00110101", "00110100", 
"00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101011", "00101010", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", 
"00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001001", 
"00001000", "00000111", "00000110", "00000101", "00000100", "00000010", "00000001", "00000000", "11111111", "11111110", "11111100", "11111011", "11111010", "11111001", "11111000", "11110111", "11110101", "11110100", "11110011", "11110010", 
"11110001", "11110000", "11101111", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", 
"11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001100", "11001011", "11001010", "11001001", 
"11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", 
"10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", 
"01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "10101110", "10101110", "10101101", "10101101", "10101101", 
"10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", 
"01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", 
"01001101", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000001", "01000001", 
"01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110100", "00110100", "00110011", "00110010", "00110001", "00110000", 
"00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", 
"00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001001", "00001000", "00000111", "00000110", "00000101", 
"00000100", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111011", "11111010", "11111001", "11111000", "11110111", "11110110", "11110100", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", 
"11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", 
"11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11001000", "11000111", "11000110", 
"11000101", "11000100", "11000100", "11000011", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", 
"10110111", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", 
"10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", 
"01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101011", 
"10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", 
"01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", 
"01001011", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111101", 
"00111100", "00111100", "00111011", "00111010", "00111001", "00111000", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00110000", "00101111", "00101110", "00101101", "00101100", 
"00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", 
"00010110", "00010101", "00010100", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000011", "00000010", "00000001", "00000000", 
"11111111", "11111110", "11111101", "11111011", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101011", "11101010", "11101001", 
"11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011010", "11011001", "11011000", "11011000", "11010111", "11010110", "11010101", 
"11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", 
"11000010", "11000010", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110101", 
"10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", 
"10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", 
"01010101", "01010101", "01010101", "01010100", "01010100", "01010100", "01010011", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", 
"10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010100", 
"01010011", "01010011", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", 
"01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111010", "00111010", 
"00111001", "00111000", "00110111", "00110110", "00110101", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00101000", 
"00100111", "00100110", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010011", "00010010", 
"00010001", "00010000", "00001111", "00001110", "00001101", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111011", 
"11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101001", "11101000", "11100111", "11100110", "11100101", 
"11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", 
"11010000", "11001111", "11001110", "11001110", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11001000", "11000111", "11000110", "11000101", "11000100", "11000100", "11000011", "11000010", "11000001", "11000001", 
"11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110011", 
"10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", 
"10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", 
"01010100", "01010100", "01010100", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", 
"01010001", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", 
"01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111001", "00111000", "00111000", "00110111", "00110110", 
"00110101", "00110100", "00110011", "00110010", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", 
"00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", 
"00001101", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111011", "11111010", "11111001", "11111000", "11110111", 
"11110110", "11110101", "11110100", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", 
"11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010010", "11010001", "11010000", "11001111", "11001110", 
"11001101", "11001100", "11001011", "11001011", "11001010", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", 
"10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", 
"10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", 
"10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "10101100", 
"10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", 
"01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001110", 
"01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", 
"01000001", "01000000", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110110", "00110101", "00110101", "00110100", "00110011", "00110010", 
"00110001", "00110000", "00101111", "00101110", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", 
"00011110", "00011101", "00011100", "00011011", "00011010", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001100", "00001011", "00001010", "00001001", 
"00001000", "00000111", "00000110", "00000101", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110100", "11110011", 
"11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", 
"11011100", "11011011", "11011010", "11011001", "11011000", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001101", "11001100", "11001011", 
"11001010", "11001001", "11001000", "11001000", "11000111", "11000110", "11000101", "11000100", "11000100", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111100", "10111100", 
"10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10110000", 
"10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "10101100", "10101100", "10101011", "10101011", "10101010", 
"10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", 
"01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", "01001100", 
"01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", 
"00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111001", "00111000", "00111000", "00110111", "00110110", "00110101", "00110100", "00110011", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", 
"00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011100", "00011011", "00011010", 
"00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000100", 
"00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11101111", "11101110", 
"11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", 
"11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11010000", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001010", "11001001", "11001000", 
"11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", 
"10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", 
"01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101001", 
"10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", 
"01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", 
"01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", 
"00111010", "00111010", "00111001", "00111000", "00110111", "00110110", "00110110", "00110101", "00110100", "00110011", "00110010", "00110001", "00110000", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", 
"00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", 
"00010101", "00010100", "00010011", "00010010", "00010001", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000100", "00000011", "00000010", "00000001", "00000000", 
"11111111", "11111110", "11111101", "11111100", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101110", "11101101", "11101100", "11101011", "11101010", 
"11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", 
"11010101", "11010100", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001101", "11001101", "11001100", "11001011", "11001010", "11001001", "11001000", "11001000", "11000111", "11000110", "11000101", 
"11000100", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10110111", 
"10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", 
"10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", 
"01010111", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", 
"01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", 
"01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111001", "00111000", "00111000", 
"00110111", "00110110", "00110101", "00110100", "00110011", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", 
"00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", 
"00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000100", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", 
"11111011", "11111001", "11111000", "11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", 
"11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", 
"11010010", "11010001", "11010000", "11001111", "11001111", "11001110", "11001101", "11001100", "11001011", "11001010", "11001010", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000011", 
"11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110110", 
"10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", 
"10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", 
"01010110", "01010110", "01010110", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", 
"01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", 
"01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", 
"01000010", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110110", "00110110", "00110101", "00110100", 
"00110011", "00110010", "00110001", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", 
"00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", 
"00001100", "00001011", "00001010", "00001001", "00001000", "00000111", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111011", "11111001", "11111000", "11110111", 
"11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100110", "11100101", "11100100", "11100011", "11100010", 
"11100001", "11100000", "11011111", "11011110", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010010", "11010001", "11010000", 
"11001111", "11001110", "11001101", "11001100", "11001100", "11001011", "11001010", "11001001", "11001000", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", 
"10111111", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110100", 
"10110011", "10110011", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", 
"10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "10101010", 
"10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", 
"01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001101", "01001101", "01001100", 
"01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000001", "01000000", 
"00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111000", "00111000", "00110111", "00110110", "00110101", "00110100", "00110100", "00110011", "00110010", "00110001", "00110000", 
"00101111", "00101110", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100010", "00100001", "00100000", "00011111", "00011110", 
"00011101", "00011100", "00011011", "00011010", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", 
"00001000", "00000111", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111011", "11111010", "11111000", "11110111", "11110110", "11110101", "11110100", "11110011", 
"11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", 
"11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001110", "11001101", 
"11001100", "11001011", "11001010", "11001010", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111111", "10111110", 
"10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", 
"10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", 
"10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "10101010", "10101010", "10101001", "10101001", "10101000", 
"10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", 
"01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", 
"01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111101", 
"00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110110", "00110110", "00110101", "00110100", "00110011", "00110010", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", 
"00101011", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", 
"00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", "00000110", "00000101", "00000100", 
"00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111011", "11111010", "11111001", "11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101111", 
"11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", 
"11011010", "11011001", "11011000", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010000", "11010000", "11001111", "11001110", "11001101", "11001100", "11001100", "11001011", "11001010", 
"11001001", "11001000", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", 
"10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", 
"10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", 
"10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", 
"01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", 
"01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111011", "00111010", "00111001", 
"00111000", "00111000", "00110111", "00110110", "00110101", "00110100", "00110100", "00110011", "00110010", "00110001", "00110000", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", 
"00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", 
"00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", 
"11111111", "11111110", "11111101", "11111100", "11111011", "11111010", "11111001", "11111000", "11110111", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", 
"11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011100", "11011011", "11011010", "11011001", "11011000", 
"11010111", "11010110", "11010101", "11010100", "11010011", "11010011", "11010010", "11010001", "11010000", "11001111", "11001110", "11001110", "11001101", "11001100", "11001011", "11001010", "11001010", "11001001", "11001000", "11000111", 
"11000110", "11000110", "11000101", "11000100", "11000100", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", 
"10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", 
"01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", 
"01011000", "01010111", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", 
"01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", 
"01000011", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110110", "00110110", 
"00110101", "00110100", "00110011", "00110010", "00110010", "00110001", "00110000", "00101111", "00101110", "00101101", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", 
"00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", 
"00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001001", "00001000", "00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", 
"11111011", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", 
"11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010101", 
"11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001111", "11001110", "11001101", "11001100", "11001011", "11001011", "11001010", "11001001", "11001000", "11001000", "11000111", "11000110", "11000101", "11000101", 
"11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10111000", 
"10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", 
"10101101", "10101100", "10101100", "10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101001", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", 
"01011000", "01011000", "01011000", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01010111", "01010111", "01010111", "01010110", 
"01010110", "01010101", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", 
"01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000010", "01000010", "01000001", 
"01000000", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111000", "00111000", "00110111", "00110110", "00110101", "00110101", "00110100", "00110011", "00110010", 
"00110001", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101011", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", 
"00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", 
"00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111011", "11111010", "11111001", "11111000", 
"11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100111", "11100110", "11100101", "11100100", 
"11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", "11011000", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010010", 
"11010001", "11010000", "11001111", "11001110", "11001101", "11001101", "11001100", "11001011", "11001010", "11001001", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000100", "11000011", "11000010", 
"11000001", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111101", "10111100", "10111100", "10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110110", 
"10110101", "10110101", "10110100", "10110100", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", 
"10101011", "10101011", "10101011", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "10101000", 
"10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010101", "01010101", "01010101", "01010100", 
"01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", 
"01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", 
"00111101", "00111100", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110111", "00110110", "00110101", "00110100", "00110011", "00110011", "00110010", "00110001", "00110000", "00101111", "00101110", 
"00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", 
"00011011", "00011010", "00011001", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", 
"00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111011", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110100", 
"11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", 
"11011111", "11011110", "11011101", "11011100", "11011011", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010101", "11010100", "11010100", "11010011", "11010010", "11010001", "11010000", "11001111", "11001111", 
"11001110", "11001101", "11001100", "11001011", "11001011", "11001010", "11001001", "11001000", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000001", "11000000", 
"10111111", "10111111", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111010", "10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110100", "10110100", 
"10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", 
"10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "10101000", "10101000", "10100111", "10100111", "10100111", 
"10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010010", "01010010", 
"01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01001000", 
"01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", "00111011", 
"00111010", "00111001", "00111000", "00111000", "00110111", "00110110", "00110101", "00110101", "00110100", "00110011", "00110010", "00110001", "00110001", "00110000", "00101111", "00101110", "00101101", "00101100", "00101100", "00101011", 
"00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", 
"00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000100", 
"00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111011", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", 
"11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011110", "11011101", 
"11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010110", "11010101", "11010100", "11010011", "11010010", "11010001", "11010001", "11010000", "11001111", "11001110", "11001101", "11001101", "11001100", 
"11001011", "11001010", "11001001", "11001001", "11001000", "11000111", "11000110", "11000110", "11000101", "11000100", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", 
"10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10111000", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", 
"10110010", "10110001", "10110001", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", 
"10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", 
"01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", 
"01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001000", "01001000", "01000111", "01000111", "01000110", "01000101", "01000101", 
"01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", "00111110", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", 
"00110111", "00110110", "00110101", "00110100", "00110011", "00110011", "00110010", "00110001", "00110000", "00101111", "00101111", "00101110", "00101101", "00101100", "00101011", "00101010", "00101010", "00101001", "00101000", "00100111", 
"00100110", "00100101", "00100100", "00100011", "00100010", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", 
"00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", 
"11111111", "11111110", "11111101", "11111100", "11111011", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", 
"11101011", "11101010", "11101001", "11101000", "11100111", "11100110", "11100101", "11100100", "11100011", "11100010", "11100001", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011001", 
"11011000", "11011000", "11010111", "11010110", "11010101", "11010100", "11010011", "11010010", "11010010", "11010001", "11010000", "11001111", "11001110", "11001110", "11001101", "11001100", "11001011", "11001011", "11001010", "11001001", 
"11001000", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", "11000011", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111111", "10111110", "10111101", "10111101", "10111100", "10111100", 
"10111011", "10111010", "10111010", "10111001", "10111001", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", 
"10110000", "10110000", "10101111", "10101111", "10101110", "10101110", "10101101", "10101101", "10101101", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", 
"10101000", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "10100111", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", 
"01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010011", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", 
"01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001010", "01001001", "01001001", "01001000", "01000111", "01000111", "01000110", "01000110", "01000101", "01000100", "01000100", "01000011", "01000011", "01000010", 
"01000001", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111101", "00111100", "00111011", "00111011", "00111010", "00111001", "00111000", "00111000", "00110111", "00110110", "00110101", "00110101", "00110100", 
"00110011", "00110010", "00110010", "00110001", "00110000", "00101111", "00101110", "00101110", "00101101", "00101100", "00101011", "00101010", "00101001", "00101000", "00101000", "00100111", "00100110", "00100101", "00100100", "00100011", 
"00100010", "00100001", "00100000", "00011111", "00011111", "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", 
"00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", 
"11111011", "11111010", "11111001", "11111000", "11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", 
"11100111", "11100110", "11100101", "11100100", "11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011011", "11011010", "11011010", "11011001", "11011000", "11010111", "11010110", 
"11010101", "11010100", "11010100", "11010011", "11010010", "11010001", "11010000", "11010000", "11001111", "11001110", "11001101", "11001100", "11001100", "11001011", "11001010", "11001001", "11001001", "11001000", "11000111", "11000110", 
"11000110", "11000101", "11000100", "11000100", "11000011", "11000010", "11000010", "11000001", "11000000", "11000000", "10111111", "10111110", "10111110", "10111101", "10111101", "10111100", "10111011", "10111011", "10111010", "10111010", 
"10111001", "10111000", "10111000", "10110111", "10110111", "10110110", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10101111", 
"10101111", "10101110", "10101110", "10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", 
"10100111", "10100110", "01011001", "10100111", "10100111", "10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", 
"01010100", "01010100", "01010011", "01010011", "01010010", "01010010", "01010001", "01010001", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", 
"01001010", "01001010", "01001001", "01001001", "01001000", "01001000", "01000111", "01000110", "01000110", "01000101", "01000101", "01000100", "01000011", "01000011", "01000010", "01000010", "01000001", "01000000", "01000000", "00111111", 
"00111110", "00111110", "00111101", "00111100", "00111100", "00111011", "00111010", "00111010", "00111001", "00111000", "00110111", "00110111", "00110110", "00110101", "00110100", "00110100", "00110011", "00110010", "00110001", "00110000", 
"00110000", "00101111", "00101110", "00101101", "00101100", "00101100", "00101011", "00101010", "00101001", "00101000", "00100111", "00100110", "00100110", "00100101", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", 
"00011110", "00011101", "00011100", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", 
"00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "11111111", "11111110", "11111101", "11111100", "11111011", "11111010", "11111001", "11111000", 
"11110111", "11110110", "11110101", "11110100", "11110011", "11110010", "11110001", "11110000", "11101111", "11101110", "11101101", "11101100", "11101011", "11101010", "11101001", "11101000", "11100111", "11100111", "11100110", "11100101", 
"11100100", "11100011", "11100010", "11100001", "11100000", "11011111", "11011110", "11011101", "11011100", "11011100", "11011011", "11011010", "11011001", "11011000", "11010111", "11010110", "11010110", "11010101", "11010100", "11010011", 
"11010010", "11010001", "11010001", "11010000", "11001111", "11001110", "11001110", "11001101", "11001100", "11001011", "11001010", "11001010", "11001001", "11001000", "11001000", "11000111", "11000110", "11000101", "11000101", "11000100", 
"11000011", "11000011", "11000010", "11000001", "11000001", "11000000", "10111111", "10111111", "10111110", "10111110", "10111101", "10111100", "10111100", "10111011", "10111011", "10111010", "10111001", "10111001", "10111000", "10111000", 
"10110111", "10110111", "10110110", "10110101", "10110101", "10110100", "10110100", "10110011", "10110011", "10110010", "10110010", "10110001", "10110001", "10110000", "10110000", "10110000", "10101111", "10101111", "10101110", "10101110", 
"10101101", "10101101", "10101100", "10101100", "10101100", "10101011", "10101011", "10101010", "10101010", "10101010", "10101001", "10101001", "10101000", "10101000", "10101000", "10100111", "10100111", "10100111", "10100110", "10100111", 
"10100110", "01011001", "01011001", "01011001", "01011000", "01011000", "01011000", "01010111", "01010111", "01010110", "01010110", "01010110", "01010101", "01010101", "01010100", "01010100", "01010100", "01010011", "01010011", "01010010", 
"01010010", "01010001", "01010001", "01010000", "01010000", "01010000", "01001111", "01001111", "01001110", "01001110", "01001101", "01001101", "01001100", "01001100", "01001011", "01001011", "01001010", "01001001", "01001001", "01001000", 
"01001000", "01000111", "01000111", "01000110", "01000101", "01000101", "01000100", "01000100", "01000011", "01000010", "01000010", "01000001", "01000001", "01000000", "00111111", "00111111", "00111110", "00111101", "00111101", "00111100", 
"00111011", "00111011", "00111010", "00111001", "00111000", "00111000", "00110111", "00110110", "00110110", "00110101", "00110100", "00110011", "00110010", "00110010", "00110001", "00110000", "00101111", "00101111", "00101110", "00101101", 
"00101100", "00101011", "00101010", "00101010", "00101001", "00101000", "00100111", "00100110", "00100101", "00100100", "00100100", "00100011", "00100010", "00100001", "00100000", "00011111", "00011110", "00011101", "00011100", "00011011", 
"00011010", "00011001", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", 
"00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", 
"00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", 
"00100000", "00100001", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101101", "00101110", "00101111", "00110000", 
"00110001", "00110001", "00110010", "00110011", "00110100", "00110100", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", "00111110", 
"00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001010", 
"01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", 
"01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", 
"10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10101111", "10110000", 
"10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", 
"10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000110", "11000111", 
"11001000", "11001001", "11001001", "11001010", "11001011", "11001100", "11001100", "11001101", "11001110", "11001111", "11001111", "11010000", "11010001", "11010010", "11010011", "11010011", "11010100", "11010101", "11010110", "11010111", 
"11011000", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", 
"11101010", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", 
"11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", 
"00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", 
"00100100", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00101111", "00110000", "00110001", "00110010", "00110010", "00110011", 
"00110100", "00110101", "00110110", "00110110", "00110111", "00111000", "00111000", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", 
"01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", 
"01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", 
"01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", 
"10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110000", "10110001", "10110001", 
"10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111100", 
"10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11001000", "11001000", "11001001", "11001010", 
"11001010", "11001011", "11001100", "11001101", "11001110", "11001110", "11001111", "11010000", "11010001", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010110", "11010111", "11011000", "11011001", "11011010", 
"11011011", "11011100", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", 
"11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", 
"00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", 
"00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100110", 
"00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101100", "00101101", "00101110", "00101111", "00110000", "00110000", "00110001", "00110010", "00110011", "00110100", "00110100", "00110101", "00110110", "00110111", 
"00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", 
"01000101", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", 
"01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", 
"01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", 
"10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", 
"10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111110", 
"10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001001", "11001010", "11001011", "11001100", "11001100", 
"11001101", "11001110", "11001111", "11010000", "11010000", "11010001", "11010010", "11010011", "11010100", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011010", "11011011", "11011100", "11011101", 
"11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", 
"11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", 
"00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", 
"00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101000", "00101001", "00101010", 
"00101011", "00101100", "00101101", "00101110", "00101110", "00101111", "00110000", "00110001", "00110010", "00110010", "00110011", "00110100", "00110101", "00110101", "00110110", "00110111", "00111000", "00111000", "00111001", "00111010", 
"00111011", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", 
"01000111", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", 
"01010010", "01010010", "01010011", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", 
"01011010", "10100111", "10100111", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", 
"10101100", "10101100", "10101101", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", 
"10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", 
"11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11001000", "11001000", "11001001", "11001010", "11001011", "11001011", "11001100", "11001101", "11001110", "11001110", "11001111", 
"11010000", "11010001", "11010010", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", 
"11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", 
"11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", 
"00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", 
"00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101010", "00101011", "00101100", "00101101", "00101110", 
"00101111", "00101111", "00110000", "00110001", "00110010", "00110011", "00110011", "00110100", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111100", "00111101", 
"00111110", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001010", 
"01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010011", 
"01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "01011000", 
"01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", 
"10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", 
"10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", 
"11000100", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001001", "11001010", "11001011", "11001100", "11001101", "11001101", "11001110", "11001111", "11010000", "11010001", "11010001", "11010010", 
"11010011", "11010100", "11010101", "11010110", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", 
"11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", 
"11111001", "11111010", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", 
"00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", 
"00100001", "00100010", "00100011", "00100100", "00100101", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110001", 
"00110010", "00110011", "00110100", "00110101", "00110101", "00110110", "00110111", "00111000", "00111000", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "00111111", "01000000", 
"01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", 
"01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", 
"01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "01011000", "01011000", "01011001", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", 
"10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000101", 
"11000110", "11000111", "11001000", "11001000", "11001001", "11001010", "11001011", "11001011", "11001100", "11001101", "11001110", "11001111", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010100", "11010101", 
"11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", 
"11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", 
"11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010001", 
"00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", 
"00100101", "00100110", "00100111", "00101000", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110011", "00110100", "00110101", 
"00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", 
"01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", 
"01001111", "01010000", "01010000", "01010001", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", 
"01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", 
"10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10101111", 
"10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", 
"10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", 
"11001001", "11001001", "11001010", "11001011", "11001100", "11001101", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011000", 
"11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11100111", "11101000", "11101001", "11101010", "11101011", 
"11101100", "11101101", "11101110", "11101111", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", 
"00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", 
"00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", 
"00101001", "00101010", "00101011", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110001", "00110010", "00110011", "00110100", "00110101", "00110101", "00110110", "00110111", "00111000", "00111000", 
"00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", 
"01000111", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", 
"01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", 
"10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", 
"10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111100", 
"10111101", "10111110", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11001000", "11001000", "11001001", "11001010", "11001011", 
"11001011", "11001100", "11001101", "11001110", "11001111", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", 
"11011101", "11011110", "11011111", "11100000", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", 
"11110000", "11110001", "11110010", "11110011", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", 
"00000101", "00000110", "00000111", "00001000", "00001001", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", 
"00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", 
"00101101", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110010", "00110011", "00110100", "00110101", "00110110", "00110110", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", 
"00111100", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", 
"01001001", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", 
"01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", 
"10101000", "10101000", "10101001", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", 
"10101010", "10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", 
"10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", 
"10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001010", "11001010", "11001011", "11001100", "11001101", "11001110", 
"11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011100", "11011101", "11011110", "11011111", 
"11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", 
"11110100", "11110101", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001001", 
"00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", 
"00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", 
"00110000", "00110001", "00110010", "00110011", "00110100", "00110100", "00110101", "00110110", "00110111", "00111000", "00111000", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", 
"01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001100", 
"01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", 
"01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "01010110", 
"01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", 
"10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", 
"10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000000", "11000001", 
"11000010", "11000010", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11001000", "11001000", "11001001", "11001010", "11001011", "11001100", "11001100", "11001101", "11001110", "11001111", "11010000", "11010000", 
"11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", 
"11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", 
"11111001", "11111010", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", 
"00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", 
"00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110010", "00110011", 
"00110100", "00110101", "00110110", "00110110", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", 
"01000011", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", 
"01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", 
"01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "01010110", "01010110", "01010111", "01010111", "01011000", 
"01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", 
"10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", 
"10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000011", 
"11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001010", "11001010", "11001011", "11001100", "11001101", "11001110", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", 
"11010101", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", 
"11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111010", "11111011", "11111100", 
"11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", 
"00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100010", "00100011", "00100100", "00100101", 
"00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110100", "00110101", "00110110", "00110111", 
"00111000", "00111000", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", 
"01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", 
"01010001", "01010010", "01010010", "01010011", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", 
"01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101101", 
"10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000101", "11000101", "11000110", 
"11000111", "11001000", "11001000", "11001001", "11001010", "11001011", "11001100", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", 
"11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11101000", "11101001", "11101010", "11101011", 
"11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", 
"00000001", "00000010", "00000011", "00000100", "00000101", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010101", "00010110", 
"00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101000", "00101001", 
"00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110110", "00110111", "00111000", "00111001", "00111010", "00111010", 
"00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", 
"01001001", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", 
"01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", 
"10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", 
"10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", 
"10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", 
"10111011", "10111100", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", 
"11001010", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011000", "11011001", "11011010", 
"11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101101", "11101110", "11101111", 
"11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111011", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", 
"00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", 
"00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101100", "00101101", 
"00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111000", "00111001", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", 
"00111110", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", 
"01001011", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", 
"01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", 
"10101010", "10101010", "10101011", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", 
"10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", 
"10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", 
"10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", "11001000", "11001000", "11001001", "11001010", "11001011", "11001100", 
"11001101", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", 
"11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11110000", "11110001", "11110010", "11110011", 
"11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000110", "00000111", "00001000", "00001001", 
"00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", 
"00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110000", "00110001", 
"00110010", "00110011", "00110100", "00110101", "00110110", "00110110", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "01000000", "01000000", "01000001", 
"01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001110", 
"01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", 
"01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "01010100", 
"01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", 
"10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", 
"10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111110", "10111111", 
"11000000", "11000000", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001010", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", 
"11010000", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", 
"11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", 
"11111000", "11111001", "11111010", "11111100", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000100", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", 
"00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", 
"00100100", "00100101", "00100110", "00100111", "00101000", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110011", "00110100", "00110101", 
"00110110", "00110111", "00111000", "00111000", "00111001", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000100", "01000100", 
"01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", 
"01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "01010100", "01010100", "01010101", "01010101", "01010110", 
"01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", 
"10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110100", 
"10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000001", 
"11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", "11001000", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", 
"11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100100", "11100101", "11100110", 
"11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111100", 
"11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001110", "00001111", "00010000", "00010001", "00010010", 
"00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", 
"00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110101", "00110110", "00110111", "00111000", "00111001", 
"00111010", "00111010", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", 
"01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", 
"01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", 
"10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", 
"01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", 
"10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", 
"10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", 
"11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010010", "11010011", "11010100", "11010101", 
"11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11101000", "11101001", "11101010", 
"11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111101", "11111110", "11111111", "00000000", 
"00000001", "00000010", "00000011", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010111", 
"00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", 
"00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111000", "00111001", "00111010", "00111011", "00111100", "00111100", 
"00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", 
"01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", 
"01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", 
"10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101100", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", 
"01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", 
"10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", 
"11001000", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", 
"11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101011", "11101100", "11101101", "11101110", 
"11101111", "11110000", "11110001", "11110010", "11110011", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000101", 
"00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", 
"00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100110", "00100111", "00101000", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", 
"00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", 
"01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", 
"01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", 
"01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101011", "10101100", 
"10101100", "10101100", "10101101", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", 
"01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101111", 
"10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", 
"10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001010", 
"11001011", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011000", "11011001", "11011010", "11011100", "11011101", 
"11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101101", "11101110", "11101111", "11110000", "11110001", "11110010", 
"11110011", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000011", "00000101", "00000110", "00000111", "00001000", "00001001", 
"00001010", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011111", "00100000", 
"00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110000", "00110001", "00110010", "00110011", 
"00110100", "00110101", "00110110", "00110111", "00111000", "00111000", "00111001", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", "01000011", 
"01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", 
"01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101101", "01010010", 
"01010011", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", 
"10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", 
"10110001", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", 
"10111101", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", "11001000", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", 
"11001110", "11001111", "11010000", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", 
"11100001", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101110", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110110", "11110111", 
"11111000", "11111001", "11111010", "11111011", "11111101", "11111110", "11111111", "00000000", "00000001", "00000010", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001011", "00001100", "00001101", "00001110", 
"00001111", "00010000", "00010001", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", 
"00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110100", "00110101", "00110110", "00110111", 
"00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", 
"01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", 
"01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", 
"10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101101", "10101110", "01010010", "01010010", "01010011", "01010011", "01010011", 
"01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", 
"10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", 
"10110011", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111111", "10111111", 
"11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001100", "11001101", "11001110", "11001111", "11010000", 
"11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", 
"11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101111", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110111", "11111000", "11111001", "11111010", "11111011", 
"11111100", "11111110", "11111111", "00000000", "00000001", "00000010", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010010", "00010011", 
"00010100", "00010101", "00010110", "00010111", "00011000", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", 
"00101010", "00101011", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111000", "00111001", "00111010", "00111011", 
"00111100", "00111101", "00111101", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", 
"01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", 
"01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", 
"10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101101", "10101110", "10101110", "01010001", "01010010", "01010010", "01010011", "01010011", "01010011", "01010100", "01010100", "01010101", 
"01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", 
"10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", 
"10110101", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", 
"11000011", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", 
"11010101", "11010101", "11010110", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11101000", "11101001", 
"11101010", "11101011", "11101100", "11101101", "11101110", "11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110111", "11111000", "11111001", "11111010", "11111011", "11111100", "11111110", "11111111", "00000000", 
"00000001", "00000010", "00000100", "00000101", "00000110", "00000111", "00001000", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00011000", 
"00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", 
"00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", 
"00111111", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", 
"01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", 
"01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", 
"10101100", "10101101", "10101101", "10101101", "10101110", "10101110", "10101111", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", 
"01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", 
"10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", 
"10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000101", 
"11000110", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", 
"11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101010", "11101011", "11101100", "11101101", 
"11101110", "11101111", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11111000", "11111001", "11111010", "11111011", "11111100", "11111110", "11111111", "00000000", "00000001", "00000010", "00000100", "00000101", 
"00000110", "00000111", "00001000", "00001010", "00001011", "00001100", "00001101", "00001110", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", 
"00011101", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", 
"00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "01000000", "01000001", "01000001", "01000010", 
"01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", "01001111", 
"01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", 
"10101110", "10101111", "10101111", "01010001", "01010001", "01010001", "01010010", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", 
"01010111", "01011000", "01011000", "01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", 
"10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", 
"11001001", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", 
"11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110010", 
"11110011", "11110100", "11110101", "11110110", "11111000", "11111001", "11111010", "11111011", "11111100", "11111110", "11111111", "00000000", "00000001", "00000010", "00000100", "00000101", "00000110", "00000111", "00001001", "00001010", 
"00001011", "00001100", "00001101", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011101", "00011110", "00011111", "00100000", "00100001", 
"00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110001", "00110010", "00110011", "00110100", "00110101", 
"00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", 
"01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", 
"01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", 
"10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101110", "10101111", "10101111", "10110000", "01010000", 
"01010000", "01010001", "01010001", "01010010", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", 
"01011001", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", 
"10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", 
"10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", 
"11001100", "11001101", "11001110", "11001111", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", 
"11100000", "11100001", "11100010", "11100011", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101100", "11101101", "11101110", "11101111", "11110000", "11110001", "11110011", "11110100", "11110101", "11110110", 
"11110111", "11111001", "11111010", "11111011", "11111100", "11111110", "11111111", "00000000", "00000001", "00000010", "00000100", "00000101", "00000110", "00000111", "00001001", "00001010", "00001011", "00001100", "00001101", "00001111", 
"00010000", "00010001", "00010010", "00010011", "00010101", "00010110", "00010111", "00011000", "00011001", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100100", "00100101", "00100110", 
"00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", 
"00111010", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001001", 
"01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", 
"01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", 
"10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "01010000", "01010000", "01010000", "01010001", "01010001", 
"01010010", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", 
"10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", 
"10111110", "10111111", "10111111", "11000000", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", 
"11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", 
"11100100", "11100101", "11100111", "11101000", "11101001", "11101010", "11101011", "11101101", "11101110", "11101111", "11110000", "11110001", "11110011", "11110100", "11110101", "11110110", "11110111", "11111001", "11111010", "11111011", 
"11111100", "11111110", "11111111", "00000000", "00000001", "00000010", "00000100", "00000101", "00000110", "00000111", "00001001", "00001010", "00001011", "00001100", "00001110", "00001111", "00010000", "00010001", "00010010", "00010100", 
"00010101", "00010110", "00010111", "00011000", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", 
"00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", 
"00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", 
"01001101", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", 
"01011000", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", 
"10101101", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10101111", "10110000", "10110000", "10110000", "01001111", "01010000", "01010000", "01010000", "01010001", "01010001", "01010001", "01010010", "01010010", 
"01010011", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", 
"10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110010", 
"10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "11000000", 
"11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", 
"11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11101000", 
"11101001", "11101010", "11101011", "11101100", "11101110", "11101111", "11110000", "11110001", "11110010", "11110100", "11110101", "11110110", "11110111", "11111001", "11111010", "11111011", "11111100", "11111110", "11111111", "00000000", 
"00000001", "00000011", "00000100", "00000101", "00000110", "00001000", "00001001", "00001010", "00001011", "00001101", "00001110", "00001111", "00010000", "00010001", "00010011", "00010100", "00010101", "00010110", "00010111", "00011001", 
"00011010", "00011011", "00011100", "00011101", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", 
"00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000001", 
"01000010", "01000010", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", 
"01001111", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101101", "10101110", "10101110", 
"10101111", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "01001111", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010011", 
"01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", 
"10101001", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110100", 
"10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000010", "11000010", 
"11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", 
"11010110", "11010111", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100011", "11100100", "11100101", "11100110", "11100111", "11101001", "11101010", "11101011", "11101100", 
"11101101", "11101111", "11110000", "11110001", "11110010", "11110011", "11110101", "11110110", "11110111", "11111000", "11111010", "11111011", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000101", 
"00000110", "00001000", "00001001", "00001010", "00001011", "00001101", "00001110", "00001111", "00010000", "00010010", "00010011", "00010100", "00010101", "00010110", "00011000", "00011001", "00011010", "00011011", "00011100", "00011110", 
"00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", 
"00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000100", "01000100", 
"01000101", "01000110", "01000111", "01000111", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", 
"01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", 
"10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10101111", "10110000", "10110000", 
"10110001", "10110001", "10110001", "01001110", "01001111", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010011", "01010100", "01010100", "01010101", 
"01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", 
"10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110110", 
"10110110", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000101", 
"11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", 
"11011010", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100100", "11100101", "11100110", "11100111", "11101000", "11101010", "11101011", "11101100", "11101101", "11101110", "11110000", "11110001", 
"11110010", "11110011", "11110101", "11110110", "11110111", "11111000", "11111010", "11111011", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000101", "00000110", "00001000", "00001001", "00001010", 
"00001011", "00001101", "00001110", "00001111", "00010001", "00010010", "00010011", "00010100", "00010101", "00010111", "00011000", "00011001", "00011010", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100011", 
"00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110110", "00110111", 
"00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", 
"01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", 
"01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", 
"10101011", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "01001110", 
"01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010101", "01010110", 
"01010110", "01010111", "01010111", "01011000", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", 
"10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", 
"11001010", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", 
"11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100110", "11100111", "11101000", "11101001", "11101011", "11101100", "11101101", "11101110", "11101111", "11110001", "11110010", "11110011", "11110101", "11110110", 
"11110111", "11111000", "11111010", "11111011", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000101", "00000110", "00001000", "00001001", "00001010", "00001100", "00001101", "00001110", "00001111", 
"00010001", "00010010", "00010011", "00010100", "00010110", "00010111", "00011000", "00011001", "00011011", "00011100", "00011101", "00011110", "00011111", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", 
"00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", 
"00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001011", "01001011", 
"01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", 
"01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", 
"10101101", "10101101", "10101110", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110010", "01001101", "01001110", "01001110", "01001110", "01001111", 
"01001111", "01010000", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", 
"01011000", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", 
"10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111011", 
"10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", 
"11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100001", "11100010", 
"11100011", "11100100", "11100101", "11100111", "11101000", "11101001", "11101010", "11101100", "11101101", "11101110", "11101111", "11110001", "11110010", "11110011", "11110100", "11110110", "11110111", "11111000", "11111010", "11111011", 
"11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000101", "00000111", "00001000", "00001001", "00001010", "00001100", "00001101", "00001110", "00010000", "00010001", "00010010", "00010011", "00010101", 
"00010110", "00010111", "00011000", "00011010", "00011011", "00011100", "00011101", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", 
"00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "00111111", 
"01000000", "01000001", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000111", "01000111", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", 
"01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", 
"10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "01001101", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01001111", "01010000", 
"01010000", "01010001", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011000", 
"01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101111", "10101111", 
"10110000", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111100", "10111100", "10111101", 
"10111110", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", 
"11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100011", "11100100", "11100101", "11100110", 
"11101000", "11101001", "11101010", "11101011", "11101101", "11101110", "11101111", "11110000", "11110010", "11110011", "11110100", "11110110", "11110111", "11111000", "11111001", "11111011", "11111100", "11111101", "11111111", "00000000", 
"00000001", "00000011", "00000100", "00000101", "00000111", "00001000", "00001001", "00001011", "00001100", "00001101", "00001110", "00010000", "00010001", "00010010", "00010100", "00010101", "00010110", "00010111", "00011001", "00011010", 
"00011011", "00011100", "00011110", "00011111", "00100000", "00100001", "00100010", "00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", 
"00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000010", "01000011", 
"01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", 
"01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", 
"10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10101111", "10110000", "10110000", "10110001", 
"10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110011", "01001100", "01001101", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", 
"01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", 
"10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", 
"10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", 
"11000001", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", 
"11010100", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011110", "11011111", "11100000", "11100001", "11100010", "11100100", "11100101", "11100110", "11100111", "11101001", "11101010", "11101011", 
"11101100", "11101110", "11101111", "11110000", "11110010", "11110011", "11110100", "11110101", "11110111", "11111000", "11111001", "11111011", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000101", 
"00000111", "00001000", "00001001", "00001011", "00001100", "00001101", "00001111", "00010000", "00010001", "00010011", "00010100", "00010101", "00010110", "00011000", "00011001", "00011010", "00011011", "00011101", "00011110", "00011111", 
"00100000", "00100010", "00100011", "00100100", "00100101", "00100110", "00100111", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", 
"00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", 
"01001000", "01001000", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", 
"01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", 
"10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110010", "10110011", 
"10110011", "10110100", "10110100", "01001100", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", 
"01010011", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", 
"10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", 
"10110100", "10110101", "10110101", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000011", 
"11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", 
"11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11100000", "11100001", "11100010", "11100011", "11100101", "11100110", "11100111", "11101000", "11101010", "11101011", "11101100", "11101101", "11101111", "11110000", 
"11110001", "11110011", "11110100", "11110101", "11110111", "11111000", "11111001", "11111011", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000101", "00000111", "00001000", "00001001", "00001011", 
"00001100", "00001101", "00001111", "00010000", "00010001", "00010011", "00010100", "00010101", "00010111", "00011000", "00011001", "00011010", "00011100", "00011101", "00011110", "00011111", "00100001", "00100010", "00100011", "00100100", 
"00100101", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", 
"00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000111", "01000111", "01001000", "01001001", "01001010", "01001010", 
"01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", 
"01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", 
"10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110100", "01001011", 
"01001100", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010011", 
"01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", 
"10101010", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110110", 
"10110110", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000110", 
"11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011011", "11011100", 
"11011101", "11011110", "11011111", "11100001", "11100010", "11100011", "11100100", "11100110", "11100111", "11101000", "11101001", "11101011", "11101100", "11101101", "11101111", "11110000", "11110001", "11110011", "11110100", "11110101", 
"11110111", "11111000", "11111001", "11111011", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000101", "00000111", "00001000", "00001010", "00001011", "00001100", "00001110", "00001111", "00010000", 
"00010010", "00010011", "00010100", "00010110", "00010111", "00011000", "00011001", "00011011", "00011100", "00011101", "00011110", "00100000", "00100001", "00100010", "00100011", "00100101", "00100110", "00100111", "00101000", "00101001", 
"00101010", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", 
"00111111", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", 
"01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101110", "10101111", 
"10101111", "10110000", "10110000", "10110001", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "01001011", "01001011", "01001011", "01001100", "01001100", 
"01001101", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", 
"01010101", "01010110", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", 
"10101011", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", 
"11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011101", "11011110", "11011111", "11100000", 
"11100010", "11100011", "11100100", "11100101", "11100111", "11101000", "11101001", "11101010", "11101100", "11101101", "11101110", "11110000", "11110001", "11110010", "11110100", "11110101", "11110110", "11111000", "11111001", "11111011", 
"11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000110", "00000111", "00001000", "00001010", "00001011", "00001100", "00001110", "00001111", "00010000", "00010010", "00010011", "00010100", "00010110", 
"00010111", "00011000", "00011010", "00011011", "00011100", "00011110", "00011111", "00100000", "00100001", "00100011", "00100100", "00100101", "00100110", "00100111", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", 
"00101111", "00110000", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000001", "01000010", 
"01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", "01010001", 
"01010010", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", 
"10101001", "10101001", "10101010", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", 
"10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110100", "10110101", "10110101", "10110101", "01001010", "01001011", "01001011", "01001011", "01001100", "01001100", "01001100", "01001101", "01001101", 
"01001110", "01001110", "01001111", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", 
"01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101101", 
"10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", "10111011", 
"10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", 
"11001110", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011001", "11011010", "11011011", "11011100", "11011101", "11011111", "11100000", "11100001", "11100010", "11100100", "11100101", 
"11100110", "11101000", "11101001", "11101010", "11101100", "11101101", "11101110", "11110000", "11110001", "11110010", "11110100", "11110101", "11110110", "11111000", "11111001", "11111010", "11111100", "11111101", "11111111", "00000000", 
"00000001", "00000011", "00000100", "00000110", "00000111", "00001000", "00001010", "00001011", "00001100", "00001110", "00001111", "00010001", "00010010", "00010011", "00010101", "00010110", "00010111", "00011001", "00011010", "00011011", 
"00011101", "00011110", "00011111", "00100000", "00100010", "00100011", "00100100", "00100101", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", 
"00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", 
"01000111", "01001000", "01001000", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", 
"01010100", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", 
"10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110010", "10110011", "10110011", 
"10110100", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "01001010", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001110", 
"01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", 
"01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101111", 
"10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111101", 
"10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", 
"11010010", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011011", "11011100", "11011101", "11011110", "11100000", "11100001", "11100010", "11100011", "11100101", "11100110", "11100111", "11101001", "11101010", 
"11101011", "11101101", "11101110", "11101111", "11110001", "11110010", "11110100", "11110101", "11110110", "11111000", "11111001", "11111010", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000110", 
"00000111", "00001000", "00001010", "00001011", "00001101", "00001110", "00001111", "00010001", "00010010", "00010100", "00010101", "00010110", "00011000", "00011001", "00011010", "00011100", "00011101", "00011110", "00011111", "00100001", 
"00100010", "00100011", "00100100", "00100110", "00100111", "00101000", "00101001", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110100", "00110101", "00110110", "00110111", "00111000", 
"00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001010", 
"01001010", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010110", "01010110", "01010111", 
"01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101100", "10101101", 
"10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110101", 
"10110110", "10110110", "10110111", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", 
"01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", 
"01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", 
"10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000000", 
"11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", 
"11010111", "11011000", "11011001", "11011010", "11011100", "11011101", "11011110", "11011111", "11100001", "11100010", "11100011", "11100100", "11100110", "11100111", "11101000", "11101010", "11101011", "11101100", "11101110", "11101111", 
"11110001", "11110010", "11110011", "11110101", "11110110", "11111000", "11111001", "11111010", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000110", "00000111", "00001001", "00001010", "00001011", 
"00001101", "00001110", "00010000", "00010001", "00010010", "00010100", "00010101", "00010110", "00011000", "00011001", "00011011", "00011100", "00011101", "00011110", "00100000", "00100001", "00100010", "00100100", "00100101", "00100110", 
"00100111", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", 
"00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001100", "01001100", "01001101", 
"01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", 
"10110000", "10110000", "10110001", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110110", "10110111", "10110111", "01001001", 
"01001001", "01001001", "01001010", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01001111", "01010000", "01010000", "01010001", 
"01010001", "01010010", "01010010", "01010011", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", 
"10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", 
"10110100", "10110100", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", 
"11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011001", "11011010", 
"11011011", "11011100", "11011110", "11011111", "11100000", "11100010", "11100011", "11100100", "11100101", "11100111", "11101000", "11101010", "11101011", "11101100", "11101110", "11101111", "11110000", "11110010", "11110011", "11110101", 
"11110110", "11110111", "11111001", "11111010", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000110", "00000111", "00001001", "00001010", "00001011", "00001101", "00001110", "00010000", "00010001", 
"00010011", "00010100", "00010101", "00010111", "00011000", "00011001", "00011011", "00011100", "00011101", "00011111", "00100000", "00100001", "00100011", "00100100", "00100101", "00100111", "00101000", "00101001", "00101010", "00101011", 
"00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", 
"01000010", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", 
"01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", 
"10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", 
"10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110110", "10110111", "10110111", "10111000", "01001000", "01001000", "01001001", "01001001", "01001010", 
"01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", 
"01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", 
"10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110101", "10110101", 
"10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", 
"11001000", "11001001", "11001010", "11001011", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010101", "11010110", "11010111", "11011000", "11011001", "11011011", "11011100", "11011101", "11011111", 
"11100000", "11100001", "11100011", "11100100", "11100101", "11100111", "11101000", "11101001", "11101011", "11101100", "11101101", "11101111", "11110000", "11110010", "11110011", "11110101", "11110110", "11110111", "11111001", "11111010", 
"11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000110", "00000111", "00001001", "00001010", "00001100", "00001101", "00001111", "00010000", "00010001", "00010011", "00010100", "00010110", "00010111", 
"00011000", "00011010", "00011011", "00011100", "00011110", "00011111", "00100000", "00100010", "00100011", "00100100", "00100110", "00100111", "00101000", "00101001", "00101011", "00101100", "00101101", "00101110", "00101111", "00110001", 
"00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", 
"01000110", "01000110", "01000111", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", 
"01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", 
"10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110011", "10110100", 
"10110100", "10110101", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10110111", "10111000", "10111000", "01000111", "01001000", "01001000", "01001001", "01001001", "01001001", "01001010", "01001010", "01001011", 
"01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", 
"01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", 
"10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", 
"11001100", "11001101", "11001110", "11001111", "11010001", "11010010", "11010011", "11010100", "11010101", "11010111", "11011000", "11011001", "11011010", "11011100", "11011101", "11011110", "11100000", "11100001", "11100010", "11100100", 
"11100101", "11100110", "11101000", "11101001", "11101010", "11101100", "11101101", "11101111", "11110000", "11110001", "11110011", "11110100", "11110110", "11110111", "11111001", "11111010", "11111100", "11111101", "11111111", "00000000", 
"00000001", "00000011", "00000100", "00000110", "00000111", "00001001", "00001010", "00001100", "00001101", "00001111", "00010000", "00010010", "00010011", "00010100", "00010110", "00010111", "00011001", "00011010", "00011011", "00011101", 
"00011110", "00011111", "00100001", "00100010", "00100011", "00100101", "00100110", "00100111", "00101001", "00101010", "00101011", "00101100", "00101101", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110110", 
"00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", 
"01001001", "01001010", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", 
"01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", 
"10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", 
"10110110", "10110111", "10110111", "10111000", "10111000", "10111000", "10111001", "01000111", "01000111", "01001000", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001010", "01001011", "01001011", "01001100", 
"01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", 
"01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", 
"10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", "10111011", 
"10111100", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001100", "11001101", "11001110", "11001111", 
"11010000", "11010001", "11010011", "11010100", "11010101", "11010110", "11010111", "11011001", "11011010", "11011011", "11011101", "11011110", "11011111", "11100001", "11100010", "11100011", "11100101", "11100110", "11100111", "11101001", 
"11101010", "11101100", "11101101", "11101110", "11110000", "11110001", "11110011", "11110100", "11110110", "11110111", "11111001", "11111010", "11111100", "11111101", "11111111", "00000000", "00000001", "00000011", "00000100", "00000110", 
"00000111", "00001001", "00001010", "00001100", "00001101", "00001111", "00010000", "00010010", "00010011", "00010101", "00010110", "00010111", "00011001", "00011010", "00011100", "00011101", "00011110", "00100000", "00100001", "00100011", 
"00100100", "00100101", "00100110", "00101000", "00101001", "00101010", "00101100", "00101101", "00101110", "00101111", "00110000", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", 
"00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001011", "01001100", "01001100", 
"01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", 
"10110000", "10110001", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10110111", "10111000", "10111000", 
"10111001", "10111001", "10111001", "01000110", "01000111", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001011", "01001100", "01001100", "01001101", 
"01001101", "01001110", "01001110", "01001111", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", 
"01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", 
"10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", 
"10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11010000", "11010001", "11010010", "11010011", 
"11010100", "11010110", "11010111", "11011000", "11011010", "11011011", "11011100", "11011101", "11011111", "11100000", "11100010", "11100011", "11100100", "11100110", "11100111", "11101001", "11101010", "11101011", "11101101", "11101110", 
"11110000", "11110001", "11110011", "11110100", "11110110", "11110111", "11111001", "11111010", "11111100", "11111101", "11111111", "00000000", "00000010", "00000011", "00000101", "00000110", "00001000", "00001001", "00001011", "00001100", 
"00001110", "00001111", "00010000", "00010010", "00010011", "00010101", "00010110", "00011000", "00011001", "00011011", "00011100", "00011101", "00011111", "00100000", "00100010", "00100011", "00100100", "00100110", "00100111", "00101000", 
"00101001", "00101011", "00101100", "00101101", "00101110", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", 
"01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", 
"01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", 
"10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", 
"10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "01000110", 
"01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", 
"01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", 
"01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10101111", "10110000", 
"10110001", "10110010", "10110010", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", 
"11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010010", "11010011", "11010100", "11010101", "11010111", "11011000", 
"11011001", "11011010", "11011100", "11011101", "11011110", "11100000", "11100001", "11100011", "11100100", "11100101", "11100111", "11101000", "11101010", "11101011", "11101101", "11101110", "11110000", "11110001", "11110010", "11110100", 
"11110101", "11110111", "11111000", "11111010", "11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000110", "00001000", "00001001", "00001011", "00001100", "00001110", "00001111", "00010001", "00010010", 
"00010100", "00010101", "00010111", "00011000", "00011001", "00011011", "00011100", "00011110", "00011111", "00100001", "00100010", "00100011", "00100101", "00100110", "00100111", "00101001", "00101010", "00101011", "00101100", "00101110", 
"00101111", "00110000", "00110001", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000010", "01000011", 
"01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010011", "01010011", 
"01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", 
"10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110100", 
"10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111001", "10111010", "10111010", "10111011", "01000101", "01000101", "01000110", "01000110", "01000111", 
"01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", 
"01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110010", 
"10110011", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000101", 
"11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001111", "11010000", "11010001", "11010010", "11010100", "11010101", "11010110", "11010111", "11011001", "11011010", "11011011", "11011101", 
"11011110", "11011111", "11100001", "11100010", "11100100", "11100101", "11100111", "11101000", "11101001", "11101011", "11101100", "11101110", "11101111", "11110001", "11110010", "11110100", "11110101", "11110111", "11111000", "11111010", 
"11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000110", "00001000", "00001001", "00001011", "00001100", "00001110", "00001111", "00010001", "00010010", "00010100", "00010101", "00010111", "00011000", 
"00011010", "00011011", "00011101", "00011110", "00100000", "00100001", "00100010", "00100100", "00100101", "00100110", "00101000", "00101001", "00101010", "00101100", "00101101", "00101110", "00101111", "00110001", "00110010", "00110011", 
"00110100", "00110101", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", 
"01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010110", 
"01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", 
"10101110", "10101111", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110101", "10110110", "10110110", "10110111", 
"10110111", "10111000", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111010", "10111011", "10111011", "01000101", "01000101", "01000101", "01000110", "01000110", "01000110", "01000111", "01000111", "01001000", 
"01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", 
"01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", 
"10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", 
"10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", 
"11001001", "11001011", "11001100", "11001101", "11001110", "11001111", "11010001", "11010010", "11010011", "11010100", "11010110", "11010111", "11011000", "11011010", "11011011", "11011100", "11011110", "11011111", "11100000", "11100010", 
"11100011", "11100101", "11100110", "11101000", "11101001", "11101011", "11101100", "11101110", "11101111", "11110001", "11110010", "11110100", "11110101", "11110111", "11111000", "11111010", "11111011", "11111101", "11111110", "00000000", 
"00000010", "00000011", "00000101", "00000110", "00001000", "00001001", "00001011", "00001100", "00001110", "00010000", "00010001", "00010011", "00010100", "00010110", "00010111", "00011001", "00011010", "00011100", "00011101", "00011110", 
"00100000", "00100001", "00100011", "00100100", "00100101", "00100111", "00101000", "00101001", "00101011", "00101100", "00101101", "00101111", "00110000", "00110001", "00110010", "00110100", "00110101", "00110110", "00110111", "00111000", 
"00111001", "00111010", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", 
"01001100", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", 
"10110001", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", 
"10111001", "10111010", "10111010", "10111011", "10111011", "10111011", "10111100", "01000100", "01000100", "01000101", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01000111", "01001000", "01001000", "01001001", 
"01001001", "01001010", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", 
"01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", 
"10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110111", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", 
"11001110", "11001111", "11010000", "11010001", "11010011", "11010100", "11010101", "11010111", "11011000", "11011001", "11011011", "11011100", "11011101", "11011111", "11100000", "11100010", "11100011", "11100100", "11100110", "11100111", 
"11101001", "11101010", "11101100", "11101101", "11101111", "11110000", "11110010", "11110100", "11110101", "11110111", "11111000", "11111010", "11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000110", 
"00001000", "00001001", "00001011", "00001101", "00001110", "00010000", "00010001", "00010011", "00010100", "00010110", "00010111", "00011001", "00011010", "00011100", "00011101", "00011111", "00100000", "00100010", "00100011", "00100100", 
"00100110", "00100111", "00101001", "00101010", "00101011", "00101101", "00101110", "00101111", "00110000", "00110010", "00110011", "00110100", "00110101", "00110110", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", 
"00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001110", "01001111", "01001111", 
"01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", 
"10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", 
"10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111010", "10111011", "10111011", 
"10111100", "10111100", "10111100", "01000011", "01000100", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001001", "01001010", 
"01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", 
"01010100", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", 
"10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", 
"10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001010", "11001011", "11001100", "11001101", "11001110", "11010000", "11010001", 
"11010010", "11010011", "11010101", "11010110", "11010111", "11011001", "11011010", "11011100", "11011101", "11011110", "11100000", "11100001", "11100011", "11100100", "11100110", "11100111", "11101001", "11101010", "11101100", "11101101", 
"11101111", "11110000", "11110010", "11110011", "11110101", "11110111", "11111000", "11111010", "11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000110", "00001000", "00001010", "00001011", "00001101", 
"00001110", "00010000", "00010010", "00010011", "00010101", "00010110", "00011000", "00011001", "00011011", "00011100", "00011110", "00011111", "00100001", "00100010", "00100100", "00100101", "00100110", "00101000", "00101001", "00101010", 
"00101100", "00101101", "00101110", "00110000", "00110001", "00110010", "00110011", "00110101", "00110110", "00110111", "00111000", "00111001", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", 
"01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", 
"01010100", "01010100", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101011", 
"10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", 
"10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "01000011", 
"01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", 
"01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", 
"01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", 
"10101110", "10101111", "10101111", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", 
"10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000111", "11001000", "11001001", "11001010", "11001011", "11001101", "11001110", "11001111", "11010000", "11010010", "11010011", "11010100", "11010110", 
"11010111", "11011000", "11011010", "11011011", "11011100", "11011110", "11011111", "11100001", "11100010", "11100100", "11100101", "11100111", "11101000", "11101010", "11101011", "11101101", "11101110", "11110000", "11110010", "11110011", 
"11110101", "11110110", "11111000", "11111010", "11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000111", "00001000", "00001010", "00001011", "00001101", "00001111", "00010000", "00010010", "00010011", 
"00010101", "00010110", "00011000", "00011010", "00011011", "00011101", "00011110", "00100000", "00100001", "00100010", "00100100", "00100101", "00100111", "00101000", "00101010", "00101011", "00101100", "00101110", "00101111", "00110000", 
"00110001", "00110011", "00110100", "00110101", "00110110", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000110", 
"01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", 
"01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", 
"10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10110111", 
"10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111100", "10111101", "10111101", "10111110", "01000010", "01000010", "01000011", "01000011", "01000100", 
"01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", 
"01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", 
"01010111", "01011000", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10101111", 
"10110000", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000001", "11000010", 
"11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001010", "11001011", "11001100", "11001101", "11001111", "11010000", "11010001", "11010010", "11010100", "11010101", "11010110", "11011000", "11011001", "11011011", 
"11011100", "11011110", "11011111", "11100000", "11100010", "11100011", "11100101", "11100110", "11101000", "11101010", "11101011", "11101101", "11101110", "11110000", "11110001", "11110011", "11110101", "11110110", "11111000", "11111001", 
"11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000111", "00001000", "00001010", "00001011", "00001101", "00001111", "00010000", "00010010", "00010100", "00010101", "00010111", "00011000", "00011010", 
"00011011", "00011101", "00011110", "00100000", "00100001", "00100011", "00100100", "00100110", "00100111", "00101001", "00101010", "00101011", "00101101", "00101110", "00101111", "00110001", "00110010", "00110011", "00110101", "00110110", 
"00110111", "00111000", "00111001", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", 
"01001100", "01001100", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", 
"10110001", "10110010", "10110010", "10110011", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111000", "10111001", "10111001", "10111010", 
"10111010", "10111011", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111101", "10111110", "10111110", "01000001", "01000010", "01000010", "01000011", "01000011", "01000011", "01000100", "01000100", "01000101", 
"01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001101", 
"01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", 
"01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", 
"10110011", "10110100", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", 
"11000111", "11001000", "11001001", "11001010", "11001011", "11001101", "11001110", "11001111", "11010001", "11010010", "11010011", "11010101", "11010110", "11010111", "11011001", "11011010", "11011100", "11011101", "11011111", "11100000", 
"11100010", "11100011", "11100101", "11100110", "11101000", "11101001", "11101011", "11101100", "11101110", "11110000", "11110001", "11110011", "11110101", "11110110", "11111000", "11111001", "11111011", "11111101", "11111110", "00000000", 
"00000010", "00000011", "00000101", "00000111", "00001000", "00001010", "00001100", "00001101", "00001111", "00010001", "00010010", "00010100", "00010101", "00010111", "00011001", "00011010", "00011100", "00011101", "00011111", "00100000", 
"00100010", "00100011", "00100101", "00100110", "00101000", "00101001", "00101011", "00101100", "00101101", "00101111", "00110000", "00110001", "00110011", "00110100", "00110101", "00110110", "00111000", "00111001", "00111010", "00111011", 
"00111100", "00111101", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", 
"01001111", "01010000", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", 
"10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", 
"10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", 
"10111100", "10111101", "10111101", "10111110", "10111110", "10111110", "10111111", "01000001", "01000001", "01000010", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000100", "01000101", "01000101", "01000110", 
"01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", 
"01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", 
"10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110100", "10110101", 
"10110110", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001010", 
"11001011", "11001100", "11001101", "11001111", "11010000", "11010001", "11010011", "11010100", "11010101", "11010111", "11011000", "11011010", "11011011", "11011101", "11011110", "11100000", "11100001", "11100011", "11100100", "11100110", 
"11100111", "11101001", "11101011", "11101100", "11101110", "11101111", "11110001", "11110011", "11110100", "11110110", "11111000", "11111001", "11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000111", 
"00001000", "00001010", "00001100", "00001101", "00001111", "00010001", "00010010", "00010100", "00010110", "00010111", "00011001", "00011010", "00011100", "00011110", "00011111", "00100001", "00100010", "00100100", "00100101", "00100111", 
"00101000", "00101010", "00101011", "00101100", "00101110", "00101111", "00110001", "00110010", "00110011", "00110100", "00110110", "00110111", "00111000", "00111001", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", 
"01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010010", "01010010", 
"01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", 
"10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", 
"10110110", "10110111", "10110111", "10111000", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111101", "10111110", "10111110", 
"10111111", "10111111", "10111111", "01000000", "01000001", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000101", "01000110", "01000110", "01000111", 
"01000111", "01001000", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", 
"01010001", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", 
"10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", 
"10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000111", "11001000", "11001001", "11001010", "11001100", "11001101", "11001110", 
"11001111", "11010001", "11010010", "11010100", "11010101", "11010110", "11011000", "11011001", "11011011", "11011100", "11011110", "11011111", "11100001", "11100010", "11100100", "11100110", "11100111", "11101001", "11101010", "11101100", 
"11101110", "11101111", "11110001", "11110011", "11110100", "11110110", "11111000", "11111001", "11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000111", "00001001", "00001010", "00001100", "00001110", 
"00001111", "00010001", "00010011", "00010100", "00010110", "00011000", "00011001", "00011011", "00011100", "00011110", "00100000", "00100001", "00100011", "00100100", "00100110", "00100111", "00101001", "00101010", "00101100", "00101101", 
"00101110", "00110000", "00110001", "00110010", "00110100", "00110101", "00110110", "00111000", "00111001", "00111010", "00111011", "00111100", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", 
"01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010101", "01010101", "01010110", 
"01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101110", 
"10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", 
"10111001", "10111001", "10111010", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "10111111", "11000000", "11000000", "01000000", 
"01000000", "01000000", "01000001", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000110", "01000111", "01000111", "01001000", 
"01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", 
"01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", 
"10101011", "10101011", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", 
"10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000100", "11000101", "11000110", "11000111", "11001000", "11001010", "11001011", "11001100", "11001110", "11001111", "11010000", "11010010", "11010011", 
"11010100", "11010110", "11010111", "11011001", "11011010", "11011100", "11011101", "11011111", "11100000", "11100010", "11100100", "11100101", "11100111", "11101000", "11101010", "11101100", "11101101", "11101111", "11110001", "11110010", 
"11110100", "11110110", "11110111", "11111001", "11111011", "11111101", "11111110", "00000000", "00000010", "00000011", "00000101", "00000111", "00001001", "00001010", "00001100", "00001110", "00010000", "00010001", "00010011", "00010101", 
"00010110", "00011000", "00011010", "00011011", "00011101", "00011110", "00100000", "00100010", "00100011", "00100101", "00100110", "00101000", "00101001", "00101011", "00101100", "00101101", "00101111", "00110000", "00110010", "00110011", 
"00110100", "00110110", "00110111", "00111000", "00111001", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", 
"01001011", "01001100", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", 
"10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", 
"10111011", "10111100", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000000", "11000001", "00111111", "00111111", "01000000", "01000000", "01000000", 
"01000001", "01000001", "01000010", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001000", "01001001", 
"01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010011", 
"01010100", "01010100", "01010101", "01010110", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101100", "10101100", 
"10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", 
"11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000111", "11001000", "11001001", "11001010", "11001100", "11001101", "11001110", "11010000", "11010001", "11010011", "11010100", "11010101", "11010111", "11011000", 
"11011010", "11011011", "11011101", "11011110", "11100000", "11100010", "11100011", "11100101", "11100110", "11101000", "11101010", "11101011", "11101101", "11101111", "11110000", "11110010", "11110100", "11110110", "11110111", "11111001", 
"11111011", "11111101", "11111110", "00000000", "00000010", "00000100", "00000101", "00000111", "00001001", "00001011", "00001100", "00001110", "00010000", "00010001", "00010011", "00010101", "00010111", "00011000", "00011010", "00011100", 
"00011101", "00011111", "00100000", "00100010", "00100100", "00100101", "00100111", "00101000", "00101010", "00101011", "00101101", "00101110", "00101111", "00110001", "00110010", "00110100", "00110101", "00110110", "00111000", "00111001", 
"00111010", "00111011", "00111100", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", 
"01001111", "01010000", "01010000", "01010001", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", 
"10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", 
"10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", 
"10111101", "10111110", "10111110", "10111111", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000001", "00111110", "00111111", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000001", 
"01000010", "01000010", "01000011", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", 
"01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", 
"01010110", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101111", 
"10110000", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", 
"11000100", "11000101", "11000110", "11000111", "11001000", "11001010", "11001011", "11001100", "11001110", "11001111", "11010001", "11010010", "11010011", "11010101", "11010110", "11011000", "11011001", "11011011", "11011100", "11011110", 
"11100000", "11100001", "11100011", "11100100", "11100110", "11101000", "11101001", "11101011", "11101101", "11101111", "11110000", "11110010", "11110100", "11110101", "11110111", "11111001", "11111011", "11111100", "11111110", "00000000", 
"00000010", "00000100", "00000101", "00000111", "00001001", "00001011", "00001100", "00001110", "00010000", "00010010", "00010011", "00010101", "00010111", "00011001", "00011010", "00011100", "00011110", "00011111", "00100001", "00100010", 
"00100100", "00100110", "00100111", "00101001", "00101010", "00101100", "00101101", "00101111", "00110000", "00110001", "00110011", "00110100", "00110110", "00110111", "00111000", "00111001", "00111011", "00111100", "00111101", "00111110", 
"01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", 
"01010011", "01010100", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", 
"10101100", "10101101", "10101101", "10101110", "10101111", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", 
"10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "10111111", 
"11000000", "11000000", "11000001", "11000001", "11000001", "11000010", "11000010", "00111110", "00111110", "00111110", "00111111", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000001", "01000010", "01000010", 
"01000011", "01000011", "01000100", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", 
"01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010111", 
"01010111", "01011000", "01011001", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101111", "10110000", "10110000", "10110001", 
"10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000010", "11000011", "11000100", "11000101", "11000111", 
"11001000", "11001001", "11001010", "11001100", "11001101", "11001111", "11010000", "11010001", "11010011", "11010100", "11010110", "11010111", "11011001", "11011010", "11011100", "11011110", "11011111", "11100001", "11100010", "11100100", 
"11100110", "11100111", "11101001", "11101011", "11101101", "11101110", "11110000", "11110010", "11110100", "11110101", "11110111", "11111001", "11111011", "11111100", "11111110", "00000000", "00000010", "00000100", "00000101", "00000111", 
"00001001", "00001011", "00001101", "00001110", "00010000", "00010010", "00010100", "00010101", "00010111", "00011001", "00011011", "00011100", "00011110", "00100000", "00100001", "00100011", "00100100", "00100110", "00101000", "00101001", 
"00101011", "00101100", "00101110", "00101111", "00110001", "00110010", "00110011", "00110101", "00110110", "00110111", "00111001", "00111010", "00111011", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000100", 
"01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010110", 
"01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", 
"10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", 
"10111010", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000000", "11000001", "11000001", "11000010", 
"11000010", "11000010", "11000011", "00111101", "00111101", "00111110", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000010", "01000011", "01000011", 
"01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", 
"01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", 
"01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", 
"10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000101", "11000110", "11000111", "11001001", "11001010", "11001011", 
"11001101", "11001110", "11001111", "11010001", "11010010", "11010100", "11010101", "11010111", "11011000", "11011010", "11011100", "11011101", "11011111", "11100000", "11100010", "11100100", "11100101", "11100111", "11101001", "11101011", 
"11101100", "11101110", "11110000", "11110010", "11110011", "11110101", "11110111", "11111001", "11111011", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00000111", "00001001", "00001011", "00001101", "00001111", 
"00010000", "00010010", "00010100", "00010110", "00011000", "00011001", "00011011", "00011101", "00011110", "00100000", "00100010", "00100011", "00100101", "00100111", "00101000", "00101010", "00101011", "00101101", "00101110", "00110000", 
"00110001", "00110011", "00110100", "00110101", "00110111", "00111000", "00111001", "00111011", "00111100", "00111101", "00111110", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001001", 
"01001010", "01001011", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", 
"01011010", "10100111", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", 
"10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", 
"10111100", "10111101", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000011", "00111100", 
"00111101", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000011", "01000100", "01000100", 
"01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", 
"01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011001", "01011010", "10100111", 
"10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", 
"10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000010", "11000011", "11000100", "11000101", "11000111", "11001000", "11001001", "11001011", "11001100", "11001101", "11001111", "11010000", 
"11010010", "11010011", "11010101", "11010110", "11011000", "11011001", "11011011", "11011101", "11011110", "11100000", "11100010", "11100011", "11100101", "11100111", "11101000", "11101010", "11101100", "11101110", "11110000", "11110001", 
"11110011", "11110101", "11110111", "11111001", "11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00000111", "00001001", "00001011", "00001101", "00001111", "00010001", "00010010", "00010100", "00010110", 
"00011000", "00011010", "00011011", "00011101", "00011111", "00100000", "00100010", "00100100", "00100101", "00100111", "00101001", "00101010", "00101100", "00101101", "00101111", "00110000", "00110010", "00110011", "00110101", "00110110", 
"00110111", "00111001", "00111010", "00111011", "00111101", "00111110", "00111111", "01000000", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", 
"01001110", "01001111", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", 
"10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110101", 
"10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", 
"10111111", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000011", "11000100", "11000100", "00111100", "00111100", "00111100", "00111101", "00111101", 
"00111101", "00111110", "00111110", "00111111", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", 
"01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", 
"01010000", "01010001", "01010010", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", 
"10101010", "10101010", "10101011", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", 
"10111100", "10111101", "10111110", "11000000", "11000001", "11000010", "11000011", "11000101", "11000110", "11000111", "11001001", "11001010", "11001011", "11001101", "11001110", "11010000", "11010001", "11010011", "11010100", "11010110", 
"11010111", "11011001", "11011011", "11011100", "11011110", "11100000", "11100001", "11100011", "11100101", "11100110", "11101000", "11101010", "11101100", "11101110", "11101111", "11110001", "11110011", "11110101", "11110111", "11111001", 
"11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00001000", "00001001", "00001011", "00001101", "00001111", "00010001", "00010011", "00010101", "00010110", "00011000", "00011010", "00011100", "00011101", 
"00011111", "00100001", "00100011", "00100100", "00100110", "00101000", "00101001", "00101011", "00101100", "00101110", "00101111", "00110001", "00110010", "00110100", "00110101", "00110111", "00111000", "00111001", "00111011", "00111100", 
"00111101", "00111111", "01000000", "01000001", "01000010", "01000011", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010001", 
"01010010", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101001", "10101010", "10101011", "10101011", "10101100", 
"10101101", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", 
"10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000000", 
"11000001", "11000001", "11000010", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000100", "11000101", "00111011", "00111011", "00111100", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", 
"00111110", "00111111", "00111111", "01000000", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", 
"01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010010", 
"01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101011", "10101011", 
"10101100", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111101", "10111110", "10111111", 
"11000000", "11000001", "11000011", "11000100", "11000101", "11000111", "11001000", "11001001", "11001011", "11001100", "11001110", "11001111", "11010001", "11010010", "11010100", "11010101", "11010111", "11011000", "11011010", "11011100", 
"11011101", "11011111", "11100001", "11100011", "11100100", "11100110", "11101000", "11101010", "11101011", "11101101", "11101111", "11110001", "11110011", "11110101", "11110111", "11111000", "11111010", "11111100", "11111110", "00000000", 
"00000010", "00000100", "00000110", "00001000", "00001010", "00001011", "00001101", "00001111", "00010001", "00010011", "00010101", "00010111", "00011001", "00011010", "00011100", "00011110", "00100000", "00100001", "00100011", "00100101", 
"00100111", "00101000", "00101010", "00101011", "00101101", "00101111", "00110000", "00110010", "00110011", "00110101", "00110110", "00110111", "00111001", "00111010", "00111011", "00111101", "00111110", "00111111", "01000001", "01000010", 
"01000011", "01000100", "01000101", "01000110", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010101", 
"01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10101111", 
"10110000", "10110000", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", 
"10111011", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000010", "11000011", 
"11000011", "11000100", "11000100", "11000100", "11000101", "11000101", "11000101", "00111010", "00111011", "00111011", "00111011", "00111100", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111110", "00111111", 
"00111111", "01000000", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", 
"01001000", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", 
"01010100", "01010101", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101110", 
"10101111", "10110000", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000001", "11000010", "11000011", 
"11000101", "11000110", "11000111", "11001001", "11001010", "11001011", "11001101", "11001110", "11010000", "11010001", "11010011", "11010101", "11010110", "11011000", "11011001", "11011011", "11011101", "11011111", "11100000", "11100010", 
"11100100", "11100110", "11100111", "11101001", "11101011", "11101101", "11101111", "11110001", "11110011", "11110101", "11110110", "11111000", "11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00001000", 
"00001010", "00001100", "00001110", "00010000", "00010001", "00010011", "00010101", "00010111", "00011001", "00011011", "00011101", "00011110", "00100000", "00100010", "00100100", "00100101", "00100111", "00101001", "00101010", "00101100", 
"00101110", "00101111", "00110001", "00110010", "00110100", "00110101", "00110111", "00111000", "00111001", "00111011", "00111100", "00111110", "00111111", "01000000", "01000001", "01000011", "01000100", "01000101", "01000110", "01000111", 
"01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01011000", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110010", 
"10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", 
"10111101", "10111110", "10111110", "10111111", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000100", "11000101", "11000101", 
"11000101", "11000110", "11000110", "00111010", "00111010", "00111010", "00111011", "00111011", "00111011", "00111100", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111110", "00111111", "00111111", "01000000", 
"01000000", "01000001", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", 
"01001010", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010100", "01010101", 
"01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", 
"10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111111", "11000000", "11000001", "11000010", "11000100", "11000101", "11000111", "11001000", 
"11001001", "11001011", "11001100", "11001110", "11001111", "11010001", "11010010", "11010100", "11010110", "11010111", "11011001", "11011011", "11011100", "11011110", "11100000", "11100010", "11100011", "11100101", "11100111", "11101001", 
"11101011", "11101101", "11101111", "11110000", "11110010", "11110100", "11110110", "11111000", "11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00001000", "00001010", "00001100", "00001110", "00010000", 
"00010010", "00010100", "00010110", "00010111", "00011001", "00011011", "00011101", "00011111", "00100001", "00100010", "00100100", "00100110", "00101000", "00101001", "00101011", "00101101", "00101110", "00110000", "00110001", "00110011", 
"00110100", "00110110", "00110111", "00111001", "00111010", "00111100", "00111101", "00111110", "01000000", "01000001", "01000010", "01000011", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", 
"01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", 
"10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110101", 
"10110110", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", 
"11000000", "11000000", "11000001", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000101", "11000110", "11000110", "11000110", "11000111", "00111001", 
"00111001", "00111010", "00111010", "00111010", "00111011", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "00111111", "01000000", "01000000", "01000001", 
"01000001", "01000010", "01000010", "01000011", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", 
"01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010110", "01010111", 
"01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", 
"10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111101", "10111110", "10111111", "11000000", "11000010", "11000011", "11000100", "11000110", "11000111", "11001001", "11001010", "11001100", "11001101", 
"11001111", "11010000", "11010010", "11010011", "11010101", "11010111", "11011000", "11011010", "11011100", "11011110", "11011111", "11100001", "11100011", "11100101", "11100111", "11101001", "11101010", "11101100", "11101110", "11110000", 
"11110010", "11110100", "11110110", "11111000", "11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00001000", "00001010", "00001100", "00001110", "00010000", "00010010", "00010100", "00010110", "00011000", 
"00011010", "00011100", "00011101", "00011111", "00100001", "00100011", "00100101", "00100110", "00101000", "00101010", "00101100", "00101101", "00101111", "00110000", "00110010", "00110100", "00110101", "00110111", "00111000", "00111010", 
"00111011", "00111100", "00111110", "00111111", "01000000", "01000010", "01000011", "01000100", "01000101", "01000110", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", 
"01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", 
"10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", 
"10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000000", "11000001", "11000001", "11000010", 
"11000010", "11000011", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000101", "11000110", "11000110", "11000110", "11000111", "11000111", "11001000", "00111000", "00111000", "00111001", "00111001", "00111010", 
"00111010", "00111010", "00111011", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000000", "01000001", "01000001", "01000010", 
"01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", 
"01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", 
"10111000", "10111010", "10111011", "10111100", "10111101", "10111110", "11000000", "11000001", "11000010", "11000100", "11000101", "11000110", "11001000", "11001001", "11001011", "11001100", "11001110", "11010000", "11010001", "11010011", 
"11010100", "11010110", "11011000", "11011010", "11011011", "11011101", "11011111", "11100001", "11100011", "11100100", "11100110", "11101000", "11101010", "11101100", "11101110", "11110000", "11110010", "11110100", "11110110", "11111000", 
"11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00001000", "00001010", "00001100", "00001110", "00010000", "00010010", "00010100", "00010110", "00011000", "00011010", "00011100", "00011110", "00100000", 
"00100010", "00100011", "00100101", "00100111", "00101001", "00101010", "00101100", "00101110", "00101111", "00110001", "00110011", "00110100", "00110110", "00110111", "00111001", "00111010", "00111100", "00111101", "00111110", "01000000", 
"01000001", "01000010", "01000100", "01000101", "01000110", "01000111", "01001000", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", 
"01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", 
"10110000", "10110001", "10110010", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111011", 
"10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", 
"11000101", "11000101", "11000101", "11000110", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001000", "00110111", "00111000", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111010", 
"00111011", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000001", "01000010", "01000010", "01000011", 
"01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", 
"01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", 
"10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10111000", "10111001", "10111010", "10111011", 
"10111100", "10111110", "10111111", "11000000", "11000010", "11000011", "11000100", "11000110", "11000111", "11001001", "11001010", "11001100", "11001101", "11001111", "11010001", "11010010", "11010100", "11010110", "11010111", "11011001", 
"11011011", "11011101", "11011110", "11100000", "11100010", "11100100", "11100110", "11101000", "11101010", "11101100", "11101110", "11110000", "11110010", "11110100", "11110110", "11111000", "11111010", "11111100", "11111110", "00000000", 
"00000010", "00000100", "00000110", "00001000", "00001010", "00001100", "00001110", "00010001", "00010011", "00010101", "00010111", "00011001", "00011010", "00011100", "00011110", "00100000", "00100010", "00100100", "00100110", "00101000", 
"00101001", "00101011", "00101101", "00101110", "00110000", "00110010", "00110011", "00110101", "00110111", "00111000", "00111010", "00111011", "00111100", "00111110", "00111111", "01000001", "01000010", "01000011", "01000100", "01000110", 
"01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001110", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110010", "10110011", 
"10110100", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", 
"10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000110", 
"11000111", "11000111", "11001000", "11001000", "11001000", "11001001", "11001001", "00110111", "00110111", "00110111", "00111000", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111010", "00111011", "00111011", 
"00111100", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", 
"01000101", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", "01001111", 
"01010000", "01010001", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", 
"10101011", "10101100", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110010", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111100", "10111101", "10111110", "10111111", 
"11000001", "11000010", "11000100", "11000101", "11000110", "11001000", "11001001", "11001011", "11001101", "11001110", "11010000", "11010010", "11010011", "11010101", "11010111", "11011000", "11011010", "11011100", "11011110", "11100000", 
"11100010", "11100100", "11100110", "11100111", "11101001", "11101011", "11101101", "11101111", "11110010", "11110100", "11110110", "11111000", "11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00001000", 
"00001011", "00001101", "00001111", "00010001", "00010011", "00010101", "00010111", "00011001", "00011011", "00011101", "00011111", "00100001", "00100011", "00100100", "00100110", "00101000", "00101010", "00101100", "00101101", "00101111", 
"00110001", "00110010", "00110100", "00110110", "00110111", "00111001", "00111010", "00111100", "00111101", "00111111", "01000000", "01000001", "01000011", "01000100", "01000101", "01000110", "01001000", "01001001", "01001010", "01001011", 
"01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", 
"10101010", "10101011", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", 
"10110111", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000001", 
"11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001000", "11001001", 
"11001001", "11001001", "11001010", "00110110", "00110110", "00110111", "00110111", "00110111", "00111000", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", 
"00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", 
"01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", 
"01010010", "01010011", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101100", "10101101", 
"10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111010", "10111011", "10111100", "10111101", "10111111", "11000000", "11000001", "11000011", "11000100", 
"11000110", "11000111", "11001001", "11001010", "11001100", "11001110", "11001111", "11010001", "11010011", "11010100", "11010110", "11011000", "11011010", "11011100", "11011101", "11011111", "11100001", "11100011", "11100101", "11100111", 
"11101001", "11101011", "11101101", "11101111", "11110001", "11110011", "11110101", "11111000", "11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000110", "00001001", "00001011", "00001101", "00001111", "00010001", 
"00010011", "00010101", "00010111", "00011001", "00011011", "00011101", "00011111", "00100001", "00100011", "00100101", "00100111", "00101001", "00101011", "00101100", "00101110", "00110000", "00110010", "00110011", "00110101", "00110110", 
"00111000", "00111010", "00111011", "00111101", "00111110", "00111111", "01000001", "01000010", "01000011", "01000101", "01000110", "01000111", "01001000", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", 
"01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", 
"10101101", "10101110", "10101111", "10110000", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111001", 
"10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111110", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", 
"11000100", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001000", "11001001", "11001001", "11001001", "11001010", "11001010", "11001010", "00110101", 
"00110110", "00110110", "00110110", "00110111", "00110111", "00110111", "00111000", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111100", "00111101", 
"00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", 
"01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010000", "01010001", "01010010", "01010011", "01010011", 
"01010100", "01010101", "01010101", "01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", 
"10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10111000", "10111001", "10111010", "10111011", "10111101", "10111110", "10111111", "11000001", "11000010", "11000011", "11000101", "11000110", "11001000", "11001010", 
"11001011", "11001101", "11001110", "11010000", "11010010", "11010100", "11010101", "11010111", "11011001", "11011011", "11011101", "11011111", "11100001", "11100011", "11100101", "11100111", "11101001", "11101011", "11101101", "11101111", 
"11110001", "11110011", "11110101", "11110111", "11111010", "11111100", "11111110", "00000000", "00000010", "00000100", "00000111", "00001001", "00001011", "00001101", "00001111", "00010001", "00010011", "00010110", "00011000", "00011010", 
"00011100", "00011110", "00100000", "00100010", "00100100", "00100110", "00101000", "00101001", "00101011", "00101101", "00101111", "00110001", "00110010", "00110100", "00110110", "00110111", "00111001", "00111010", "00111100", "00111101", 
"00111111", "01000000", "01000010", "01000011", "01000100", "01000110", "01000111", "01001000", "01001001", "01001010", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", 
"01010110", "01010111", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101000", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", 
"10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", 
"10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", 
"11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001000", "11001001", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001011", "00110100", "00110101", "00110101", "00110101", "00110110", 
"00110110", "00110111", "00110111", "00110111", "00111000", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111101", "00111110", 
"00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", 
"01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010101", "01010101", 
"01010110", "01010111", "01011000", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", 
"10110100", "10110110", "10110111", "10111000", "10111001", "10111010", "10111100", "10111101", "10111110", "11000000", "11000001", "11000011", "11000100", "11000110", "11000111", "11001001", "11001010", "11001100", "11001110", "11001111", 
"11010001", "11010011", "11010101", "11010111", "11011000", "11011010", "11011100", "11011110", "11100000", "11100010", "11100100", "11100110", "11101000", "11101010", "11101101", "11101111", "11110001", "11110011", "11110101", "11110111", 
"11111001", "11111100", "11111110", "00000000", "00000010", "00000100", "00000111", "00001001", "00001011", "00001101", "00001111", "00010010", "00010100", "00010110", "00011000", "00011010", "00011100", "00011110", "00100000", "00100010", 
"00100100", "00100110", "00101000", "00101010", "00101100", "00101110", "00110000", "00110001", "00110011", "00110101", "00110110", "00111000", "00111010", "00111011", "00111101", "00111110", "01000000", "01000001", "01000010", "01000100", 
"01000101", "01000110", "01001000", "01001001", "01001010", "01001011", "01001100", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110011", "10110011", "10110100", 
"10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", 
"11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", 
"11001000", "11001001", "11001001", "11001010", "11001010", "11001010", "11001011", "11001011", "11001011", "11001100", "11001100", "00110100", "00110100", "00110100", "00110101", "00110101", "00110101", "00110110", "00110110", "00110110", 
"00110111", "00110111", "00111000", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111101", "00111110", "00111110", "00111111", 
"00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001000", "01001001", "01001010", 
"01001010", "01001011", "01001100", "01001100", "01001101", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01010111", 
"01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110100", "10110101", "10110110", "10110111", 
"10111000", "10111010", "10111011", "10111100", "10111110", "10111111", "11000000", "11000010", "11000011", "11000101", "11000110", "11001000", "11001010", "11001011", "11001101", "11001111", "11010000", "11010010", "11010100", "11010110", 
"11011000", "11011010", "11011100", "11011110", "11100000", "11100010", "11100100", "11100110", "11101000", "11101010", "11101100", "11101110", "11110001", "11110011", "11110101", "11110111", "11111001", "11111100", "11111110", "00000000", 
"00000010", "00000101", "00000111", "00001001", "00001011", "00001110", "00010000", "00010010", "00010100", "00010110", "00011000", "00011011", "00011101", "00011111", "00100001", "00100011", "00100101", "00100111", "00101001", "00101011", 
"00101101", "00101110", "00110000", "00110010", "00110100", "00110101", "00110111", "00111001", "00111010", "00111100", "00111110", "00111111", "01000000", "01000010", "01000011", "01000101", "01000110", "01000111", "01001001", "01001010", 
"01001011", "01001100", "01001101", "01001110", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101001", 
"10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", 
"10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "11000000", "11000000", "11000001", "11000001", "11000001", "11000010", 
"11000010", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001010", 
"11001011", "11001011", "11001011", "11001100", "11001100", "11001100", "11001101", "00110011", "00110011", "00110100", "00110100", "00110100", "00110101", "00110101", "00110101", "00110110", "00110110", "00110110", "00110111", "00110111", 
"00111000", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "00111111", "01000000", 
"01000000", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", 
"01001100", "01001101", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011010", 
"10100111", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111001", "10111010", "10111011", 
"10111101", "10111110", "11000000", "11000001", "11000010", "11000100", "11000110", "11000111", "11001001", "11001011", "11001100", "11001110", "11010000", "11010010", "11010011", "11010101", "11010111", "11011001", "11011011", "11011101", 
"11011111", "11100001", "11100011", "11100101", "11101000", "11101010", "11101100", "11101110", "11110000", "11110010", "11110101", "11110111", "11111001", "11111011", "11111110", "00000000", "00000010", "00000101", "00000111", "00001001", 
"00001011", "00001110", "00010000", "00010010", "00010101", "00010111", "00011001", "00011011", "00011101", "00011111", "00100001", "00100011", "00100110", "00101000", "00101001", "00101011", "00101101", "00101111", "00110001", "00110011", 
"00110101", "00110110", "00111000", "00111010", "00111011", "00111101", "00111110", "01000000", "01000001", "01000011", "01000100", "01000110", "01000111", "01001000", "01001001", "01001011", "01001100", "01001101", "01001110", "01001111", 
"01010000", "01010001", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101100", "10101100", "10101101", 
"10101110", "10101111", "10101111", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", 
"10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000101", 
"11000101", "11000110", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001010", "11001011", "11001011", "11001011", "11001100", "11001100", "11001101", 
"11001101", "11001101", "11001110", "00110010", "00110010", "00110011", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", "00110101", "00110110", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", 
"00111000", "00111001", "00111001", "00111010", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", 
"01000010", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", 
"01001110", "01001110", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", 
"10101010", "10101011", "10101100", "10101100", "10101101", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110111", "10111000", "10111001", "10111010", "10111100", "10111101", "10111111", "11000000", 
"11000010", "11000011", "11000101", "11000110", "11001000", "11001010", "11001011", "11001101", "11001111", "11010001", "11010011", "11010101", "11010111", "11011000", "11011010", "11011101", "11011111", "11100001", "11100011", "11100101", 
"11100111", "11101001", "11101011", "11101110", "11110000", "11110010", "11110101", "11110111", "11111001", "11111011", "11111110", "00000000", "00000010", "00000101", "00000111", "00001001", "00001100", "00001110", "00010000", "00010011", 
"00010101", "00010111", "00011001", "00011100", "00011110", "00100000", "00100010", "00100100", "00100110", "00101000", "00101010", "00101100", "00101110", "00110000", "00110010", "00110100", "00110101", "00110111", "00111001", "00111010", 
"00111100", "00111110", "00111111", "01000001", "01000010", "01000100", "01000101", "01000110", "01001000", "01001001", "01001010", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", 
"01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101001", "10101010", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10110000", "10110000", "10110001", 
"10110010", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111110", 
"10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000101", "11000110", "11000110", "11000111", "11000111", 
"11001000", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001100", "11001101", "11001101", "11001101", "11001110", "11001110", "11001110", "00110001", 
"00110010", "00110010", "00110010", "00110011", "00110011", "00110011", "00110100", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", "00111000", "00111001", 
"00111001", "00111010", "00111010", "00111011", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", 
"01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", "01001110", "01001111", 
"01010000", "01010000", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010110", "01010111", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", 
"10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110110", "10110111", "10111000", "10111010", "10111011", "10111100", "10111110", "10111111", "11000001", "11000010", "11000100", "11000110", 
"11000111", "11001001", "11001011", "11001100", "11001110", "11010000", "11010010", "11010100", "11010110", "11011000", "11011010", "11011100", "11011110", "11100000", "11100010", "11100100", "11100111", "11101001", "11101011", "11101101", 
"11110000", "11110010", "11110100", "11110111", "11111001", "11111011", "11111110", "00000000", "00000010", "00000101", "00000111", "00001010", "00001100", "00001110", "00010001", "00010011", "00010101", "00011000", "00011010", "00011100", 
"00011110", "00100000", "00100011", "00100101", "00100111", "00101001", "00101011", "00101101", "00101111", "00110001", "00110011", "00110100", "00110110", "00111000", "00111010", "00111011", "00111101", "00111111", "01000000", "01000010", 
"01000011", "01000101", "01000110", "01000111", "01001001", "01001010", "01001011", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101101", "10101101", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", 
"10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "11000000", "11000000", "11000001", 
"11000001", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001000", "11001001", "11001001", "11001010", 
"11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001100", "11001101", "11001101", "11001101", "11001110", "11001110", "11001110", "11001111", "11001111", "00110001", "00110001", "00110001", "00110010", "00110010", 
"00110010", "00110011", "00110011", "00110011", "00110100", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", "00111000", "00111001", "00111001", "00111010", 
"00111010", "00111011", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", 
"01000100", "01000101", "01000110", "01000110", "01000111", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", 
"01010010", "01010011", "01010011", "01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", 
"10110000", "10110001", "10110010", "10110011", "10110101", "10110110", "10110111", "10111001", "10111010", "10111011", "10111101", "10111110", "11000000", "11000001", "11000011", "11000101", "11000110", "11001000", "11001010", "11001100", 
"11001101", "11001111", "11010001", "11010011", "11010101", "11010111", "11011001", "11011011", "11011101", "11100000", "11100010", "11100100", "11100110", "11101000", "11101011", "11101101", "11101111", "11110010", "11110100", "11110110", 
"11111001", "11111011", "11111110", "00000000", "00000010", "00000101", "00000111", "00001010", "00001100", "00001111", "00010001", "00010011", "00010110", "00011000", "00011010", "00011101", "00011111", "00100001", "00100011", "00100101", 
"00100111", "00101010", "00101100", "00101110", "00110000", "00110001", "00110011", "00110101", "00110111", "00111001", "00111011", "00111100", "00111110", "00111111", "01000001", "01000011", "01000100", "01000110", "01000111", "01001000", 
"01001010", "01001011", "01001100", "01001101", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", 
"10101010", "10101011", "10101100", "10101101", "10101110", "10101110", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111000", 
"10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", 
"11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001011", "11001100", "11001100", 
"11001100", "11001101", "11001101", "11001110", "11001110", "11001110", "11001111", "11001111", "11001111", "11010000", "11010000", "00110000", "00110000", "00110000", "00110001", "00110001", "00110001", "00110010", "00110010", "00110010", 
"00110011", "00110011", "00110100", "00110100", "00110100", "00110101", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111011", 
"00111011", "00111100", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", 
"01000110", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010010", "01010010", "01010011", 
"01010100", "01010101", "01010110", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110011", 
"10110100", "10110101", "10110110", "10111000", "10111001", "10111010", "10111100", "10111101", "10111111", "11000001", "11000010", "11000100", "11000101", "11000111", "11001001", "11001011", "11001101", "11001111", "11010000", "11010010", 
"11010100", "11010110", "11011001", "11011011", "11011101", "11011111", "11100001", "11100011", "11100110", "11101000", "11101010", "11101101", "11101111", "11110001", "11110100", "11110110", "11111001", "11111011", "11111110", "00000000", 
"00000010", "00000101", "00000111", "00001010", "00001100", "00001111", "00010001", "00010100", "00010110", "00011000", "00011011", "00011101", "00011111", "00100010", "00100100", "00100110", "00101000", "00101010", "00101100", "00101110", 
"00110000", "00110010", "00110100", "00110110", "00111000", "00111010", "00111011", "00111101", "00111111", "01000000", "01000010", "01000011", "01000101", "01000110", "01001000", "01001001", "01001011", "01001100", "01001101", "01001110", 
"01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101010", "10101011", "10101100", "10101101", "10101110", 
"10101111", "10101111", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111001", "10111010", "10111010", "10111011", "10111100", 
"10111100", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", 
"11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001101", "11001110", "11001110", "11001110", 
"11001111", "11001111", "11001111", "11010000", "11010000", "11010000", "11010001", "00101111", "00101111", "00110000", "00110000", "00110000", "00110001", "00110001", "00110001", "00110010", "00110010", "00110010", "00110011", "00110011", 
"00110011", "00110100", "00110100", "00110101", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111011", "00111011", "00111100", 
"00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", 
"01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", 
"01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110010", "10110011", "10110100", "10110101", "10110111", 
"10111000", "10111010", "10111011", "10111101", "10111110", "11000000", "11000001", "11000011", "11000101", "11000110", "11001000", "11001010", "11001100", "11001110", "11010000", "11010010", "11010100", "11010110", "11011000", "11011010", 
"11011100", "11011110", "11100001", "11100011", "11100101", "11101000", "11101010", "11101100", "11101111", "11110001", "11110100", "11110110", "11111001", "11111011", "11111110", "00000000", "00000011", "00000101", "00001000", "00001010", 
"00001101", "00001111", "00010010", "00010100", "00010110", "00011001", "00011011", "00011110", "00100000", "00100010", "00100100", "00100111", "00101001", "00101011", "00101101", "00101111", "00110001", "00110011", "00110101", "00110111", 
"00111001", "00111011", "00111100", "00111110", "01000000", "01000001", "01000011", "01000100", "01000110", "01000111", "01001001", "01001010", "01001100", "01001101", "01001110", "01001111", "01010001", "01010010", "01010011", "01010100", 
"01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101011", "10101100", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110010", 
"10110011", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111110", "10111111", 
"11000000", "11000000", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", 
"11001001", "11001010", "11001010", "11001011", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001101", "11001110", "11001110", "11001110", "11001111", "11001111", "11001111", "11010000", "11010000", "11010001", 
"11010001", "11010001", "11010001", "00101110", "00101111", "00101111", "00101111", "00101111", "00110000", "00110000", "00110001", "00110001", "00110001", "00110010", "00110010", "00110010", "00110011", "00110011", "00110011", "00110100", 
"00110100", "00110101", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", 
"00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", "01000110", "01000110", "01000111", "01001000", "01001000", 
"01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001101", "01001110", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010100", "01010101", "01010101", "01010110", "01010111", "01011000", 
"01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110001", "10110010", "10110011", "10110100", "10110110", "10110111", "10111001", "10111010", "10111100", 
"10111101", "10111111", "11000000", "11000010", "11000100", "11000101", "11000111", "11001001", "11001011", "11001101", "11001111", "11010001", "11010011", "11010101", "11010111", "11011001", "11011100", "11011110", "11100000", "11100010", 
"11100101", "11100111", "11101010", "11101100", "11101110", "11110001", "11110011", "11110110", "11111000", "11111011", "11111101", "00000000", "00000011", "00000101", "00001000", "00001010", "00001101", "00001111", "00010010", "00010100", 
"00010111", "00011001", "00011100", "00011110", "00100001", "00100011", "00100101", "00100111", "00101010", "00101100", "00101110", "00110000", "00110010", "00110100", "00110110", "00111000", "00111010", "00111100", "00111101", "00111111", 
"01000001", "01000010", "01000100", "01000101", "01000111", "01001000", "01001010", "01001011", "01001101", "01001110", "01001111", "01010000", "01010001", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101100", "10101101", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", 
"10110110", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111100", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000001", "11000001", "11000010", "11000010", 
"11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001100", 
"11001100", "11001100", "11001101", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11001111", "11010000", "11010000", "11010000", "11010001", "11010001", "11010001", "11010010", "11010010", "11010010", "00101101", 
"00101110", "00101110", "00101110", "00101111", "00101111", "00101111", "00110000", "00110000", "00110000", "00110001", "00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110011", "00110100", "00110100", "00110100", 
"00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", 
"00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001001", "01001010", "01001010", 
"01001011", "01001100", "01001100", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", 
"10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101111", "10110000", "10110001", "10110010", "10110011", "10110101", "10110110", "10111000", "10111001", "10111011", "10111100", "10111110", "10111111", "11000001", 
"11000011", "11000100", "11000110", "11001000", "11001010", "11001100", "11001110", "11010000", "11010010", "11010100", "11010110", "11011001", "11011011", "11011101", "11011111", "11100010", "11100100", "11100111", "11101001", "11101100", 
"11101110", "11110001", "11110011", "11110110", "11111000", "11111011", "11111101", "00000000", "00000011", "00000101", "00001000", "00001011", "00001101", "00010000", "00010010", "00010101", "00010111", "00011010", "00011100", "00011111", 
"00100001", "00100100", "00100110", "00101000", "00101010", "00101101", "00101111", "00110001", "00110011", "00110101", "00110111", "00111001", "00111011", "00111100", "00111110", "01000000", "01000010", "01000011", "01000101", "01000110", 
"01001000", "01001001", "01001011", "01001100", "01001110", "01001111", "01010000", "01010001", "01010010", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", 
"10101011", "10101100", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110001", "10110010", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", 
"10111010", "10111011", "10111100", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", 
"11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001100", "11001101", "11001101", "11001110", "11001110", 
"11001110", "11001111", "11001111", "11001111", "11010000", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010010", "11010010", "11010011", "11010011", "00101101", "00101101", "00101101", "00101110", "00101110", 
"00101110", "00101110", "00101111", "00101111", "00110000", "00110000", "00110000", "00110001", "00110001", "00110001", "00110010", "00110010", "00110010", "00110011", "00110011", "00110100", "00110100", "00110100", "00110101", "00110101", 
"00110110", "00110110", "00110111", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", "00111110", "00111111", 
"01000000", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001011", "01001100", 
"01001101", "01001110", "01001111", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", 
"10101011", "10101100", "10101110", "10101111", "10110000", "10110001", "10110010", "10110100", "10110101", "10110111", "10111000", "10111010", "10111011", "10111101", "10111110", "11000000", "11000010", "11000100", "11000101", "11000111", 
"11001001", "11001011", "11001101", "11001111", "11010001", "11010011", "11010110", "11011000", "11011010", "11011100", "11011111", "11100001", "11100100", "11100110", "11101001", "11101011", "11101110", "11110000", "11110011", "11110101", 
"11111000", "11111011", "11111101", "00000000", "00000011", "00000101", "00001000", "00001011", "00001101", "00010000", "00010011", "00010101", "00011000", "00011010", "00011101", "00011111", "00100010", "00100100", "00100111", "00101001", 
"00101011", "00101101", "00110000", "00110010", "00110100", "00110110", "00111000", "00111010", "00111100", "00111101", "00111111", "01000001", "01000011", "01000100", "01000110", "01000111", "01001001", "01001010", "01001100", "01001101", 
"01001111", "01010000", "01010001", "01010010", "01010011", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101101", "10101110", 
"10101111", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111001", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", 
"10111110", "10111110", "10111111", "11000000", "11000000", "11000001", "11000001", "11000010", "11000011", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", 
"11001001", "11001001", "11001010", "11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001101", "11001110", "11001110", "11001110", "11001111", "11001111", "11010000", "11010000", "11010000", 
"11010001", "11010001", "11010001", "11010010", "11010010", "11010010", "11010011", "11010011", "11010011", "11010100", "11010100", "00101100", "00101100", "00101100", "00101101", "00101101", "00101101", "00101110", "00101110", "00101110", 
"00101111", "00101111", "00101111", "00110000", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110010", "00110011", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", 
"00110110", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", "00111111", "00111111", "01000000", "01000000", 
"01000001", "01000010", "01000010", "01000011", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01000111", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001101", "01001110", "01001110", 
"01001111", "01010000", "01010001", "01010010", "01010011", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101101", "10101110", 
"10101111", "10110000", "10110001", "10110011", "10110100", "10110110", "10110111", "10111001", "10111010", "10111100", "10111101", "10111111", "11000001", "11000011", "11000100", "11000110", "11001000", "11001010", "11001100", "11001110", 
"11010000", "11010011", "11010101", "11010111", "11011001", "11011100", "11011110", "11100001", "11100011", "11100110", "11101000", "11101011", "11101101", "11110000", "11110011", "11110101", "11111000", "11111011", "11111101", "00000000", 
"00000011", "00000110", "00001000", "00001011", "00001110", "00010000", "00010011", "00010110", "00011000", "00011011", "00011110", "00100000", "00100011", "00100101", "00100111", "00101010", "00101100", "00101110", "00110000", "00110011", 
"00110101", "00110111", "00111001", "00111011", "00111101", "00111110", "01000000", "01000010", "01000100", "01000101", "01000111", "01001001", "01001010", "01001011", "01001101", "01001110", "01010000", "01010001", "01010010", "01010011", 
"01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110010", "10110011", 
"10110100", "10110100", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111110", "10111111", "10111111", "11000000", "11000001", 
"11000001", "11000010", "11000010", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001010", "11001011", 
"11001011", "11001100", "11001100", "11001101", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11001111", "11010000", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010010", "11010011", 
"11010011", "11010011", "11010100", "11010100", "11010100", "11010100", "11010101", "00101011", "00101011", "00101100", "00101100", "00101100", "00101100", "00101101", "00101101", "00101101", "00101110", "00101110", "00101110", "00101111", 
"00101111", "00110000", "00110000", "00110000", "00110001", "00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", "00110110", "00110111", 
"00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", 
"01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", 
"01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101101", "10101110", "10101111", "10110000", "10110010", 
"10110011", "10110101", "10110110", "10110111", "10111001", "10111011", "10111100", "10111110", "11000000", "11000010", "11000011", "11000101", "11000111", "11001001", "11001011", "11001101", "11010000", "11010010", "11010100", "11010110", 
"11011001", "11011011", "11011101", "11100000", "11100010", "11100101", "11101000", "11101010", "11101101", "11110000", "11110010", "11110101", "11111000", "11111010", "11111101", "00000000", "00000011", "00000110", "00001000", "00001011", 
"00001110", "00010001", "00010100", "00010110", "00011001", "00011100", "00011110", "00100001", "00100011", "00100110", "00101000", "00101011", "00101101", "00101111", "00110001", "00110100", "00110110", "00111000", "00111010", "00111100", 
"00111110", "01000000", "01000001", "01000011", "01000101", "01000110", "01001000", "01001010", "01001011", "01001101", "01001110", "01001111", "01010001", "01010010", "01010011", "01010100", "01010110", "01010111", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110101", "10110110", "10110111", 
"10111000", "10111000", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", 
"11000101", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001110", 
"11001110", "11001110", "11001111", "11001111", "11010000", "11010000", "11010000", "11010001", "11010001", "11010001", "11010010", "11010010", "11010010", "11010011", "11010011", "11010011", "11010100", "11010100", "11010100", "11010101", 
"11010101", "11010101", "11010110", "00101010", "00101010", "00101011", "00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", "00101101", "00101110", "00101110", "00101110", "00101111", "00101111", "00101111", 
"00110000", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110010", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", 
"00111000", "00111001", "00111001", "00111010", "00111010", "00111011", "00111011", "00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", 
"01000100", "01000101", "01000101", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001011", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010000", "01010001", "01010010", "01010011", 
"01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101100", "10101101", "10101110", "10101111", "10110001", "10110010", "10110011", "10110101", "10110110", 
"10111000", "10111010", "10111011", "10111101", "10111111", "11000000", "11000010", "11000100", "11000110", "11001000", "11001010", "11001100", "11001111", "11010001", "11010011", "11010101", "11011000", "11011010", "11011101", "11011111", 
"11100010", "11100100", "11100111", "11101010", "11101100", "11101111", "11110010", "11110101", "11111000", "11111010", "11111101", "00000000", "00000011", "00000110", "00001001", "00001011", "00001110", "00010001", "00010100", "00010111", 
"00011001", "00011100", "00011111", "00100001", "00100100", "00100111", "00101001", "00101011", "00101110", "00110000", "00110010", "00110101", "00110111", "00111001", "00111011", "00111101", "00111111", "01000001", "01000010", "01000100", 
"01000110", "01001000", "01001001", "01001011", "01001100", "01001110", "01001111", "01010000", "01010010", "01010011", "01010100", "01010101", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", 
"10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110010", "10110011", "10110100", "10110101", "10110110", "10110110", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", 
"10111100", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000011", "11000100", "11000101", "11000101", "11000110", "11000110", "11000111", "11000111", 
"11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11001111", "11010000", "11010000", 
"11010000", "11010001", "11010001", "11010010", "11010010", "11010010", "11010011", "11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010101", "11010110", "11010110", "11010110", "11010110", "00101001", 
"00101010", "00101010", "00101010", "00101010", "00101011", "00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", "00101101", "00101110", "00101110", "00101110", "00101111", "00101111", "00110000", "00110000", 
"00110000", "00110001", "00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110100", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", "00111001", 
"00111001", "00111010", "00111010", "00111011", "00111011", "00111100", "00111101", "00111101", "00111110", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000100", "01000101", 
"01000110", "01000110", "01000111", "01001000", "01001001", "01001010", "01001010", "01001011", "01001100", "01001101", "01001110", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", 
"01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101011", "10101100", "10101101", "10101110", "10110000", "10110001", "10110010", "10110100", "10110101", "10110111", "10111000", "10111010", "10111100", 
"10111110", "10111111", "11000001", "11000011", "11000101", "11000111", "11001001", "11001011", "11001110", "11010000", "11010010", "11010101", "11010111", "11011001", "11011100", "11011111", "11100001", "11100100", "11100111", "11101001", 
"11101100", "11101111", "11110010", "11110101", "11110111", "11111010", "11111101", "00000000", "00000011", "00000110", "00001001", "00001100", "00001111", "00010010", "00010100", "00010111", "00011010", "00011101", "00011111", "00100010", 
"00100101", "00100111", "00101010", "00101100", "00101111", "00110001", "00110011", "00110110", "00111000", "00111010", "00111100", "00111110", "01000000", "01000010", "01000100", "01000101", "01000111", "01001001", "01001010", "01001100", 
"01001101", "01001111", "01010000", "01010010", "01010011", "01010100", "01010101", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", 
"10110000", "10110001", "10110010", "10110011", "10110100", "10110100", "10110101", "10110110", "10110111", "10111000", "10111000", "10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", 
"11000000", "11000000", "11000001", "11000001", "11000010", "11000011", "11000011", "11000100", "11000100", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", 
"11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11001111", "11010000", "11010000", "11010001", "11010001", "11010001", "11010010", "11010010", "11010010", 
"11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010101", "11010101", "11010110", "11010110", "11010110", "11010111", "11010111", "11010111", "00101000", "00101001", "00101001", "00101001", "00101010", 
"00101010", "00101010", "00101011", "00101011", "00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", "00101110", "00101110", "00101110", "00101111", "00101111", "00101111", "00110000", "00110000", "00110001", 
"00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", 
"00111010", "00111011", "00111100", "00111100", "00111101", "00111101", "00111110", "00111111", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", 
"01001000", "01001000", "01001001", "01001010", "01001011", "01001100", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101001", "10101011", "10101100", "10101101", "10101110", "10110000", "10110001", "10110011", "10110100", "10110110", "10110111", "10111001", "10111011", "10111100", "10111110", "11000000", "11000010", 
"11000100", "11000110", "11001000", "11001010", "11001101", "11001111", "11010001", "11010100", "11010110", "11011001", "11011011", "11011110", "11100001", "11100011", "11100110", "11101001", "11101100", "11101110", "11110001", "11110100", 
"11110111", "11111010", "11111101", "00000000", "00000011", "00000110", "00001001", "00001100", "00001111", "00010010", "00010101", "00011000", "00011011", "00011101", "00100000", "00100011", "00100110", "00101000", "00101011", "00101101", 
"00110000", "00110010", "00110100", "00110111", "00111001", "00111011", "00111101", "00111111", "01000001", "01000011", "01000101", "01000110", "01001000", "01001010", "01001011", "01001101", "01001110", "01010000", "01010001", "01010011", 
"01010100", "01010101", "01010110", "01011000", "01011001", "01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", 
"10110101", "10110110", "10110110", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", 
"11000011", "11000100", "11000100", "11000101", "11000110", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", 
"11001110", "11001110", "11001110", "11001111", "11001111", "11010000", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010010", "11010011", "11010011", "11010011", "11010100", "11010100", "11010100", "11010101", 
"11010101", "11010101", "11010110", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", "11011000", "00101000", "00101000", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", 
"00101010", "00101011", "00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", "00101101", "00101110", "00101110", "00101110", "00101111", "00101111", "00110000", "00110000", "00110000", "00110001", "00110001", 
"00110010", "00110010", "00110010", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111010", "00111011", 
"00111100", "00111100", "00111101", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", 
"01001010", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", 
"10101010", "10101011", "10101100", "10101101", "10101111", "10110000", "10110010", "10110011", "10110101", "10110110", "10111000", "10111010", "10111011", "10111101", "10111111", "11000001", "11000011", "11000101", "11000111", "11001001", 
"11001100", "11001110", "11010000", "11010011", "11010101", "11011000", "11011010", "11011101", "11100000", "11100011", "11100101", "11101000", "11101011", "11101110", "11110001", "11110100", "11110111", "11111010", "11111101", "00000000", 
"00000011", "00000110", "00001001", "00001100", "00001111", "00010010", "00010101", "00011000", "00011011", "00011110", "00100001", "00100100", "00100110", "00101001", "00101100", "00101110", "00110001", "00110011", "00110101", "00111000", 
"00111010", "00111100", "00111110", "01000000", "01000010", "01000100", "01000110", "01001000", "01001001", "01001011", "01001101", "01001110", "01010000", "01010001", "01010010", "01010100", "01010101", "01010110", "01011000", "01011001", 
"01011010", "10100111", "10101000", "10101001", "10101010", "10101011", "10101101", "10101110", "10101111", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111000", 
"10111001", "10111010", "10111011", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", 
"11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11001111", "11010000", 
"11010000", "11010001", "11010001", "11010001", "11010010", "11010010", "11010011", "11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010101", "11010110", "11010110", "11010110", "11010111", "11010111", 
"11010111", "11011000", "11011000", "11011000", "11011000", "11011001", "11011001", "00100111", "00100111", "00100111", "00101000", "00101000", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101010", 
"00101011", "00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", "00101101", "00101110", "00101110", "00101111", "00101111", "00101111", "00110000", "00110000", "00110001", "00110001", "00110001", "00110010", 
"00110010", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111011", "00111011", "00111100", "00111100", 
"00111101", "00111110", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000101", "01000101", "01000110", "01000111", "01001000", "01001000", "01001001", "01001010", "01001011", 
"01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010001", "01010010", "01010011", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "10100111", "10101000", "10101010", "10101011", "10101100", 
"10101110", "10101111", "10110000", "10110010", "10110011", "10110101", "10110111", "10111000", "10111010", "10111100", "10111110", "11000000", "11000010", "11000100", "11000110", "11001000", "11001011", "11001101", "11001111", "11010010", 
"11010100", "11010111", "11011010", "11011100", "11011111", "11100010", "11100101", "11101000", "11101011", "11101110", "11110001", "11110100", "11110111", "11111010", "11111101", "00000000", "00000011", "00000110", "00001001", "00001101", 
"00010000", "00010011", "00010110", "00011001", "00011100", "00011111", "00100010", "00100100", "00100111", "00101010", "00101101", "00101111", "00110010", "00110100", "00110110", "00111001", "00111011", "00111101", "00111111", "01000001", 
"01000011", "01000101", "01000111", "01001001", "01001011", "01001100", "01001110", "01001111", "01010001", "01010010", "01010100", "01010101", "01010110", "01010111", "01011001", "01011010", "10100111", "10101000", "10101001", "10101011", 
"10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", 
"10111101", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", 
"11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11010000", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010010", 
"11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010101", "11010110", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", "11011000", "11011000", "11011001", "11011001", 
"11011001", "11011010", "11011010", "00100110", "00100110", "00100110", "00100111", "00100111", "00100111", "00101000", "00101000", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101010", "00101011", 
"00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", "00101110", "00101110", "00101110", "00101111", "00101111", "00110000", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110011", 
"00110011", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111110", 
"00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001101", 
"01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010111", "01011000", "01011001", "01011010", "10100111", "10101001", "10101010", "10101011", "10101100", "10101110", "10101111", "10110001", 
"10110010", "10110100", "10110101", "10110111", "10111001", "10111011", "10111101", "10111111", "11000001", "11000011", "11000101", "11000111", "11001010", "11001100", "11001110", "11010001", "11010011", "11010110", "11011001", "11011100", 
"11011110", "11100001", "11100100", "11100111", "11101010", "11101101", "11110000", "11110011", "11110111", "11111010", "11111101", "00000000", "00000011", "00000111", "00001010", "00001101", "00010000", "00010011", "00010110", "00011010", 
"00011101", "00100000", "00100010", "00100101", "00101000", "00101011", "00101110", "00110000", "00110011", "00110101", "00111000", "00111010", "00111100", "00111110", "01000001", "01000011", "01000101", "01000110", "01001000", "01001010", 
"01001100", "01001101", "01001111", "01010001", "01010010", "01010011", "01010101", "01010110", "01010111", "01011001", "01011010", "10100111", "10101000", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", 
"10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111100", "10111101", "10111110", "10111111", "10111111", "11000000", "11000001", 
"11000010", "11000010", "11000011", "11000100", "11000100", "11000101", "11000101", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001001", "11001010", "11001011", "11001011", "11001100", "11001100", "11001101", 
"11001101", "11001110", "11001110", "11001110", "11001111", "11001111", "11010000", "11010000", "11010001", "11010001", "11010001", "11010010", "11010010", "11010011", "11010011", "11010011", "11010100", "11010100", "11010101", "11010101", 
"11010101", "11010110", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", "11011000", "11011000", "11011001", "11011001", "11011001", "11011010", "11011010", "11011010", "11011010", "11011011", "00100101", 
"00100101", "00100110", "00100110", "00100110", "00100110", "00100111", "00100111", "00100111", "00101000", "00101000", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101010", "00101011", "00101011", 
"00101011", "00101100", "00101100", "00101101", "00101101", "00101101", "00101110", "00101110", "00101111", "00101111", "00101111", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110010", "00110011", "00110011", 
"00110100", "00110100", "00110101", "00110101", "00110110", "00110111", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111011", "00111011", "00111100", "00111100", "00111101", "00111110", "00111110", "00111111", 
"01000000", "01000001", "01000001", "01000010", "01000011", "01000100", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", 
"01010001", "01010010", "01010011", "01010100", "01010101", "01010110", "01011000", "01011001", "01011010", "10100111", "10101001", "10101010", "10101011", "10101101", "10101110", "10101111", "10110001", "10110011", "10110100", "10110110", 
"10111000", "10111010", "10111011", "10111101", "10111111", "11000010", "11000100", "11000110", "11001000", "11001011", "11001101", "11010000", "11010010", "11010101", "11011000", "11011011", "11011110", "11100000", "11100011", "11100110", 
"11101010", "11101101", "11110000", "11110011", "11110110", "11111001", "11111101", "00000000", "00000011", "00000111", "00001010", "00001101", "00010001", "00010100", "00010111", "00011010", "00011101", "00100000", "00100011", "00100110", 
"00101001", "00101100", "00101111", "00110001", "00110100", "00110110", "00111001", "00111011", "00111101", "01000000", "01000010", "01000100", "01000110", "01001000", "01001010", "01001011", "01001101", "01001111", "01010000", "01010010", 
"01010011", "01010101", "01010110", "01010111", "01011001", "01011010", "10100111", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", 
"10110110", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", 
"11000101", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11010000", 
"11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010010", "11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010101", "11010110", "11010110", "11010111", "11010111", "11010111", 
"11011000", "11011000", "11011000", "11011000", "11011001", "11011001", "11011001", "11011010", "11011010", "11011010", "11011011", "11011011", "11011011", "11011011", "11011100", "00100100", "00100100", "00100101", "00100101", "00100101", 
"00100101", "00100110", "00100110", "00100110", "00100111", "00100111", "00100111", "00101000", "00101000", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101011", "00101011", "00101011", "00101100", 
"00101100", "00101100", "00101101", "00101101", "00101110", "00101110", "00101110", "00101111", "00101111", "00110000", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110100", "00110100", 
"00110101", "00110101", "00110110", "00110110", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", 
"01000010", "01000010", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", 
"01010100", "01010101", "01010110", "01010111", "01011001", "01011010", "10100111", "10101001", "10101010", "10101011", "10101101", "10101110", "10110000", "10110001", "10110011", "10110101", "10110110", "10111000", "10111010", "10111100", 
"10111110", "11000000", "11000011", "11000101", "11000111", "11001010", "11001100", "11001111", "11010001", "11010100", "11010111", "11011010", "11011101", "11100000", "11100011", "11100110", "11101001", "11101100", "11101111", "11110011", 
"11110110", "11111001", "11111101", "00000000", "00000011", "00000111", "00001010", "00001110", "00010001", "00010100", "00011000", "00011011", "00011110", "00100001", "00100100", "00100111", "00101010", "00101101", "00110000", "00110010", 
"00110101", "00111000", "00111010", "00111100", "00111111", "01000001", "01000011", "01000101", "01000111", "01001001", "01001011", "01001101", "01001110", "01010000", "01010010", "01010011", "01010101", "01010110", "01010111", "01011001", 
"01011010", "10100111", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", 
"10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000011", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11000111", "11001000", "11001000", 
"11001001", "11001010", "11001010", "11001011", "11001011", "11001100", "11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11010000", "11010000", "11010001", "11010001", "11010001", "11010010", "11010010", 
"11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010101", "11010110", "11010110", "11010110", "11010111", "11010111", "11011000", "11011000", "11011000", "11011000", "11011001", "11011001", "11011001", 
"11011010", "11011010", "11011010", "11011011", "11011011", "11011011", "11011011", "11011100", "11011100", "11011100", "11011100", "00100011", "00100100", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100101", 
"00100110", "00100110", "00100110", "00100111", "00100111", "00100111", "00101000", "00101000", "00101000", "00101000", "00101001", "00101001", "00101010", "00101010", "00101010", "00101011", "00101011", "00101011", "00101100", "00101100", 
"00101100", "00101101", "00101101", "00101110", "00101110", "00101111", "00101111", "00101111", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", 
"00110110", "00110110", "00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111101", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", 
"01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010100", "01010101", "01010110", 
"01010111", "01011001", "01011010", "10100111", "10101001", "10101010", "10101011", "10101101", "10101110", "10110000", "10110010", "10110011", "10110101", "10110111", "10111001", "10111011", "10111101", "10111111", "11000001", "11000100", 
"11000110", "11001000", "11001011", "11001110", "11010000", "11010011", "11010110", "11011001", "11011100", "11011111", "11100010", "11100101", "11101000", "11101100", "11101111", "11110010", "11110110", "11111001", "11111101", "00000000", 
"00000100", "00000111", "00001011", "00001110", "00010001", "00010101", "00011000", "00011100", "00011111", "00100010", "00100101", "00101000", "00101011", "00101110", "00110001", "00110100", "00110110", "00111001", "00111011", "00111110", 
"01000000", "01000010", "01000100", "01000110", "01001000", "01001010", "01001100", "01001110", "01010000", "01010001", "01010011", "01010100", "01010110", "01010111", "01011001", "01011010", "10100111", "10101001", "10101010", "10101011", 
"10101100", "10101101", "10101110", "10110000", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", 
"10111111", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001010", "11001010", "11001011", "11001011", "11001100", 
"11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010011", "11010011", "11010011", "11010100", "11010100", "11010101", "11010101", 
"11010101", "11010110", "11010110", "11010110", "11010111", "11010111", "11011000", "11011000", "11011000", "11011000", "11011001", "11011001", "11011001", "11011010", "11011010", "11011010", "11011011", "11011011", "11011011", "11011100", 
"11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011101", "00100010", "00100011", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", 
"00100110", "00100110", "00100111", "00100111", "00100111", "00101000", "00101000", "00101000", "00101000", "00101001", "00101001", "00101010", "00101010", "00101010", "00101011", "00101011", "00101011", "00101100", "00101100", "00101101", 
"00101101", "00101101", "00101110", "00101110", "00101111", "00101111", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110100", "00110100", "00110101", "00110101", "00110110", "00110110", 
"00110111", "00111000", "00111000", "00111001", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000001", "01000001", "01000010", "01000011", "01000100", "01000101", 
"01000110", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010010", "01010011", "01010100", "01010101", "01010110", "01010111", "01011001", "01011010", 
"10100111", "10101001", "10101010", "10101100", "10101101", "10101111", "10110000", "10110010", "10110100", "10110110", "10111000", "10111010", "10111100", "10111110", "11000000", "11000010", "11000101", "11000111", "11001010", "11001100", 
"11001111", "11010010", "11010101", "11011000", "11011011", "11011110", "11100001", "11100100", "11101000", "11101011", "11101111", "11110010", "11110101", "11111001", "11111100", "00000000", "00000100", "00000111", "00001011", "00001110", 
"00010010", "00010101", "00011001", "00011100", "00100000", "00100011", "00100110", "00101001", "00101100", "00101111", "00110010", "00110101", "00110111", "00111010", "00111101", "00111111", "01000001", "01000100", "01000110", "01001000", 
"01001010", "01001100", "01001110", "01001111", "01010001", "01010011", "01010100", "01010110", "01010111", "01011000", "01011010", "10100111", "10101001", "10101010", "10101011", "10101100", "10101110", "10101111", "10110000", "10110001", 
"10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111110", "10111111", "11000000", "11000001", "11000010", "11000010", "11000011", 
"11000100", "11000101", "11000101", "11000110", "11000111", "11000111", "11001000", "11001000", "11001001", "11001010", "11001010", "11001011", "11001011", "11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", 
"11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010010", "11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010110", "11010110", "11010110", "11010111", "11010111", "11010111", 
"11011000", "11011000", "11011001", "11011001", "11011001", "11011001", "11011010", "11011010", "11011010", "11011011", "11011011", "11011011", "11011100", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011110", 
"11011110", "11011110", "11011110", "00100001", "00100010", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", "00100110", 
"00100110", "00100111", "00100111", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", 
"00101110", "00101110", "00101110", "00101111", "00101111", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110100", "00110101", "00110101", "00110110", "00110110", "00110111", "00111000", 
"00111000", "00111001", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111110", "00111110", "00111111", "01000000", "01000001", "01000010", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", 
"01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010100", "01010101", "01010110", "01010111", "01011001", "01011010", "10101000", "10101001", "10101010", 
"10101100", "10101101", "10101111", "10110001", "10110010", "10110100", "10110110", "10111000", "10111010", "10111100", "10111111", "11000001", "11000011", "11000110", "11001001", "11001011", "11001110", "11010001", "11010100", "11010111", 
"11011010", "11011101", "11100000", "11100100", "11100111", "11101011", "11101110", "11110010", "11110101", "11111001", "11111100", "00000000", "00000100", "00000111", "00001011", "00001111", "00010010", "00010110", "00011010", "00011101", 
"00100000", "00100100", "00100111", "00101010", "00101101", "00110000", "00110011", "00110110", "00111001", "00111011", "00111110", "01000000", "01000011", "01000101", "01000111", "01001001", "01001011", "01001101", "01001111", "01010001", 
"01010010", "01010100", "01010110", "01010111", "01011000", "01011010", "10101000", "10101001", "10101010", "10101011", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011", "10110101", "10110110", "10110111", 
"10111000", "10111001", "10111010", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", "11000111", 
"11001000", "11001001", "11001001", "11001010", "11001010", "11001011", "11001100", "11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", 
"11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010110", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011001", "11011010", "11011010", 
"11011010", "11011010", "11011011", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011101", "11011110", "11011110", "11011110", "11011110", "11011111", "11011111", "11011111", "00100001", 
"00100001", "00100001", "00100001", "00100010", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", "00100110", "00100110", 
"00100110", "00100111", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", "00101110", 
"00101110", "00101111", "00101111", "00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110100", "00110100", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", "00111001", 
"00111001", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", "00111111", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000110", "01000111", "01001000", "01001001", 
"01001010", "01001011", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011", "01010101", "01010110", "01010111", "01011000", "01011010", "10101000", "10101001", "10101010", "10101100", "10101110", "10101111", 
"10110001", "10110011", "10110101", "10110111", "10111001", "10111011", "10111101", "11000000", "11000010", "11000101", "11000111", "11001010", "11001101", "11010000", "11010011", "11010110", "11011001", "11011100", "11100000", "11100011", 
"11100110", "11101010", "11101110", "11110001", "11110101", "11111001", "11111100", "00000000", "00000100", "00001000", "00001011", "00001111", "00010011", "00010111", "00011010", "00011110", "00100001", "00100101", "00101000", "00101011", 
"00101111", "00110010", "00110101", "00110111", "00111010", "00111101", "00111111", "01000010", "01000100", "01000110", "01001001", "01001011", "01001101", "01001111", "01010000", "01010010", "01010100", "01010101", "01010111", "01011000", 
"01011010", "10101000", "10101001", "10101010", "10101011", "10101101", "10101110", "10101111", "10110000", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", 
"10111101", "10111110", "10111111", "11000000", "11000000", "11000001", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", "11000111", "11001000", "11001001", "11001001", "11001010", "11001010", "11001011", 
"11001100", "11001100", "11001101", "11001101", "11001110", "11001111", "11001111", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010011", "11010011", "11010011", "11010100", "11010100", "11010101", "11010101", 
"11010110", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011001", "11011010", "11011010", "11011010", "11011011", "11011011", "11011011", "11011100", "11011100", "11011100", 
"11011100", "11011101", "11011101", "11011101", "11011110", "11011110", "11011110", "11011110", "11011111", "11011111", "11011111", "11011111", "11100000", "11100000", "11100000", "00100000", "00100000", "00100000", "00100000", "00100001", 
"00100001", "00100001", "00100001", "00100010", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", "00100110", "00100110", 
"00100111", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101101", "00101101", "00101101", "00101110", "00101110", 
"00101111", "00101111", "00110000", "00110000", "00110001", "00110001", "00110010", "00110011", "00110011", "00110100", "00110100", "00110101", "00110110", "00110110", "00110111", "00110111", "00111000", "00111001", "00111001", "00111010", 
"00111011", "00111100", "00111100", "00111101", "00111110", "00111111", "01000000", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001100", 
"01001101", "01001110", "01010000", "01010001", "01010010", "01010011", "01010101", "01010110", "01010111", "01011000", "01011010", "10101000", "10101001", "10101011", "10101100", "10101110", "10110000", "10110001", "10110011", "10110101", 
"10110111", "10111010", "10111100", "10111110", "11000001", "11000011", "11000110", "11001001", "11001011", "11001110", "11010001", "11010101", "11011000", "11011011", "11011111", "11100010", "11100110", "11101001", "11101101", "11110001", 
"11110101", "11111000", "11111100", "00000000", "00000100", "00001000", "00001100", "00010000", "00010100", "00010111", "00011011", "00011111", "00100010", "00100110", "00101001", "00101101", "00110000", "00110011", "00110110", "00111001", 
"00111100", "00111110", "01000001", "01000011", "01000110", "01001000", "01001010", "01001100", "01001110", "01010000", "01010010", "01010100", "01010101", "01010111", "01011000", "01011010", "10101000", "10101001", "10101010", "10101100", 
"10101101", "10101110", "10101111", "10110001", "10110010", "10110011", "10110100", "10110101", "10110110", "10110111", "10111001", "10111010", "10111011", "10111100", "10111101", "10111101", "10111110", "10111111", "11000000", "11000001", 
"11000010", "11000011", "11000011", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001001", "11001010", "11001011", "11001011", "11001100", "11001100", "11001101", "11001110", "11001110", "11001111", 
"11001111", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010011", "11010011", "11010100", "11010100", "11010101", "11010101", "11010101", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", 
"11011000", "11011001", "11011001", "11011001", "11011010", "11011010", "11011010", "11011011", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011101", "11011110", "11011110", "11011110", 
"11011110", "11011111", "11011111", "11011111", "11100000", "11100000", "11100000", "11100000", "11100001", "11100001", "11100001", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100000", "00100001", 
"00100001", "00100001", "00100010", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", "00100110", "00100110", "00100111", 
"00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101011", "00101011", "00101011", "00101100", "00101100", "00101101", "00101101", "00101110", "00101110", "00101111", "00101111", 
"00110000", "00110000", "00110001", "00110001", "00110010", "00110010", "00110011", "00110100", "00110100", "00110101", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", 
"00111101", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000011", "01000100", "01000101", "01000110", "01000111", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", 
"01010001", "01010010", "01010011", "01010100", "01010110", "01010111", "01011000", "01011010", "10101000", "10101001", "10101011", "10101100", "10101110", "10110000", "10110010", "10110100", "10110110", "10111000", "10111010", "10111101", 
"10111111", "11000010", "11000100", "11000111", "11001010", "11001101", "11010000", "11010011", "11010111", "11011010", "11011110", "11100001", "11100101", "11101001", "11101100", "11110000", "11110100", "11111000", "11111100", "00000000", 
"00000100", "00001000", "00001100", "00010000", "00010100", "00011000", "00011100", "00100000", "00100011", "00100111", "00101010", "00101110", "00110001", "00110100", "00110111", "00111010", "00111101", "01000000", "01000010", "01000101", 
"01000111", "01001010", "01001100", "01001110", "01010000", "01010010", "01010011", "01010101", "01010111", "01011000", "01011010", "10101000", "10101001", "10101010", "10101100", "10101101", "10101110", "10110000", "10110001", "10110010", 
"10110011", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000010", "11000011", "11000100", "11000101", "11000110", 
"11000110", "11000111", "11001000", "11001001", "11001001", "11001010", "11001011", "11001011", "11001100", "11001101", "11001101", "11001110", "11001110", "11001111", "11001111", "11010000", "11010001", "11010001", "11010010", "11010010", 
"11010011", "11010011", "11010100", "11010100", "11010100", "11010101", "11010101", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011001", "11011010", "11011010", "11011010", 
"11011011", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011110", "11011110", "11011110", "11011110", "11011111", "11011111", "11011111", "11011111", "11100000", "11100000", "11100000", 
"11100000", "11100001", "11100001", "11100001", "11100001", "11100010", "11100010", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100000", "00100001", "00100001", 
"00100001", "00100001", "00100010", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", "00100110", "00100110", "00100111", "00100111", 
"00100111", "00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101100", "00101101", "00101101", "00101110", "00101110", "00101111", "00101111", "00110000", 
"00110001", "00110001", "00110010", "00110010", "00110011", "00110011", "00110100", "00110101", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111110", 
"00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001010", "01001011", "01001101", "01001110", "01001111", "01010000", "01010010", "01010011", 
"01010100", "01010110", "01010111", "01011000", "01011010", "10101000", "10101001", "10101011", "10101101", "10101110", "10110000", "10110010", "10110100", "10110110", "10111001", "10111011", "10111110", "11000000", "11000011", "11000110", 
"11001001", "11001100", "11001111", "11010010", "11010110", "11011001", "11011101", "11100000", "11100100", "11101000", "11101100", "11110000", "11110100", "11111000", "11111100", "00000000", "00000100", "00001000", "00001101", "00010001", 
"00010101", "00011001", "00011101", "00100001", "00100100", "00101000", "00101100", "00101111", "00110010", "00110110", "00111001", "00111100", "00111111", "01000001", "01000100", "01000110", "01001001", "01001011", "01001101", "01001111", 
"01010001", "01010011", "01010101", "01010111", "01011000", "01011010", "10101000", "10101001", "10101011", "10101100", "10101101", "10101111", "10110000", "10110001", "10110011", "10110100", "10110101", "10110110", "10110111", "10111000", 
"10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001001", "11001010", 
"11001011", "11001011", "11001100", "11001101", "11001101", "11001110", "11001111", "11001111", "11010000", "11010000", "11010001", "11010001", "11010010", "11010010", "11010011", "11010011", "11010100", "11010100", "11010101", "11010101", 
"11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011001", "11011010", "11011010", "11011010", "11011011", "11011011", "11011100", "11011100", "11011100", "11011100", "11011101", 
"11011101", "11011101", "11011110", "11011110", "11011110", "11011111", "11011111", "11011111", "11011111", "11100000", "11100000", "11100000", "11100000", "11100001", "11100001", "11100001", "11100001", "11100010", "11100010", "11100010", 
"11100010", "11100011", "11100011", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100000", "00100001", "00100001", 
"00100001", "00100001", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100100", "00100101", "00100101", "00100110", "00100110", "00100110", "00100111", "00100111", "00100111", 
"00101000", "00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101101", "00101101", "00101110", "00101110", "00101111", "00101111", "00110000", "00110000", "00110001", 
"00110001", "00110010", "00110011", "00110011", "00110100", "00110101", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "00111111", 
"01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001111", "01010000", "01010001", "01010011", "01010100", "01010101", "01010111", 
"01011000", "01011010", "10101000", "10101001", "10101011", "10101101", "10101111", "10110001", "10110011", "10110101", "10110111", "10111010", "10111100", "10111111", "11000001", "11000100", "11000111", "11001010", "11001110", "11010001", 
"11010100", "11011000", "11011100", "11011111", "11100011", "11100111", "11101011", "11101111", "11110011", "11111000", "11111100", "00000000", "00000100", "00001001", "00001101", "00010001", "00010110", "00011010", "00011110", "00100010", 
"00100110", "00101001", "00101101", "00110001", "00110100", "00110111", "00111010", "00111101", "01000000", "01000011", "01000110", "01001000", "01001010", "01001101", "01001111", "01010001", "01010011", "01010101", "01010111", "01011000", 
"01011010", "10101000", "10101001", "10101011", "10101100", "10101110", "10101111", "10110000", "10110010", "10110011", "10110100", "10110101", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", 
"10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001001", "11001010", "11001011", "11001100", "11001100", "11001101", "11001110", "11001110", 
"11001111", "11001111", "11010000", "11010001", "11010001", "11010010", "11010010", "11010011", "11010011", "11010100", "11010100", "11010101", "11010101", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", 
"11011001", "11011001", "11011001", "11011010", "11011010", "11011011", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011110", "11011110", "11011110", "11011110", "11011111", "11011111", 
"11011111", "11100000", "11100000", "11100000", "11100000", "11100001", "11100001", "11100001", "11100001", "11100010", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100011", "11100100", "11100100", "00011100", 
"00011100", "00011100", "00011101", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100000", "00100001", "00100001", 
"00100001", "00100010", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", "00100110", "00100111", "00100111", "00100111", "00101000", 
"00101000", "00101001", "00101001", "00101001", "00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101101", "00101101", "00101110", "00101110", "00101111", "00101111", "00110000", "00110001", "00110001", "00110010", 
"00110010", "00110011", "00110100", "00110100", "00110101", "00110110", "00110111", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", 
"01000011", "01000100", "01000101", "01000110", "01000111", "01001000", "01001001", "01001011", "01001100", "01001101", "01001110", "01010000", "01010001", "01010010", "01010100", "01010101", "01010111", "01011000", "01011010", "10101000", 
"10101001", "10101011", "10101101", "10101111", "10110001", "10110011", "10110110", "10111000", "10111010", "10111101", "11000000", "11000011", "11000110", "11001001", "11001100", "11001111", "11010011", "11010111", "11011010", "11011110", 
"11100010", "11100110", "11101010", "11101111", "11110011", "11110111", "11111100", "00000000", "00000101", "00001001", "00001110", "00010010", "00010110", "00011011", "00011111", "00100011", "00100111", "00101011", "00101110", "00110010", 
"00110101", "00111001", "00111100", "00111111", "01000010", "01000101", "01000111", "01001010", "01001100", "01001110", "01010001", "01010011", "01010101", "01010110", "01011000", "01011010", "10101000", "10101001", "10101011", "10101100", 
"10101110", "10101111", "10110001", "10110010", "10110011", "10110101", "10110110", "10110111", "10111000", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", 
"11000101", "11000110", "11000110", "11000111", "11001000", "11001001", "11001010", "11001010", "11001011", "11001100", "11001100", "11001101", "11001110", "11001110", "11001111", "11010000", "11010000", "11010001", "11010001", "11010010", 
"11010011", "11010011", "11010100", "11010100", "11010101", "11010101", "11010110", "11010110", "11010111", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011001", "11011010", "11011010", "11011011", "11011011", 
"11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011110", "11011110", "11011110", "11011111", "11011111", "11011111", "11100000", "11100000", "11100000", "11100000", "11100001", "11100001", "11100001", 
"11100001", "11100010", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100100", "11100100", "11100101", "00011011", "00011011", "00011100", "00011100", "00011100", 
"00011100", "00011100", "00011101", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100000", "00100001", "00100001", 
"00100001", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", "00100110", "00100111", "00100111", "00100111", "00101000", "00101000", 
"00101001", "00101001", "00101001", "00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101101", "00101101", "00101110", "00101111", "00101111", "00110000", "00110000", "00110001", "00110010", "00110010", "00110011", 
"00110100", "00110100", "00110101", "00110110", "00110110", "00110111", "00111000", "00111001", "00111010", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", 
"01000101", "01000110", "01001000", "01001001", "01001010", "01001011", "01001101", "01001110", "01001111", "01010001", "01010010", "01010100", "01010101", "01010111", "01011000", "01011010", "10101000", "10101010", "10101011", "10101101", 
"10101111", "10110010", "10110100", "10110110", "10111001", "10111011", "10111110", "11000001", "11000100", "11000111", "11001011", "11001110", "11010010", "11010101", "11011001", "11011101", "11100001", "11100101", "11101010", "11101110", 
"11110010", "11110111", "11111011", "00000000", "00000101", "00001001", "00001110", "00010011", "00010111", "00011100", "00100000", "00100100", "00101000", "00101100", "00110000", "00110100", "00110111", "00111010", "00111110", "01000001", 
"01000100", "01000110", "01001001", "01001100", "01001110", "01010000", "01010010", "01010100", "01010110", "01011000", "01011010", "10101000", "10101001", "10101011", "10101101", "10101110", "10110000", "10110001", "10110010", "10110100", 
"10110101", "10110110", "10111000", "10111001", "10111010", "10111011", "10111100", "10111110", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000101", "11000110", "11000111", "11001000", "11001001", 
"11001010", "11001010", "11001011", "11001100", "11001101", "11001101", "11001110", "11001111", "11001111", "11010000", "11010001", "11010001", "11010010", "11010010", "11010011", "11010011", "11010100", "11010100", "11010101", "11010101", 
"11010110", "11010110", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011010", "11011010", "11011010", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011110", 
"11011110", "11011110", "11011111", "11011111", "11011111", "11100000", "11100000", "11100000", "11100000", "11100001", "11100001", "11100001", "11100001", "11100010", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", 
"11100011", "11100100", "11100100", "11100100", "11100100", "11100101", "11100101", "11100101", "11100101", "11100101", "11100110", "00011010", "00011010", "00011011", "00011011", "00011011", "00011011", "00011011", "00011100", "00011100", 
"00011100", "00011100", "00011101", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100000", "00100001", "00100001", 
"00100001", "00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100110", "00100110", "00100110", "00100111", "00100111", "00101000", "00101000", "00101001", 
"00101001", "00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101101", "00101101", "00101110", "00101110", "00101111", "00101111", "00110000", "00110001", "00110001", "00110010", "00110011", "00110011", "00110100", 
"00110101", "00110110", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000100", "01000101", "01000110", "01000111", 
"01001000", "01001010", "01001011", "01001100", "01001110", "01001111", "01010000", "01010010", "01010011", "01010101", "01010111", "01011000", "01011010", "10101000", "10101010", "10101100", "10101110", "10110000", "10110010", "10110100", 
"10110111", "10111010", "10111100", "10111111", "11000010", "11000110", "11001001", "11001100", "11010000", "11010100", "11011000", "11011100", "11100000", "11100100", "11101001", "11101101", "11110010", "11110111", "11111011", "00000000", 
"00000101", "00001010", "00001111", "00010011", "00011000", "00011101", "00100001", "00100101", "00101010", "00101110", "00110001", "00110101", "00111001", "00111100", "00111111", "01000011", "01000110", "01001000", "01001011", "01001101", 
"01010000", "01010010", "01010100", "01010110", "01011000", "01011010", "10101000", "10101010", "10101011", "10101101", "10101110", "10110000", "10110001", "10110011", "10110100", "10110110", "10110111", "10111000", "10111010", "10111011", 
"10111100", "10111101", "10111110", "10111111", "11000000", "11000010", "11000011", "11000100", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001011", "11001100", "11001101", "11001110", 
"11001110", "11001111", "11010000", "11010000", "11010001", "11010001", "11010010", "11010011", "11010011", "11010100", "11010100", "11010101", "11010101", "11010110", "11010110", "11010111", "11010111", "11011000", "11011000", "11011001", 
"11011001", "11011010", "11011010", "11011010", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011110", "11011110", "11011110", "11011111", "11011111", "11011111", "11100000", "11100000", 
"11100000", "11100001", "11100001", "11100001", "11100001", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100100", "11100100", "11100101", "11100101", "11100101", 
"11100101", "11100110", "11100110", "11100110", "11100110", "11100110", "11100111", "00011001", "00011001", "00011010", "00011010", "00011010", "00011010", "00011010", "00011011", "00011011", "00011011", "00011011", "00011100", "00011100", 
"00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100001", "00100001", "00100001", 
"00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100110", "00100110", "00100110", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", 
"00101010", "00101010", "00101011", "00101011", "00101100", "00101100", "00101101", "00101101", "00101110", "00101111", "00101111", "00110000", "00110000", "00110001", "00110010", "00110010", "00110011", "00110100", "00110101", "00110101", 
"00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111100", "00111101", "00111110", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01001000", "01001001", "01001010", 
"01001100", "01001101", "01001111", "01010000", "01010010", "01010011", "01010101", "01010110", "01011000", "01011010", "10101000", "10101010", "10101100", "10101110", "10110000", "10110011", "10110101", "10111000", "10111010", "10111101", 
"11000001", "11000100", "11000111", "11001011", "11001111", "11010010", "11010110", "11011011", "11011111", "11100011", "11101000", "11101101", "11110001", "11110110", "11111011", "00000000", "00000101", "00001010", "00001111", "00010100", 
"00011001", "00011110", "00100010", "00100111", "00101011", "00101111", "00110011", "00110111", "00111011", "00111110", "01000001", "01000100", "01000111", "01001010", "01001101", "01001111", "01010010", "01010100", "01010110", "01011000", 
"01011010", "10101000", "10101010", "10101011", "10101101", "10101111", "10110000", "10110010", "10110011", "10110101", "10110110", "10111000", "10111001", "10111010", "10111011", "10111101", "10111110", "10111111", "11000000", "11000001", 
"11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001011", "11001100", "11001101", "11001110", "11001110", "11001111", "11010000", "11010001", "11010001", "11010010", 
"11010010", "11010011", "11010100", "11010100", "11010101", "11010101", "11010110", "11010110", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011010", "11011010", "11011011", "11011011", "11011011", "11011100", 
"11011100", "11011101", "11011101", "11011101", "11011110", "11011110", "11011110", "11011111", "11011111", "11011111", "11100000", "11100000", "11100000", "11100001", "11100001", "11100001", "11100001", "11100010", "11100010", "11100010", 
"11100011", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100100", "11100101", "11100101", "11100101", "11100101", "11100101", "11100110", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", 
"11100111", "11100111", "11100111", "00011000", "00011001", "00011001", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", "00011010", "00011011", "00011011", "00011011", "00011011", "00011011", "00011100", 
"00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100001", "00100001", "00100001", 
"00100010", "00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100101", "00100101", "00100101", "00100110", "00100110", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101010", 
"00101010", "00101011", "00101011", "00101100", "00101100", "00101101", "00101110", "00101110", "00101111", "00101111", "00110000", "00110001", "00110010", "00110010", "00110011", "00110100", "00110101", "00110101", "00110110", "00110111", 
"00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000101", "01000110", "01000111", "01001000", "01001010", "01001011", "01001101", "01001110", 
"01010000", "01010001", "01010011", "01010101", "01010110", "01011000", "01011010", "10101000", "10101010", "10101100", "10101110", "10110001", "10110011", "10110110", "10111001", "10111100", "10111111", "11000010", "11000101", "11001001", 
"11001101", "11010001", "11010101", "11011001", "11011110", "11100010", "11100111", "11101100", "11110001", "11110110", "11111011", "00000000", "00000101", "00001011", "00010000", "00010101", "00011010", "00011111", "00100100", "00101000", 
"00101101", "00110001", "00110101", "00111001", "00111100", "01000000", "01000011", "01000110", "01001001", "01001100", "01001111", "01010001", "01010100", "01010110", "01011000", "01011010", "10101000", "10101010", "10101100", "10101101", 
"10101111", "10110001", "10110010", "10110100", "10110101", "10110111", "10111000", "10111010", "10111011", "10111100", "10111101", "10111111", "11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", 
"11001000", "11001001", "11001010", "11001011", "11001100", "11001100", "11001101", "11001110", "11001111", "11001111", "11010000", "11010001", "11010010", "11010010", "11010011", "11010011", "11010100", "11010101", "11010101", "11010110", 
"11010110", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011010", "11011010", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011101", "11011110", "11011110", "11011111", 
"11011111", "11011111", "11100000", "11100000", "11100000", "11100001", "11100001", "11100001", "11100001", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100100", 
"11100101", "11100101", "11100101", "11100101", "11100110", "11100110", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101000", "11101000", "00010111", 
"00011000", "00011000", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", "00011010", "00011010", "00011011", "00011011", "00011011", "00011011", "00011100", 
"00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100001", "00100001", "00100001", 
"00100010", "00100010", "00100011", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100110", "00100110", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101010", "00101010", 
"00101011", "00101011", "00101100", "00101101", "00101101", "00101110", "00101110", "00101111", "00110000", "00110001", "00110001", "00110010", "00110011", "00110100", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", 
"00111010", "00111011", "00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000011", "01000100", "01000101", "01000110", "01001000", "01001001", "01001011", "01001100", "01001110", "01001111", "01010001", "01010011", 
"01010100", "01010110", "01011000", "01011010", "10101000", "10101010", "10101100", "10101111", "10110001", "10110100", "10110111", "10111010", "10111101", "11000000", "11000100", "11000111", "11001011", "11001111", "11010011", "11011000", 
"11011100", "11100001", "11100110", "11101011", "11110000", "11110101", "11111011", "00000000", "00000110", "00001011", "00010000", "00010110", "00011011", "00100000", "00100101", "00101010", "00101110", "00110011", "00110111", "00111011", 
"00111110", "01000010", "01000101", "01001001", "01001011", "01001110", "01010001", "01010011", "01010110", "01011000", "01011010", "10101000", "10101010", "10101100", "10101110", "10101111", "10110001", "10110011", "10110100", "10110110", 
"10110111", "10111001", "10111010", "10111100", "10111101", "10111110", "10111111", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", 
"11001101", "11001110", "11001111", "11010000", "11010000", "11010001", "11010010", "11010011", "11010011", "11010100", "11010100", "11010101", "11010110", "11010110", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", 
"11011010", "11011010", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011110", "11011110", "11011110", "11011111", "11011111", "11100000", "11100000", "11100000", "11100001", "11100001", "11100001", 
"11100010", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100100", "11100101", "11100101", "11100101", "11100101", "11100110", "11100110", "11100110", "11100110", "11100110", 
"11100111", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101000", "11101000", "11101000", "11101001", "11101001", "11101001", "11101001", "11101001", "00010110", "00010111", "00010111", "00010111", "00010111", 
"00010111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", "00011010", "00011010", "00011011", "00011011", "00011011", "00011011", 
"00011100", "00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00100000", "00100000", "00100000", "00100001", "00100001", "00100010", 
"00100010", "00100010", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100110", "00100110", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101010", "00101010", "00101011", 
"00101100", "00101100", "00101101", "00101101", "00101110", "00101111", "00110000", "00110000", "00110001", "00110010", "00110011", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", 
"00111100", "00111101", "00111110", "00111111", "01000001", "01000010", "01000011", "01000100", "01000110", "01000111", "01001001", "01001010", "01001100", "01001101", "01001111", "01010001", "01010010", "01010100", "01010110", "01011000", 
"01011010", "10101000", "10101010", "10101101", "10101111", "10110010", "10110101", "10110111", "10111011", "10111110", "11000010", "11000101", "11001001", "11001101", "11010010", "11010110", "11011011", "11100000", "11100101", "11101010", 
"11110000", "11110101", "11111010", "00000000", "00000110", "00001011", "00010001", "00010111", "00011100", "00100001", "00100111", "00101011", "00110000", "00110101", "00111001", "00111101", "01000001", "01000100", "01001000", "01001011", 
"01001110", "01010000", "01010011", "01010101", "01011000", "01011010", "10101000", "10101010", "10101100", "10101110", "10110000", "10110010", "10110011", "10110101", "10110110", "10111000", "10111010", "10111011", "10111100", "10111110", 
"10111111", "11000000", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11001111", "11010000", "11010001", "11010010", 
"11010010", "11010011", "11010100", "11010100", "11010101", "11010110", "11010110", "11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011010", "11011010", "11011011", "11011011", "11011100", "11011100", "11011101", 
"11011101", "11011110", "11011110", "11011110", "11011111", "11011111", "11011111", "11100000", "11100000", "11100001", "11100001", "11100001", "11100010", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100100", 
"11100100", "11100100", "11100100", "11100101", "11100101", "11100101", "11100101", "11100110", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101000", "11101000", 
"11101001", "11101001", "11101001", "11101001", "11101001", "11101001", "11101010", "11101010", "11101010", "11101010", "11101010", "00010110", "00010110", "00010110", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", 
"00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", "00011010", "00011011", "00011011", "00011011", "00011011", 
"00011100", "00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011110", "00011111", "00011111", "00011111", "00100000", "00100000", "00100001", "00100001", "00100001", "00100010", 
"00100010", "00100010", "00100011", "00100011", "00100100", "00100100", "00100101", "00100101", "00100110", "00100110", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101010", "00101010", "00101011", "00101100", 
"00101100", "00101101", "00101110", "00101110", "00101111", "00110000", "00110001", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", 
"00111110", "01000000", "01000001", "01000010", "01000100", "01000101", "01000110", "01001000", "01001010", "01001011", "01001101", "01001110", "01010000", "01010010", "01010100", "01010110", "01011000", "01011010", "10101000", "10101011", 
"10101101", "10110000", "10110010", "10110101", "10111000", "10111100", "10111111", "11000011", "11000111", "11001011", "11010000", "11010101", "11011001", "11011111", "11100100", "11101001", "11101111", "11110101", "11111010", "00000000", 
"00000110", "00001100", "00010010", "00011000", "00011101", "00100011", "00101000", "00101101", "00110010", "00110111", "00111011", "00111111", "01000011", "01000110", "01001010", "01001101", "01010000", "01010011", "01010101", "01011000", 
"01011010", "10101000", "10101010", "10101100", "10101110", "10110000", "10110010", "10110100", "10110110", "10110111", "10111001", "10111010", "10111100", "10111101", "10111111", "11000000", "11000001", "11000011", "11000100", "11000101", 
"11000110", "11000111", "11001000", "11001001", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010000", "11010001", "11010010", "11010011", "11010011", "11010100", "11010101", "11010101", "11010110", 
"11010111", "11010111", "11011000", "11011000", "11011001", "11011001", "11011010", "11011011", "11011011", "11011100", "11011100", "11011100", "11011101", "11011101", "11011110", "11011110", "11011111", "11011111", "11011111", "11100000", 
"11100000", "11100000", "11100001", "11100001", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100101", "11100101", "11100101", "11100101", "11100110", "11100110", 
"11100110", "11100110", "11100111", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101000", "11101000", "11101001", "11101001", "11101001", "11101001", "11101001", "11101010", "11101010", "11101010", "11101010", 
"11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101011", "00010101", "00010101", "00010101", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010110", "00010110", "00010110", "00010111", 
"00010111", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", "00011010", "00011011", "00011011", "00011011", 
"00011011", "00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011111", "00011111", "00100000", "00100000", "00100000", "00100001", "00100001", "00100001", "00100010", 
"00100010", "00100011", "00100011", "00100100", "00100100", "00100100", "00100101", "00100101", "00100110", "00100111", "00100111", "00101000", "00101000", "00101001", "00101001", "00101010", "00101011", "00101011", "00101100", "00101101", 
"00101101", "00101110", "00101111", "00110000", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111101", "00111111", "01000000", 
"01000001", "01000011", "01000100", "01000110", "01000111", "01001001", "01001010", "01001100", "01001110", "01010000", "01010010", "01010100", "01010110", "01011000", "01011010", "10101000", "10101011", "10101101", "10110000", "10110011", 
"10110110", "10111010", "10111101", "11000001", "11000101", "11001001", "11001110", "11010011", "11011000", "11011101", "11100011", "11101000", "11101110", "11110100", "11111010", "00000000", "00000110", "00001101", "00010011", "00011001", 
"00011111", "00100100", "00101010", "00101111", "00110100", "00111001", "00111101", "01000001", "01000101", "01001001", "01001100", "01001111", "01010010", "01010101", "01010111", "01011010", "10101000", "10101011", "10101101", "10101111", 
"10110001", "10110011", "10110100", "10110110", "10111000", "10111010", "10111011", "10111101", "10111110", "11000000", "11000001", "11000010", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011", 
"11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010010", "11010011", "11010100", "11010101", "11010101", "11010110", "11010111", "11010111", "11011000", "11011000", "11011001", "11011010", "11011010", 
"11011011", "11011011", "11011100", "11011100", "11011101", "11011101", "11011110", "11011110", "11011110", "11011111", "11011111", "11100000", "11100000", "11100000", "11100001", "11100001", "11100010", "11100010", "11100010", "11100011", 
"11100011", "11100011", "11100100", "11100100", "11100100", "11100100", "11100101", "11100101", "11100101", "11100110", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", 
"11101000", "11101000", "11101001", "11101001", "11101001", "11101001", "11101001", "11101010", "11101010", "11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", 
"11101100", "11101100", "11101100", "00010100", "00010100", "00010100", "00010100", "00010100", "00010100", "00010101", "00010101", "00010101", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010110", "00010110", 
"00010111", "00010111", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", "00011010", "00011011", "00011011", 
"00011011", "00011100", "00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011111", "00011111", "00100000", "00100000", "00100000", "00100001", "00100001", "00100010", "00100010", 
"00100010", "00100011", "00100011", "00100100", "00100100", "00100101", "00100101", "00100110", "00100110", "00100111", "00101000", "00101000", "00101001", "00101001", "00101010", "00101011", "00101011", "00101100", "00101101", "00101110", 
"00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011", "00111100", "00111110", "00111111", "01000000", "01000010", "01000011", 
"01000101", "01000110", "01001000", "01001010", "01001100", "01001101", "01001111", "01010001", "01010011", "01010101", "01011000", "01011010", "10101001", "10101011", "10101110", "10110001", "10110100", "10110111", "10111011", "10111111", 
"11000011", "11000111", "11001100", "11010001", "11010110", "11011100", "11100001", "11100111", "11101101", "11110011", "11111010", "00000000", "00000111", "00001101", "00010100", "00011010", "00100000", "00100110", "00101100", "00110001", 
"00110110", "00111011", "01000000", "01000100", "01001000", "01001011", "01001111", "01010010", "01010101", "01010111", "01011010", "10101001", "10101011", "10101101", "10101111", "10110001", "10110011", "10110101", "10110111", "10111001", 
"10111010", "10111100", "10111110", "10111111", "11000001", "11000010", "11000011", "11000101", "11000110", "11000111", "11001000", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010000", "11010001", 
"11010010", "11010011", "11010100", "11010100", "11010101", "11010110", "11010111", "11010111", "11011000", "11011000", "11011001", "11011010", "11011010", "11011011", "11011011", "11011100", "11011100", "11011101", "11011101", "11011110", 
"11011110", "11011111", "11011111", "11100000", "11100000", "11100000", "11100001", "11100001", "11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100101", "11100101", "11100101", 
"11100101", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101000", "11101001", "11101001", "11101001", "11101001", "11101001", "11101010", "11101010", "11101010", 
"11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", "11101100", "11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101101", "00010011", 
"00010011", "00010011", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", "00010100", "00010100", "00010100", "00010101", "00010101", "00010101", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", 
"00010110", "00010110", "00010111", "00010111", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", "00011011", "00011011", 
"00011011", "00011011", "00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011111", "00011111", "00100000", "00100000", "00100000", "00100001", "00100001", "00100010", "00100010", 
"00100011", "00100011", "00100100", "00100100", "00100101", "00100101", "00100110", "00100110", "00100111", "00101000", "00101000", "00101001", "00101001", "00101010", "00101011", "00101100", "00101100", "00101101", "00101110", "00101111", 
"00110000", "00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00111000", "00111001", "00111010", "00111011", "00111101", "00111110", "00111111", "01000001", "01000010", "01000100", "01000110", "01000111", 
"01001001", "01001011", "01001101", "01001111", "01010001", "01010011", "01010101", "01010111", "01011010", "10101001", "10101011", "10101110", "10110001", "10110101", "10111000", "10111100", "11000000", "11000101", "11001010", "11001111", 
"11010100", "11011010", "11100000", "11100110", "11101100", "11110011", "11111001", "00000000", "00000111", "00001110", "00010101", "00011100", "00100010", "00101000", "00101110", "00110100", "00111001", "00111110", "01000010", "01000110", 
"01001010", "01001110", "01010001", "01010100", "01010111", "01011010", "10101001", "10101011", "10101101", "10110000", "10110010", "10110100", "10110110", "10111000", "10111010", "10111011", "10111101", "10111111", "11000000", "11000010", 
"11000011", "11000101", "11000110", "11000111", "11001000", "11001010", "11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010011", "11010100", "11010101", "11010110", "11010110", 
"11010111", "11011000", "11011000", "11011001", "11011010", "11011010", "11011011", "11011100", "11011100", "11011101", "11011101", "11011110", "11011110", "11011111", "11011111", "11100000", "11100000", "11100000", "11100001", "11100001", 
"11100010", "11100010", "11100010", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100101", "11100101", "11100101", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", "11100111", "11101000", 
"11101000", "11101000", "11101000", "11101001", "11101001", "11101001", "11101001", "11101010", "11101010", "11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", 
"11101100", "11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101110", "11101110", "11101110", "11101110", "11101110", "00010010", "00010010", "00010010", "00010010", "00010010", 
"00010010", "00010011", "00010011", "00010011", "00010011", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", "00010100", "00010100", "00010101", "00010101", "00010101", "00010101", "00010101", "00010101", "00010110", 
"00010110", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", "00011011", 
"00011011", "00011011", "00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011110", "00011110", "00011110", "00011111", "00011111", "00100000", "00100000", "00100000", "00100001", "00100001", "00100010", "00100010", 
"00100011", "00100011", "00100100", "00100100", "00100101", "00100110", "00100110", "00100111", "00101000", "00101000", "00101001", "00101010", "00101010", "00101011", "00101100", "00101101", "00101101", "00101110", "00101111", "00110000", 
"00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00111000", "00111001", "00111010", "00111011", "00111101", "00111110", "01000000", "01000001", "01000011", "01000101", "01000110", "01001000", "01001010", "01001100", 
"01001110", "01010000", "01010011", "01010101", "01010111", "01011010", "10101001", "10101100", "10101111", "10110010", "10110110", "10111010", "10111110", "11000010", "11000111", "11001100", "11010010", "11011000", "11011110", "11100100", 
"11101011", "11110010", "11111001", "00000000", "00000111", "00001111", "00010110", "00011101", "00100100", "00101010", "00110000", "00110110", "00111011", "01000000", "01000101", "01001001", "01001101", "01010001", "01010100", "01010111", 
"01011010", "10101001", "10101011", "10101110", "10110000", "10110010", "10110101", "10110111", "10111001", "10111010", "10111100", "10111110", "11000000", "11000001", "11000011", "11000100", "11000110", "11000111", "11001001", "11001010", 
"11001011", "11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010110", "11010111", "11011000", "11011001", "11011001", "11011010", "11011010", "11011011", 
"11011100", "11011100", "11011101", "11011101", "11011110", "11011110", "11011111", "11011111", "11100000", "11100000", "11100001", "11100001", "11100010", "11100010", "11100010", "11100011", "11100011", "11100100", "11100100", "11100100", 
"11100101", "11100101", "11100101", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101000", "11101001", "11101001", "11101001", "11101001", "11101010", "11101010", 
"11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", "11101100", "11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101110", 
"11101110", "11101110", "11101110", "11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11101111", "11101111", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", 
"00010010", "00010010", "00010010", "00010010", "00010011", "00010011", "00010011", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", "00010100", "00010100", "00010100", "00010101", "00010101", "00010101", "00010101", 
"00010101", "00010110", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", 
"00011011", "00011011", "00011011", "00011100", "00011100", "00011100", "00011101", "00011101", "00011110", "00011110", "00011110", "00011111", "00011111", "00100000", "00100000", "00100001", "00100001", "00100010", "00100010", "00100011", 
"00100011", "00100100", "00100100", "00100101", "00100110", "00100110", "00100111", "00100111", "00101000", "00101001", "00101010", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", 
"00110011", "00110100", "00110101", "00110110", "00110111", "00111001", "00111010", "00111100", "00111101", "00111111", "01000000", "01000010", "01000100", "01000110", "01000111", "01001001", "01001011", "01001110", "01010000", "01010010", 
"01010101", "01010111", "01011010", "10101001", "10101100", "10101111", "10110011", "10110111", "10111011", "11000000", "11000101", "11001010", "11010000", "11010110", "11011100", "11100011", "11101010", "11110001", "11111001", "00000000", 
"00001000", "00010000", "00010111", "00011111", "00100110", "00101101", "00110011", "00111001", "00111110", "01000011", "01001000", "01001100", "01010000", "01010100", "01010111", "01011010", "10101001", "10101100", "10101110", "10110001", 
"10110011", "10110101", "10110111", "10111010", "10111100", "10111101", "10111111", "11000001", "11000011", "11000100", "11000110", "11000111", "11001001", "11001010", "11001011", "11001100", "11001110", "11001111", "11010000", "11010001", 
"11010010", "11010011", "11010100", "11010101", "11010101", "11010110", "11010111", "11011000", "11011001", "11011001", "11011010", "11011011", "11011011", "11011100", "11011101", "11011101", "11011110", "11011110", "11011111", "11011111", 
"11100000", "11100000", "11100001", "11100001", "11100010", "11100010", "11100011", "11100011", "11100011", "11100100", "11100100", "11100100", "11100101", "11100101", "11100110", "11100110", "11100110", "11100110", "11100111", "11100111", 
"11100111", "11101000", "11101000", "11101000", "11101001", "11101001", "11101001", "11101001", "11101010", "11101010", "11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", 
"11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101101", "11101101", "11101110", "11101110", "11101110", "11101110", "11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11101111", "11101111", 
"11101111", "11101111", "11110000", "11110000", "11110000", "11110000", "11110000", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", 
"00010010", "00010010", "00010010", "00010010", "00010010", "00010010", "00010010", "00010011", "00010011", "00010011", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", "00010100", "00010100", "00010101", "00010101", 
"00010101", "00010101", "00010110", "00010110", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011010", "00011010", "00011010", 
"00011010", "00011011", "00011011", "00011100", "00011100", "00011100", "00011101", "00011101", "00011101", "00011110", "00011110", "00011111", "00011111", "00100000", "00100000", "00100001", "00100001", "00100010", "00100010", "00100011", 
"00100011", "00100100", "00100101", "00100101", "00100110", "00100111", "00100111", "00101000", "00101001", "00101010", "00101011", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110100", 
"00110101", "00110110", "00110111", "00111001", "00111010", "00111100", "00111101", "00111111", "01000001", "01000011", "01000100", "01000110", "01001001", "01001011", "01001101", "01001111", "01010010", "01010100", "01010111", "01011010", 
"10101001", "10101100", "10110000", "10110100", "10111000", "10111101", "11000010", "11000111", "11001101", "11010011", "11011010", "11100001", "11101001", "11110000", "11111000", "00000000", "00001000", "00010001", "00011001", "00100001", 
"00101000", "00101111", "00110110", "00111100", "01000001", "01000110", "01001011", "01001111", "01010011", "01010111", "01011010", "10101001", "10101100", "10101111", "10110001", "10110100", "10110110", "10111000", "10111011", "10111101", 
"10111111", "11000001", "11000010", "11000100", "11000110", "11000111", "11001001", "11001010", "11001011", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", 
"11011000", "11011001", "11011001", "11011010", "11011011", "11011100", "11011100", "11011101", "11011101", "11011110", "11011111", "11011111", "11100000", "11100000", "11100001", "11100001", "11100010", "11100010", "11100011", "11100011", 
"11100011", "11100100", "11100100", "11100101", "11100101", "11100101", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101001", "11101001", "11101001", "11101001", "11101010", 
"11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", "11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101101", "11101110", "11101110", "11101110", 
"11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110001", "11110001", "11110001", 
"11110001", "11110001", "11110001", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", 
"00010001", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010010", "00010010", "00010011", "00010011", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", "00010100", "00010100", 
"00010101", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011010", "00011010", 
"00011010", "00011011", "00011011", "00011011", "00011100", "00011100", "00011101", "00011101", "00011101", "00011110", "00011110", "00011111", "00011111", "00100000", "00100000", "00100001", "00100001", "00100010", "00100011", "00100011", 
"00100100", "00100100", "00100101", "00100110", "00100111", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110001", "00110010", "00110011", "00110101", "00110110", 
"00110111", "00111001", "00111010", "00111100", "00111110", "00111111", "01000001", "01000011", "01000101", "01001000", "01001010", "01001100", "01001111", "01010001", "01010100", "01010111", "01011010", "10101001", "10101101", "10110001", 
"10110101", "10111010", "10111111", "11000100", "11001010", "11010001", "11011000", "11011111", "11100111", "11101111", "11111000", "00000000", "00001001", "00010010", "00011011", "00100011", "00101011", "00110010", "00111001", "00111111", 
"01000101", "01001010", "01001110", "01010011", "01010110", "01011010", "10101001", "10101100", "10101111", "10110010", "10110101", "10110111", "10111010", "10111100", "10111110", "11000000", "11000010", "11000100", "11000110", "11000111", 
"11001001", "11001010", "11001100", "11001101", "11001110", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011001", "11011010", "11011011", "11011100", "11011100", 
"11011101", "11011110", "11011110", "11011111", "11100000", "11100000", "11100001", "11100001", "11100010", "11100010", "11100011", "11100011", "11100100", "11100100", "11100100", "11100101", "11100101", "11100110", "11100110", "11100110", 
"11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101001", "11101001", "11101001", "11101010", "11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", 
"11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101101", "11101110", "11101110", "11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11110000", "11110000", 
"11110000", "11110000", "11110000", "11110000", "11110000", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "00001110", 
"00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", 
"00010000", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010010", "00010011", "00010011", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", 
"00010100", "00010100", "00010101", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", "00011010", 
"00011010", "00011010", "00011011", "00011011", "00011100", "00011100", "00011100", "00011101", "00011101", "00011110", "00011110", "00011111", "00011111", "00100000", "00100000", "00100001", "00100010", "00100010", "00100011", "00100100", 
"00100100", "00100101", "00100110", "00100111", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111", "00110000", "00110010", "00110011", "00110100", "00110110", "00110111", "00111001", 
"00111010", "00111100", "00111110", "01000000", "01000010", "01000100", "01000110", "01001001", "01001011", "01001110", "01010001", "01010100", "01010111", "01011010", "10101010", "10101101", "10110010", "10110110", "10111011", "11000001", 
"11000111", "11001110", "11010101", "11011101", "11100101", "11101110", "11110111", "00000000", "00001010", "00010011", "00011101", "00100101", "00101110", "00110101", "00111100", "01000011", "01001000", "01001101", "01010010", "01010110", 
"01011010", "10101010", "10101101", "10110000", "10110011", "10110110", "10111000", "10111011", "10111101", "10111111", "11000010", "11000100", "11000101", "11000111", "11001001", "11001011", "11001100", "11001110", "11001111", "11010000", 
"11010001", "11010011", "11010100", "11010101", "11010110", "11010111", "11011000", "11011001", "11011010", "11011010", "11011011", "11011100", "11011101", "11011101", "11011110", "11011111", "11011111", "11100000", "11100001", "11100001", 
"11100010", "11100010", "11100011", "11100011", "11100100", "11100100", "11100101", "11100101", "11100110", "11100110", "11100110", "11100111", "11100111", "11100111", "11101000", "11101000", "11101000", "11101001", "11101001", "11101001", 
"11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101101", "11101110", "11101110", "11101110", "11101110", 
"11101110", "11101111", "11101111", "11101111", "11101111", "11101111", "11101111", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", 
"11110001", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "00001101", "00001101", "00001101", "00001101", "00001101", 
"00001101", "00001101", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00010000", "00010000", 
"00010000", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010010", "00010011", "00010011", "00010011", "00010011", "00010011", 
"00010100", "00010100", "00010100", "00010100", "00010101", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", "00011001", "00011001", "00011001", 
"00011010", "00011010", "00011010", "00011011", "00011011", "00011100", "00011100", "00011101", "00011101", "00011110", "00011110", "00011111", "00011111", "00100000", "00100001", "00100001", "00100010", "00100011", "00100011", "00100100", 
"00100101", "00100110", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101111", "00110000", "00110001", "00110010", "00110100", "00110101", "00110111", "00111001", "00111011", "00111100", 
"00111110", "01000001", "01000011", "01000101", "01001000", "01001010", "01001101", "01010000", "01010011", "01010110", "01011010", "10101010", "10101110", "10110011", "10111000", "10111101", "11000100", "11001011", "11010010", "11011011", 
"11100011", "11101101", "11110110", "00000000", "00001011", "00010101", "00011111", "00101000", "00110001", "00111001", "01000000", "01000110", "01001100", "01010001", "01010110", "01011010", "10101010", "10101101", "10110001", "10110100", 
"10110111", "10111010", "10111100", "10111111", "11000001", "11000011", "11000101", "11000111", "11001001", "11001011", "11001100", "11001110", "11001111", "11010001", "11010010", "11010011", "11010101", "11010110", "11010111", "11011000", 
"11011001", "11011010", "11011011", "11011100", "11011100", "11011101", "11011110", "11011111", "11011111", "11100000", "11100001", "11100001", "11100010", "11100010", "11100011", "11100011", "11100100", "11100100", "11100101", "11100101", 
"11100110", "11100110", "11100111", "11100111", "11100111", "11101000", "11101000", "11101001", "11101001", "11101001", "11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", 
"11101100", "11101101", "11101101", "11101101", "11101101", "11101110", "11101110", "11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11101111", "11101111", "11110000", "11110000", "11110000", "11110000", "11110000", 
"11110000", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110011", "11110011", "11110011", "11110011", 
"11110011", "11110011", "11110011", "11110011", "11110011", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001101", "00001101", 
"00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", "00001111", 
"00001111", "00001111", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", "00010010", "00010011", "00010011", 
"00010011", "00010011", "00010100", "00010100", "00010100", "00010100", "00010101", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", "00011000", "00011000", "00011001", "00011001", 
"00011001", "00011010", "00011010", "00011011", "00011011", "00011100", "00011100", "00011101", "00011101", "00011110", "00011110", "00011111", "00011111", "00100000", "00100001", "00100001", "00100010", "00100011", "00100100", "00100100", 
"00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101101", "00101110", "00101111", "00110001", "00110010", "00110100", "00110101", "00110111", "00111001", "00111011", "00111101", "00111111", "01000001", 
"01000100", "01000110", "01001001", "01001100", "01001111", "01010011", "01010110", "01011010", "10101010", "10101111", "10110100", "10111010", "11000000", "11000111", "11001111", "11011000", "11100001", "11101011", "11110101", "00000000", 
"00001011", "00010111", "00100001", "00101011", "00110101", "00111101", "01000100", "01001011", "01010000", "01010101", "01011010", "10101010", "10101110", "10110010", "10110101", "10111000", "10111011", "10111110", "11000000", "11000011", 
"11000101", "11000111", "11001001", "11001011", "11001101", "11001111", "11010000", "11010010", "11010011", "11010100", "11010110", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011110", 
"11011111", "11100000", "11100001", "11100001", "11100010", "11100010", "11100011", "11100100", "11100100", "11100101", "11100101", "11100110", "11100110", "11100111", "11100111", "11101000", "11101000", "11101000", "11101001", "11101001", 
"11101001", "11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101110", "11101110", "11101110", "11101110", "11101110", "11101111", 
"11101111", "11101111", "11101111", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110001", "11110001", "11110001", "11110001", "11110001", "11110001", "11110010", "11110010", "11110010", "11110010", "11110010", 
"11110010", "11110010", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", 
"11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001100", "00001100", "00001100", "00001100", "00001100", 
"00001100", "00001100", "00001100", "00001100", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", 
"00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010010", 
"00010010", "00010011", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010111", "00010111", "00010111", "00011000", "00011000", "00011000", 
"00011001", "00011001", "00011010", "00011010", "00011011", "00011011", "00011100", "00011100", "00011101", "00011110", "00011110", "00011111", "00011111", "00100000", "00100001", "00100010", "00100010", "00100011", "00100100", "00100101", 
"00100110", "00100111", "00101000", "00101001", "00101010", "00101100", "00101101", "00101110", "00110000", "00110001", "00110011", "00110101", "00110111", "00111001", "00111011", "00111101", "01000000", "01000010", "01000101", "01001000", 
"01001011", "01001110", "01010010", "01010110", "01011010", "10101011", "10110000", "10110101", "10111100", "11000011", "11001011", "11010101", "11011111", "11101001", "11110101", "00000000", "00001101", "00011001", "00100100", "00101111", 
"00111001", "01000001", "01001001", "01001111", "01010101", "01011010", "10101011", "10101111", "10110011", "10110110", "10111010", "10111101", "11000000", "11000010", "11000101", "11000111", "11001001", "11001011", "11001101", "11001111", 
"11010001", "11010010", "11010100", "11010101", "11010111", "11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100000", "11100001", "11100010", "11100011", "11100011", "11100100", 
"11100100", "11100101", "11100110", "11100110", "11100111", "11100111", "11101000", "11101000", "11101000", "11101001", "11101001", "11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101100", "11101100", "11101100", 
"11101101", "11101101", "11101101", "11101110", "11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11101111", "11101111", "11110000", "11110000", "11110000", "11110000", "11110000", "11110001", "11110001", "11110001", 
"11110001", "11110001", "11110001", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110100", "11110100", "11110100", 
"11110100", "11110100", "11110100", "11110100", "11110100", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110110", "11110110", "11110110", "11110110", 
"11110110", "11110110", "11110110", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", 
"00001011", "00001011", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001110", "00001110", 
"00001110", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010001", "00010001", 
"00010010", "00010010", "00010010", "00010010", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010111", "00010111", "00011000", "00011000", 
"00011000", "00011001", "00011001", "00011010", "00011010", "00011011", "00011100", "00011100", "00011101", "00011101", "00011110", "00011111", "00100000", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100110", 
"00100111", "00101000", "00101001", "00101011", "00101100", "00101110", "00101111", "00110001", "00110011", "00110101", "00110111", "00111001", "00111011", "00111110", "01000000", "01000011", "01000110", "01001010", "01001101", "01010001", 
"01010101", "01011010", "10101011", "10110001", "10110111", "10111111", "11000111", "11010001", "11011100", "11100111", "11110011", "00000000", "00001110", "00011100", "00101000", "00110100", "00111110", "01000110", "01001110", "01010100", 
"01011010", "10101011", "10110000", "10110100", "10111000", "10111011", "10111111", "11000010", "11000101", "11000111", "11001010", "11001100", "11001110", "11010000", "11010010", "11010011", "11010101", "11010110", "11011000", "11011001", 
"11011010", "11011100", "11011101", "11011110", "11011111", "11100000", "11100000", "11100001", "11100010", "11100011", "11100011", "11100100", "11100101", "11100101", "11100110", "11100111", "11100111", "11101000", "11101000", "11101001", 
"11101001", "11101010", "11101010", "11101010", "11101011", "11101011", "11101011", "11101100", "11101100", "11101101", "11101101", "11101101", "11101101", "11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11101111", 
"11110000", "11110000", "11110000", "11110000", "11110000", "11110001", "11110001", "11110001", "11110001", "11110001", "11110010", "11110010", "11110010", "11110010", "11110010", "11110010", "11110011", "11110011", "11110011", "11110011", 
"11110011", "11110011", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", 
"11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "00001001", 
"00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001011", 
"00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001101", "00001101", "00001101", 
"00001101", "00001101", "00001101", "00001110", "00001110", "00001110", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010000", "00010000", "00010001", 
"00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010011", "00010011", "00010011", "00010011", "00010100", "00010100", "00010101", "00010101", "00010101", "00010110", "00010110", "00010110", "00010111", "00010111", 
"00011000", "00011000", "00011001", "00011001", "00011010", "00011011", "00011011", "00011100", "00011101", "00011101", "00011110", "00011111", "00100000", "00100000", "00100001", "00100010", "00100011", "00100100", "00100110", "00100111", 
"00101000", "00101010", "00101011", "00101101", "00101110", "00110000", "00110010", "00110100", "00110110", "00111001", "00111011", "00111110", "01000001", "01000101", "01001000", "01001100", "01010000", "01010101", "01011010", "10101100", 
"10110010", "10111010", "11000010", "11001100", "11011000", "11100100", "11110010", "00000000", "00010000", "00011111", "00101101", "00111001", "01000011", "01001100", "01010100", "01011010", "10101100", "10110001", "10110101", "10111010", 
"10111101", "11000001", "11000100", "11000111", "11001010", "11001100", "11001111", "11010001", "11010011", "11010101", "11010110", "11011000", "11011001", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", 
"11100010", "11100011", "11100100", "11100100", "11100101", "11100110", "11100110", "11100111", "11101000", "11101000", "11101001", "11101001", "11101010", "11101010", "11101011", "11101011", "11101100", "11101100", "11101100", "11101101", 
"11101101", "11101101", "11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11101111", "11110000", "11110000", "11110000", "11110000", "11110001", "11110001", "11110001", "11110001", "11110010", "11110010", "11110010", 
"11110010", "11110010", "11110011", "11110011", "11110011", "11110011", "11110011", "11110011", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", "11110101", "11110101", "11110101", "11110101", "11110101", 
"11110101", "11110101", "11110101", "11110101", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", 
"11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "00001000", "00001000", "00001000", "00001000", "00001000", 
"00001000", "00001000", "00001000", "00001000", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001010", "00001010", "00001010", 
"00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001100", "00001100", "00001100", "00001100", 
"00001100", "00001100", "00001100", "00001101", "00001101", "00001101", "00001101", "00001101", "00001101", "00001110", "00001110", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", "00010000", "00010000", 
"00010000", "00010000", "00010001", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010011", "00010011", "00010011", "00010100", "00010100", "00010100", "00010101", "00010101", "00010110", "00010110", "00010111", 
"00010111", "00011000", "00011000", "00011001", "00011010", "00011010", "00011011", "00011100", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011", "00100100", "00100101", "00100111", "00101000", 
"00101010", "00101011", "00101101", "00101111", "00110001", "00110100", "00110110", "00111001", "00111100", "00111111", "01000011", "01000110", "01001011", "01001111", "01010100", "01011010", "10101100", "10110100", "10111101", "11000111", 
"11010011", "11100001", "11110000", "00000000", "00010010", "00100011", "00110010", "00111111", "01001010", "01010011", "01011010", "10101100", "10110010", "10110111", "10111100", "11000000", "11000100", "11000111", "11001010", "11001101", 
"11010000", "11010010", "11010100", "11010110", "11011000", "11011001", "11011011", "11011100", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100110", "11100111", "11101000", 
"11101000", "11101001", "11101010", "11101010", "11101011", "11101011", "11101100", "11101100", "11101100", "11101101", "11101101", "11101110", "11101110", "11101110", "11101111", "11101111", "11101111", "11110000", "11110000", "11110000", 
"11110001", "11110001", "11110001", "11110001", "11110010", "11110010", "11110010", "11110010", "11110010", "11110011", "11110011", "11110011", "11110011", "11110011", "11110100", "11110100", "11110100", "11110100", "11110100", "11110100", 
"11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110111", "11110111", "11110111", 
"11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", 
"11111000", "11111000", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", 
"00000111", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001001", "00001001", "00001001", "00001001", "00001001", 
"00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001011", "00001011", "00001011", "00001011", "00001011", 
"00001011", "00001011", "00001011", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001101", "00001101", "00001101", "00001101", "00001101", "00001110", "00001110", "00001110", "00001110", "00001110", "00001111", 
"00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010001", "00010001", "00010001", "00010010", "00010010", "00010010", "00010011", "00010011", "00010100", "00010100", "00010100", "00010101", "00010101", "00010110", 
"00010110", "00010111", "00011000", "00011000", "00011001", "00011010", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100100", "00100101", "00100111", "00101000", "00101010", 
"00101100", "00101110", "00110000", "00110011", "00110110", "00111001", "00111100", "01000000", "01000100", "01001001", "01001110", "01010100", "01011010", "10101101", "10110110", "11000001", "11001110", "11011101", "11101110", "00000000", 
"00010101", "00101000", "00111001", "01000110", "01010001", "01011010", "10101101", "10110100", "10111010", "10111111", "11000011", "11000111", "11001011", "11001110", "11010001", "11010011", "11010110", "11011000", "11011010", "11011100", 
"11011101", "11011111", "11100000", "11100001", "11100010", "11100011", "11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101001", "11101010", "11101011", "11101011", "11101100", "11101100", "11101101", "11101101", 
"11101110", "11101110", "11101110", "11101111", "11101111", "11110000", "11110000", "11110000", "11110001", "11110001", "11110001", "11110001", "11110010", "11110010", "11110010", "11110010", "11110011", "11110011", "11110011", "11110011", 
"11110100", "11110100", "11110100", "11110100", "11110100", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110110", "11110111", 
"11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", 
"11111000", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111010", "11111010", "11111010", 
"11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000111", "00000111", 
"00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", 
"00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001010", "00001010", "00001010", "00001010", 
"00001010", "00001010", "00001010", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001100", "00001100", "00001100", "00001100", "00001100", "00001101", "00001101", "00001101", "00001101", "00001110", 
"00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00001111", "00010000", "00010000", "00010000", "00010001", "00010001", "00010010", "00010010", "00010010", "00010011", "00010011", "00010100", "00010100", "00010101", 
"00010101", "00010110", "00010111", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100011", "00100100", "00100110", "00101000", "00101010", "00101101", 
"00101111", "00110010", "00110101", "00111001", "00111101", "01000001", "01000110", "01001100", "01010011", "01011010", "10101111", "10111010", "11000111", "11011000", "11101011", "00000000", "00011001", "00101111", "01000001", "01001111", 
"01011010", "10101111", "10110110", "10111101", "11000010", "11000111", "11001011", "11001111", "11010010", "11010101", "11011000", "11011010", "11011100", "11011110", "11100000", "11100001", "11100011", "11100100", "11100101", "11100110", 
"11100111", "11101000", "11101001", "11101010", "11101010", "11101011", "11101100", "11101100", "11101101", "11101110", "11101110", "11101111", "11101111", "11101111", "11110000", "11110000", "11110001", "11110001", "11110001", "11110010", 
"11110010", "11110010", "11110011", "11110011", "11110011", "11110011", "11110100", "11110100", "11110100", "11110100", "11110101", "11110101", "11110101", "11110101", "11110101", "11110101", "11110110", "11110110", "11110110", "11110110", 
"11110110", "11110110", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", 
"11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", 
"11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", 
"11111011", "11111011", "11111011", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000110", "00000110", "00000110", "00000110", 
"00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", 
"00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001001", "00001001", "00001001", 
"00001001", "00001001", "00001001", "00001001", "00001001", "00001010", "00001010", "00001010", "00001010", "00001010", "00001010", "00001011", "00001011", "00001011", "00001011", "00001011", "00001011", "00001100", "00001100", "00001100", 
"00001100", "00001101", "00001101", "00001101", "00001101", "00001110", "00001110", "00001110", "00001111", "00001111", "00001111", "00010000", "00010000", "00010001", "00010001", "00010001", "00010010", "00010010", "00010011", "00010100", 
"00010100", "00010101", "00010110", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011111", "00100000", "00100010", "00100100", "00100110", "00101000", "00101011", "00101110", "00110001", 
"00110101", "00111001", "00111110", "01000011", "01001010", "01010001", "01011010", "10110001", "10111111", "11010001", "11100111", "00000000", "00011111", "00111001", "01001100", "01011010", "10110001", "10111010", "11000001", "11000111", 
"11001100", "11010001", "11010101", "11011000", "11011011", "11011101", "11011111", "11100001", "11100011", "11100100", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101101", "11101110", 
"11101111", "11101111", "11110000", "11110000", "11110001", "11110001", "11110010", "11110010", "11110010", "11110011", "11110011", "11110011", "11110100", "11110100", "11110100", "11110101", "11110101", "11110101", "11110101", "11110101", 
"11110110", "11110110", "11110110", "11110110", "11110110", "11110111", "11110111", "11110111", "11110111", "11110111", "11110111", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111001", 
"11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", 
"11111010", "11111010", "11111010", "11111010", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", 
"11111011", "11111011", "11111011", "11111011", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "00000100", 
"00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000101", "00000101", "00000101", "00000101", "00000101", 
"00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000110", "00000110", "00000110", "00000110", "00000110", 
"00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", 
"00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001001", "00001001", "00001001", "00001001", "00001001", "00001001", "00001010", "00001010", "00001010", "00001010", "00001010", "00001011", 
"00001011", "00001011", "00001011", "00001011", "00001100", "00001100", "00001100", "00001101", "00001101", "00001101", "00001110", "00001110", "00001110", "00001111", "00001111", "00010000", "00010000", "00010001", "00010001", "00010010", 
"00010011", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011100", "00011101", "00011111", "00100001", "00100011", "00100101", "00101000", "00101011", "00101111", "00110100", "00111001", 
"00111111", "01000110", "01001111", "01011010", "10110100", "11000111", "11100001", "00000000", "00101000", "01000110", "01011010", "10110100", "10111111", "11000111", "11001110", "11010011", "11011000", "11011100", "11011111", "11100001", 
"11100011", "11100101", "11100111", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111", "11110000", "11110000", "11110001", "11110001", "11110010", "11110010", "11110011", "11110011", "11110100", "11110100", 
"11110101", "11110101", "11110101", "11110101", "11110110", "11110110", "11110110", "11110111", "11110111", "11110111", "11110111", "11110111", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111001", "11111001", 
"11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111011", "11111011", "11111011", 
"11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", 
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111101", "11111101", "11111101", "11111101", 
"11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "00000011", "00000011", "00000011", "00000011", "00000011", 
"00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000100", "00000100", "00000100", "00000100", "00000100", 
"00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000101", 
"00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", 
"00000110", "00000110", "00000110", "00000110", "00000110", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00001000", "00001000", "00001000", "00001000", "00001000", "00001000", "00001001", 
"00001001", "00001001", "00001001", "00001001", "00001010", "00001010", "00001010", "00001011", "00001011", "00001011", "00001011", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111", "00001111", "00010000", 
"00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011001", "00011011", "00011101", "00011111", "00100001", "00100100", "00101000", "00101101", "00110010", "00111001", "01000001", "01001100", 
"01011010", "10111010", "11011000", "00000000", "00111001", "01011010", "10111010", "11000111", "11010001", "11011000", "11011101", "11100001", "11100100", "11100111", "11101001", "11101011", "11101101", "11101110", "11101111", "11110000", 
"11110001", "11110010", "11110011", "11110011", "11110100", "11110101", "11110101", "11110101", "11110110", "11110110", "11110111", "11110111", "11110111", "11111000", "11111000", "11111000", "11111000", "11111001", "11111001", "11111001", 
"11111001", "11111001", "11111001", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111010", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", "11111011", 
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111101", "11111101", "11111101", "11111101", 
"11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", 
"11111101", "11111101", "11111101", "11111101", "11111101", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", 
"11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", 
"00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000011", "00000011", 
"00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", 
"00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", 
"00000100", "00000100", "00000100", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000101", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", 
"00000111", "00000111", "00000111", "00000111", "00000111", "00000111", "00001000", "00001000", "00001000", "00001000", "00001001", "00001001", "00001001", "00001010", "00001010", "00001011", "00001011", "00001011", "00001100", "00001101", 
"00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010101", "00010111", "00011001", "00011100", "00011111", "00100011", "00101000", "00101111", "00111001", "01000110", "01011010", "11000111", "00000000", 
"01011010", "11000111", "11011000", "11100001", "11100111", "11101011", "11101110", "11110000", "11110010", "11110011", "11110101", "11110101", "11110110", "11110111", "11111000", "11111000", "11111001", "11111001", "11111001", "11111010", 
"11111010", "11111010", "11111010", "11111011", "11111011", "11111011", "11111011", "11111011", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111101", "11111101", "11111101", "11111101", 
"11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111101", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", 
"11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", "11111110", 
"11111110", "11111110", "11111110", "11111110", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", 
"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", 
"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", 
"00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", 
"00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000001", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", 
"00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", "00000010", 
"00000010", "00000010", "00000010", "00000010", "00000010", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000100", 
"00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000100", "00000101", "00000101", "00000101", "00000101", "00000101", "00000110", "00000110", "00000110", "00000110", "00000111", "00000111", "00000111", "00001000", 
"00001000", "00001001", "00001010", "00001011", "00001011", "00001101", "00001110", "00010000", "00010010", "00010101", "00011001", "00011111", "00101000", "00111001", "01011010" );
begin
process(clk) is
begin
	if rising_edge(clk) then
		if i_ce='1' then
			sample_out_re<=mem_re(conv_integer(sample_in_im&sample_in_re));
			sample_out_im<=mem_im(conv_integer(sample_in_im&sample_in_re));
		end if;
		o_ce<=i_ce;
	end if;
end process;
end table_demod;
