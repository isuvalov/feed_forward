--
--  Copyright (c) 2003 Launchbird Design Systems, Inc.
--  All rights reserved.
--  
--  Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
--    Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
--    Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES,
--  INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
--  IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--  OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
--  OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--  (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--  
--  Overview:
--  
--    Cordics (COordinate Rotation DIgital Computers) are used to calculate
--    trigonometric functions and complex plane phase rotations.
--    This vector mode cordic rotates any complex vector to the positive real axis.
--    The resulting angle is the initial angle plus the angle of rotation.
--  
--  Interface:
--  
--    Synchronization:
--      clock_c  : Clock input.
--      enable_i : Synchronous enable.
--      reset_i  : Synchronous reset.
--  
--    Inputs:
--      real_i   : Initial real component (signed).
--      imag_i   : Initial imaginary component (signed).
--      angle_i  : Initial angle (modulo 2PI).
--  
--    Outputs:
--      real_o   : Resulting real component (signed).
--      imag_o   : Resulting imaginary component (signed).
--      angle_o  : Resulting angle (modulo 2PI).
--  
--  Built In Parameters:
--  
--    Cordic Mode    = Vector
--    Vector Width   = 32
--    Angle Width    = 32
--    Cordic Stages  = 32
--  
--  Resulting Pipeline Latency is 34 clock cycles.
--  
--  
--  
--  Generated by Confluence 0.6.3  --  Launchbird Design Systems, Inc.  --  www.launchbird.com
--  
--  Build Date : Fri Aug 22 09:44:40 CDT 2003
--  
--  Interface
--  
--    Build Name    : cf_cordic_v_32_32_32
--    Clock Domains : clock_c  
--    Vector Input  : enable_i(1)
--    Vector Input  : reset_i(1)
--    Vector Input  : real_i(32)
--    Vector Input  : imag_i(32)
--    Vector Input  : ang_i(32)
--    Vector Output : real_o(32)
--    Vector Output : imag_o(32)
--    Vector Output : ang_o(32)
--  
--  
--  

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_cordic_v_32_32_32_56;
architecture rtl of cf_cordic_v_32_32_32_56 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(30 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(32 downto 0);
signal n7 : unsigned(32 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(32 downto 0);
begin
n1 <= i1(31 downto 31);
n2 <= not n1;
n3 <= i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n4 <= n2 & n3;
n5 <= "0";
n6 <= n5 & n4;
n7 <= n9 - n6;
n8 <= n7(32 downto 32);
n9 <= "010000000000000000000000000000000";
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_55 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_55;
architecture rtl of cf_cordic_v_32_32_32_55 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(29 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(1 downto 0);
signal n12 : unsigned(29 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s23_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & n1;
n3 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3) &
  i4(2 downto 2);
n4 <= n2 & n3;
n5 <= i3 + n4;
n6 <= i3 - n4;
n7 <= n5 when s23_1 = "1" else n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n8 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
n9 <= not s23_1;
n10 <= i3(31 downto 31);
n11 <= n10 & n10;
n12 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2);
n13 <= n11 & n12;
n14 <= i4 + n13;
n15 <= i4 - n13;
n16 <= n14 when n9 = "1" else n15;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n17 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n17 <= n16;
    end if;
  end if;
end process;
n18 <= "00001001111110110011100001011011";
n19 <= i5 + n18;
n20 <= i5 - n18;
n21 <= n19 when s23_1 = "1" else n20;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n22 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n22 <= n21;
    end if;
  end if;
end process;
s23 : cf_cordic_v_32_32_32_56 port map (i4, s23_1);
o3 <= n22;
o2 <= n17;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end entity cf_cordic_v_32_32_32_54;
architecture rtl of cf_cordic_v_32_32_32_54 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(4 downto 0);
signal n5 : unsigned(5 downto 0);
signal n6 : unsigned(6 downto 0);
signal n7 : unsigned(7 downto 0);
signal n8 : unsigned(8 downto 0);
begin
n1 <= i1 & i1;
n2 <= i1 & n1;
n3 <= i1 & n2;
n4 <= i1 & n3;
n5 <= i1 & n4;
n6 <= i1 & n5;
n7 <= i1 & n6;
n8 <= i1 & n7;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_53 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_53;
architecture rtl of cf_cordic_v_32_32_32_53 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(22 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(22 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s21_1 : unsigned(8 downto 0);
signal s22_1 : unsigned(8 downto 0);
signal s23_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_v_32_32_32_54;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9);
n3 <= s21_1 & n2;
n4 <= i3 + n3;
n5 <= i3 - n3;
n6 <= n4 when s23_1 = "1" else n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= not s23_1;
n9 <= i3(31 downto 31);
n10 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9);
n11 <= s22_1 & n10;
n12 <= i4 + n11;
n13 <= i4 - n11;
n14 <= n12 when n8 = "1" else n13;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n15 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
n16 <= "00000000000101000101111100101111";
n17 <= i5 + n16;
n18 <= i5 - n16;
n19 <= n17 when s23_1 = "1" else n18;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n20 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n20 <= n19;
    end if;
  end if;
end process;
s21 : cf_cordic_v_32_32_32_54 port map (n1, s21_1);
s22 : cf_cordic_v_32_32_32_54 port map (n9, s22_1);
s23 : cf_cordic_v_32_32_32_56 port map (i4, s23_1);
o3 <= n20;
o2 <= n15;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_cordic_v_32_32_32_52;
architecture rtl of cf_cordic_v_32_32_32_52 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(10 downto 0);
signal n3 : unsigned(11 downto 0);
signal n4 : unsigned(12 downto 0);
signal n5 : unsigned(13 downto 0);
signal n6 : unsigned(14 downto 0);
signal n7 : unsigned(15 downto 0);
signal s8_1 : unsigned(8 downto 0);
component cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_v_32_32_32_54;
begin
n1 <= i1 & s8_1;
n2 <= i1 & n1;
n3 <= i1 & n2;
n4 <= i1 & n3;
n5 <= i1 & n4;
n6 <= i1 & n5;
n7 <= i1 & n6;
s8 : cf_cordic_v_32_32_32_54 port map (i1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_51 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_51;
architecture rtl of cf_cordic_v_32_32_32_51 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s21_1 : unsigned(15 downto 0);
signal s22_1 : unsigned(15 downto 0);
signal s23_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_v_32_32_32_52;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16);
n3 <= s21_1 & n2;
n4 <= i3 + n3;
n5 <= i3 - n3;
n6 <= n4 when s23_1 = "1" else n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= not s23_1;
n9 <= i3(31 downto 31);
n10 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16);
n11 <= s22_1 & n10;
n12 <= i4 + n11;
n13 <= i4 - n11;
n14 <= n12 when n8 = "1" else n13;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n15 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
n16 <= "00000000000000000010100010111110";
n17 <= i5 + n16;
n18 <= i5 - n16;
n19 <= n17 when s23_1 = "1" else n18;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n20 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n20 <= n19;
    end if;
  end if;
end process;
s21 : cf_cordic_v_32_32_32_52 port map (n1, s21_1);
s22 : cf_cordic_v_32_32_32_52 port map (n9, s22_1);
s23 : cf_cordic_v_32_32_32_56 port map (i4, s23_1);
o3 <= n20;
o2 <= n15;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end entity cf_cordic_v_32_32_32_50;
architecture rtl of cf_cordic_v_32_32_32_50 is
signal n1 : unsigned(16 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(18 downto 0);
signal n4 : unsigned(19 downto 0);
signal n5 : unsigned(20 downto 0);
signal n6 : unsigned(21 downto 0);
signal n7 : unsigned(22 downto 0);
signal s8_1 : unsigned(15 downto 0);
component cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_v_32_32_32_52;
begin
n1 <= i1 & s8_1;
n2 <= i1 & n1;
n3 <= i1 & n2;
n4 <= i1 & n3;
n5 <= i1 & n4;
n6 <= i1 & n5;
n7 <= i1 & n6;
s8 : cf_cordic_v_32_32_32_52 port map (i1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_49 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_49;
architecture rtl of cf_cordic_v_32_32_32_49 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(8 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s21_1 : unsigned(22 downto 0);
signal s22_1 : unsigned(22 downto 0);
signal s23_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_cordic_v_32_32_32_50;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23);
n3 <= s21_1 & n2;
n4 <= i3 + n3;
n5 <= i3 - n3;
n6 <= n4 when s23_1 = "1" else n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= not s23_1;
n9 <= i3(31 downto 31);
n10 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23);
n11 <= s22_1 & n10;
n12 <= i4 + n11;
n13 <= i4 - n11;
n14 <= n12 when n8 = "1" else n13;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n15 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
n16 <= "00000000000000000000000001010001";
n17 <= i5 + n16;
n18 <= i5 - n16;
n19 <= n17 when s23_1 = "1" else n18;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n20 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n20 <= n19;
    end if;
  end if;
end process;
s21 : cf_cordic_v_32_32_32_50 port map (n1, s21_1);
s22 : cf_cordic_v_32_32_32_50 port map (n9, s22_1);
s23 : cf_cordic_v_32_32_32_56 port map (i4, s23_1);
o3 <= n20;
o2 <= n15;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_48 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(29 downto 0));
end entity cf_cordic_v_32_32_32_48;
architecture rtl of cf_cordic_v_32_32_32_48 is
signal n1 : unsigned(23 downto 0);
signal n2 : unsigned(24 downto 0);
signal n3 : unsigned(25 downto 0);
signal n4 : unsigned(26 downto 0);
signal n5 : unsigned(27 downto 0);
signal n6 : unsigned(28 downto 0);
signal n7 : unsigned(29 downto 0);
signal s8_1 : unsigned(22 downto 0);
component cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_cordic_v_32_32_32_50;
begin
n1 <= i1 & s8_1;
n2 <= i1 & n1;
n3 <= i1 & n2;
n4 <= i1 & n3;
n5 <= i1 & n4;
n6 <= i1 & n5;
n7 <= i1 & n6;
s8 : cf_cordic_v_32_32_32_50 port map (i1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_47 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_47;
architecture rtl of cf_cordic_v_32_32_32_47 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(30 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(30 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s23_1 : unsigned(29 downto 0);
signal s24_1 : unsigned(29 downto 0);
signal s25_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_48 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(29 downto 0));
end component cf_cordic_v_32_32_32_48;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s23_1;
n3 <= i4(31 downto 31);
n4 <= n2 & n3;
n5 <= i3 + n4;
n6 <= i3 - n4;
n7 <= n5 when s25_1 = "1" else n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n8 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
n9 <= not s25_1;
n10 <= i3(31 downto 31);
n11 <= n10 & s24_1;
n12 <= i3(31 downto 31);
n13 <= n11 & n12;
n14 <= i4 + n13;
n15 <= i4 - n13;
n16 <= n14 when n9 = "1" else n15;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n17 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n17 <= n16;
    end if;
  end if;
end process;
n18 <= "00000000000000000000000000000000";
n19 <= i5 + n18;
n20 <= i5 - n18;
n21 <= n19 when s25_1 = "1" else n20;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n22 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n22 <= n21;
    end if;
  end if;
end process;
s23 : cf_cordic_v_32_32_32_48 port map (n1, s23_1);
s24 : cf_cordic_v_32_32_32_48 port map (n10, s24_1);
s25 : cf_cordic_v_32_32_32_56 port map (i4, s25_1);
o3 <= n22;
o2 <= n17;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_46 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_46;
architecture rtl of cf_cordic_v_32_32_32_46 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(1 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s21_1 : unsigned(29 downto 0);
signal s22_1 : unsigned(29 downto 0);
signal s23_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_48 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(29 downto 0));
end component cf_cordic_v_32_32_32_48;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= i4(31 downto 31) &
  i4(30 downto 30);
n3 <= s21_1 & n2;
n4 <= i3 + n3;
n5 <= i3 - n3;
n6 <= n4 when s23_1 = "1" else n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= not s23_1;
n9 <= i3(31 downto 31);
n10 <= i3(31 downto 31) &
  i3(30 downto 30);
n11 <= s22_1 & n10;
n12 <= i4 + n11;
n13 <= i4 - n11;
n14 <= n12 when n8 = "1" else n13;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n15 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
n16 <= "00000000000000000000000000000001";
n17 <= i5 + n16;
n18 <= i5 - n16;
n19 <= n17 when s23_1 = "1" else n18;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n20 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n20 <= n19;
    end if;
  end if;
end process;
s21 : cf_cordic_v_32_32_32_48 port map (n1, s21_1);
s22 : cf_cordic_v_32_32_32_48 port map (n9, s22_1);
s23 : cf_cordic_v_32_32_32_56 port map (i4, s23_1);
o3 <= n20;
o2 <= n15;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_45 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_45;
architecture rtl of cf_cordic_v_32_32_32_45 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(23 downto 0);
signal n3 : unsigned(24 downto 0);
signal n4 : unsigned(25 downto 0);
signal n5 : unsigned(26 downto 0);
signal n6 : unsigned(27 downto 0);
signal n7 : unsigned(28 downto 0);
signal n8 : unsigned(2 downto 0);
signal n9 : unsigned(31 downto 0);
signal s10_1 : unsigned(22 downto 0);
component cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_cordic_v_32_32_32_50;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s10_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= n1 & n6;
n8 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29);
n9 <= n7 & n8;
s10 : cf_cordic_v_32_32_32_50 port map (n1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_44 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_44;
architecture rtl of cf_cordic_v_32_32_32_44 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_45 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_45;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000000000000000000001";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_45 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_45 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_43 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_43;
architecture rtl of cf_cordic_v_32_32_32_43 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(23 downto 0);
signal n3 : unsigned(24 downto 0);
signal n4 : unsigned(25 downto 0);
signal n5 : unsigned(26 downto 0);
signal n6 : unsigned(27 downto 0);
signal n7 : unsigned(3 downto 0);
signal n8 : unsigned(31 downto 0);
signal s9_1 : unsigned(22 downto 0);
component cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_cordic_v_32_32_32_50;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s9_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28);
n8 <= n6 & n7;
s9 : cf_cordic_v_32_32_32_50 port map (n1, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_42 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_42;
architecture rtl of cf_cordic_v_32_32_32_42 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_43 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_43;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000000000000000000011";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_43 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_43 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_41 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_41;
architecture rtl of cf_cordic_v_32_32_32_41 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(23 downto 0);
signal n3 : unsigned(24 downto 0);
signal n4 : unsigned(25 downto 0);
signal n5 : unsigned(26 downto 0);
signal n6 : unsigned(4 downto 0);
signal n7 : unsigned(31 downto 0);
signal s8_1 : unsigned(22 downto 0);
component cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_cordic_v_32_32_32_50;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s8_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27);
n7 <= n5 & n6;
s8 : cf_cordic_v_32_32_32_50 port map (n1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_40 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_40;
architecture rtl of cf_cordic_v_32_32_32_40 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_41 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_41;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000000000000000000101";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_41 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_41 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_39 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_39;
architecture rtl of cf_cordic_v_32_32_32_39 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(23 downto 0);
signal n3 : unsigned(24 downto 0);
signal n4 : unsigned(25 downto 0);
signal n5 : unsigned(5 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0);
signal n10 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(23 downto 0);
signal n14 : unsigned(24 downto 0);
signal n15 : unsigned(25 downto 0);
signal n16 : unsigned(5 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s27_1 : unsigned(22 downto 0);
signal s28_1 : unsigned(22 downto 0);
signal s29_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_cordic_v_32_32_32_50;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s27_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26);
n6 <= n4 & n5;
n7 <= i3 + n6;
n8 <= i3 - n6;
n9 <= n7 when s29_1 = "1" else n8;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n10 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
n11 <= not s29_1;
n12 <= i3(31 downto 31);
n13 <= n12 & s28_1;
n14 <= n12 & n13;
n15 <= n12 & n14;
n16 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26);
n17 <= n15 & n16;
n18 <= i4 + n17;
n19 <= i4 - n17;
n20 <= n18 when n11 = "1" else n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n21 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= "00000000000000000000000000001010";
n23 <= i5 + n22;
n24 <= i5 - n22;
n25 <= n23 when s29_1 = "1" else n24;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n26 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n26 <= n25;
    end if;
  end if;
end process;
s27 : cf_cordic_v_32_32_32_50 port map (n1, s27_1);
s28 : cf_cordic_v_32_32_32_50 port map (n12, s28_1);
s29 : cf_cordic_v_32_32_32_56 port map (i4, s29_1);
o3 <= n26;
o2 <= n21;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_38 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_38;
architecture rtl of cf_cordic_v_32_32_32_38 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(23 downto 0);
signal n3 : unsigned(24 downto 0);
signal n4 : unsigned(6 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(23 downto 0);
signal n13 : unsigned(24 downto 0);
signal n14 : unsigned(6 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s25_1 : unsigned(22 downto 0);
signal s26_1 : unsigned(22 downto 0);
signal s27_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_cordic_v_32_32_32_50;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s25_1;
n3 <= n1 & n2;
n4 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25);
n5 <= n3 & n4;
n6 <= i3 + n5;
n7 <= i3 - n5;
n8 <= n6 when s27_1 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= not s27_1;
n11 <= i3(31 downto 31);
n12 <= n11 & s26_1;
n13 <= n11 & n12;
n14 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25);
n15 <= n13 & n14;
n16 <= i4 + n15;
n17 <= i4 - n15;
n18 <= n16 when n10 = "1" else n17;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n19 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= "00000000000000000000000000010100";
n21 <= i5 + n20;
n22 <= i5 - n20;
n23 <= n21 when s27_1 = "1" else n22;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n24 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
s25 : cf_cordic_v_32_32_32_50 port map (n1, s25_1);
s26 : cf_cordic_v_32_32_32_50 port map (n11, s26_1);
s27 : cf_cordic_v_32_32_32_56 port map (i4, s27_1);
o3 <= n24;
o2 <= n19;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_37;
architecture rtl of cf_cordic_v_32_32_32_37 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(23 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(23 downto 0);
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s23_1 : unsigned(22 downto 0);
signal s24_1 : unsigned(22 downto 0);
signal s25_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_50 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_cordic_v_32_32_32_50;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s23_1;
n3 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24);
n4 <= n2 & n3;
n5 <= i3 + n4;
n6 <= i3 - n4;
n7 <= n5 when s25_1 = "1" else n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n8 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
n9 <= not s25_1;
n10 <= i3(31 downto 31);
n11 <= n10 & s24_1;
n12 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24);
n13 <= n11 & n12;
n14 <= i4 + n13;
n15 <= i4 - n13;
n16 <= n14 when n9 = "1" else n15;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n17 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n17 <= n16;
    end if;
  end if;
end process;
n18 <= "00000000000000000000000000101001";
n19 <= i5 + n18;
n20 <= i5 - n18;
n21 <= n19 when s25_1 = "1" else n20;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n22 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n22 <= n21;
    end if;
  end if;
end process;
s23 : cf_cordic_v_32_32_32_50 port map (n1, s23_1);
s24 : cf_cordic_v_32_32_32_50 port map (n10, s24_1);
s25 : cf_cordic_v_32_32_32_56 port map (i4, s25_1);
o3 <= n22;
o2 <= n17;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_36 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_36;
architecture rtl of cf_cordic_v_32_32_32_36 is
signal s1_1 : unsigned(31 downto 0);
signal s1_2 : unsigned(31 downto 0);
signal s1_3 : unsigned(31 downto 0);
signal s2_1 : unsigned(31 downto 0);
signal s2_2 : unsigned(31 downto 0);
signal s2_3 : unsigned(31 downto 0);
signal s3_1 : unsigned(31 downto 0);
signal s3_2 : unsigned(31 downto 0);
signal s3_3 : unsigned(31 downto 0);
signal s4_1 : unsigned(31 downto 0);
signal s4_2 : unsigned(31 downto 0);
signal s4_3 : unsigned(31 downto 0);
signal s5_1 : unsigned(31 downto 0);
signal s5_2 : unsigned(31 downto 0);
signal s5_3 : unsigned(31 downto 0);
signal s6_1 : unsigned(31 downto 0);
signal s6_2 : unsigned(31 downto 0);
signal s6_3 : unsigned(31 downto 0);
signal s7_1 : unsigned(31 downto 0);
signal s7_2 : unsigned(31 downto 0);
signal s7_3 : unsigned(31 downto 0);
signal s8_1 : unsigned(31 downto 0);
signal s8_2 : unsigned(31 downto 0);
signal s8_3 : unsigned(31 downto 0);
component cf_cordic_v_32_32_32_47 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_47;
component cf_cordic_v_32_32_32_46 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_46;
component cf_cordic_v_32_32_32_44 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_44;
component cf_cordic_v_32_32_32_42 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_42;
component cf_cordic_v_32_32_32_40 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_40;
component cf_cordic_v_32_32_32_39 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_39;
component cf_cordic_v_32_32_32_38 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_38;
component cf_cordic_v_32_32_32_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_37;
begin
s1 : cf_cordic_v_32_32_32_47 port map (clock_c, i1, i2, s2_1, s2_2, s2_3, s1_1, s1_2, s1_3);
s2 : cf_cordic_v_32_32_32_46 port map (clock_c, i1, i2, s3_1, s3_2, s3_3, s2_1, s2_2, s2_3);
s3 : cf_cordic_v_32_32_32_44 port map (clock_c, i1, i2, s4_1, s4_2, s4_3, s3_1, s3_2, s3_3);
s4 : cf_cordic_v_32_32_32_42 port map (clock_c, i1, i2, s5_1, s5_2, s5_3, s4_1, s4_2, s4_3);
s5 : cf_cordic_v_32_32_32_40 port map (clock_c, i1, i2, s6_1, s6_2, s6_3, s5_1, s5_2, s5_3);
s6 : cf_cordic_v_32_32_32_39 port map (clock_c, i1, i2, s7_1, s7_2, s7_3, s6_1, s6_2, s6_3);
s7 : cf_cordic_v_32_32_32_38 port map (clock_c, i1, i2, s8_1, s8_2, s8_3, s7_1, s7_2, s7_3);
s8 : cf_cordic_v_32_32_32_37 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s1_3;
o2 <= s1_2;
o1 <= s1_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_35 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_35;
architecture rtl of cf_cordic_v_32_32_32_35 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(16 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(18 downto 0);
signal n5 : unsigned(19 downto 0);
signal n6 : unsigned(20 downto 0);
signal n7 : unsigned(21 downto 0);
signal n8 : unsigned(9 downto 0);
signal n9 : unsigned(31 downto 0);
signal s10_1 : unsigned(15 downto 0);
component cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_v_32_32_32_52;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s10_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= n1 & n6;
n8 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22);
n9 <= n7 & n8;
s10 : cf_cordic_v_32_32_32_52 port map (n1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_34 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_34;
architecture rtl of cf_cordic_v_32_32_32_34 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_35 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_35;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000000000000010100011";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_35 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_35 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_33 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_33;
architecture rtl of cf_cordic_v_32_32_32_33 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(16 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(18 downto 0);
signal n5 : unsigned(19 downto 0);
signal n6 : unsigned(20 downto 0);
signal n7 : unsigned(10 downto 0);
signal n8 : unsigned(31 downto 0);
signal s9_1 : unsigned(15 downto 0);
component cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_v_32_32_32_52;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s9_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21);
n8 <= n6 & n7;
s9 : cf_cordic_v_32_32_32_52 port map (n1, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_32;
architecture rtl of cf_cordic_v_32_32_32_32 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_33 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_33;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000000000000101000110";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_33 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_33 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_31 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_31;
architecture rtl of cf_cordic_v_32_32_32_31 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(16 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(18 downto 0);
signal n5 : unsigned(19 downto 0);
signal n6 : unsigned(11 downto 0);
signal n7 : unsigned(31 downto 0);
signal s8_1 : unsigned(15 downto 0);
component cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_v_32_32_32_52;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s8_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20);
n7 <= n5 & n6;
s8 : cf_cordic_v_32_32_32_52 port map (n1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_30;
architecture rtl of cf_cordic_v_32_32_32_30 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_31 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_31;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000000000001010001100";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_31 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_31 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_29 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_29;
architecture rtl of cf_cordic_v_32_32_32_29 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(16 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(18 downto 0);
signal n5 : unsigned(12 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0);
signal n10 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(16 downto 0);
signal n14 : unsigned(17 downto 0);
signal n15 : unsigned(18 downto 0);
signal n16 : unsigned(12 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s27_1 : unsigned(15 downto 0);
signal s28_1 : unsigned(15 downto 0);
signal s29_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_v_32_32_32_52;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s27_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19);
n6 <= n4 & n5;
n7 <= i3 + n6;
n8 <= i3 - n6;
n9 <= n7 when s29_1 = "1" else n8;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n10 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
n11 <= not s29_1;
n12 <= i3(31 downto 31);
n13 <= n12 & s28_1;
n14 <= n12 & n13;
n15 <= n12 & n14;
n16 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19);
n17 <= n15 & n16;
n18 <= i4 + n17;
n19 <= i4 - n17;
n20 <= n18 when n11 = "1" else n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n21 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= "00000000000000000000010100011000";
n23 <= i5 + n22;
n24 <= i5 - n22;
n25 <= n23 when s29_1 = "1" else n24;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n26 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n26 <= n25;
    end if;
  end if;
end process;
s27 : cf_cordic_v_32_32_32_52 port map (n1, s27_1);
s28 : cf_cordic_v_32_32_32_52 port map (n12, s28_1);
s29 : cf_cordic_v_32_32_32_56 port map (i4, s29_1);
o3 <= n26;
o2 <= n21;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_28;
architecture rtl of cf_cordic_v_32_32_32_28 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(16 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(13 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(16 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(13 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s25_1 : unsigned(15 downto 0);
signal s26_1 : unsigned(15 downto 0);
signal s27_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_v_32_32_32_52;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s25_1;
n3 <= n1 & n2;
n4 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18);
n5 <= n3 & n4;
n6 <= i3 + n5;
n7 <= i3 - n5;
n8 <= n6 when s27_1 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= not s27_1;
n11 <= i3(31 downto 31);
n12 <= n11 & s26_1;
n13 <= n11 & n12;
n14 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18);
n15 <= n13 & n14;
n16 <= i4 + n15;
n17 <= i4 - n15;
n18 <= n16 when n10 = "1" else n17;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n19 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= "00000000000000000000101000110000";
n21 <= i5 + n20;
n22 <= i5 - n20;
n23 <= n21 when s27_1 = "1" else n22;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n24 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
s25 : cf_cordic_v_32_32_32_52 port map (n1, s25_1);
s26 : cf_cordic_v_32_32_32_52 port map (n11, s26_1);
s27 : cf_cordic_v_32_32_32_56 port map (i4, s27_1);
o3 <= n24;
o2 <= n19;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_27;
architecture rtl of cf_cordic_v_32_32_32_27 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(16 downto 0);
signal n3 : unsigned(14 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(16 downto 0);
signal n12 : unsigned(14 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s23_1 : unsigned(15 downto 0);
signal s24_1 : unsigned(15 downto 0);
signal s25_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_52 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_cordic_v_32_32_32_52;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s23_1;
n3 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17);
n4 <= n2 & n3;
n5 <= i3 + n4;
n6 <= i3 - n4;
n7 <= n5 when s25_1 = "1" else n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n8 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
n9 <= not s25_1;
n10 <= i3(31 downto 31);
n11 <= n10 & s24_1;
n12 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17);
n13 <= n11 & n12;
n14 <= i4 + n13;
n15 <= i4 - n13;
n16 <= n14 when n9 = "1" else n15;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n17 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n17 <= n16;
    end if;
  end if;
end process;
n18 <= "00000000000000000001010001011111";
n19 <= i5 + n18;
n20 <= i5 - n18;
n21 <= n19 when s25_1 = "1" else n20;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n22 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n22 <= n21;
    end if;
  end if;
end process;
s23 : cf_cordic_v_32_32_32_52 port map (n1, s23_1);
s24 : cf_cordic_v_32_32_32_52 port map (n10, s24_1);
s25 : cf_cordic_v_32_32_32_56 port map (i4, s25_1);
o3 <= n22;
o2 <= n17;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_26;
architecture rtl of cf_cordic_v_32_32_32_26 is
signal s1_1 : unsigned(31 downto 0);
signal s1_2 : unsigned(31 downto 0);
signal s1_3 : unsigned(31 downto 0);
signal s2_1 : unsigned(31 downto 0);
signal s2_2 : unsigned(31 downto 0);
signal s2_3 : unsigned(31 downto 0);
signal s3_1 : unsigned(31 downto 0);
signal s3_2 : unsigned(31 downto 0);
signal s3_3 : unsigned(31 downto 0);
signal s4_1 : unsigned(31 downto 0);
signal s4_2 : unsigned(31 downto 0);
signal s4_3 : unsigned(31 downto 0);
signal s5_1 : unsigned(31 downto 0);
signal s5_2 : unsigned(31 downto 0);
signal s5_3 : unsigned(31 downto 0);
signal s6_1 : unsigned(31 downto 0);
signal s6_2 : unsigned(31 downto 0);
signal s6_3 : unsigned(31 downto 0);
signal s7_1 : unsigned(31 downto 0);
signal s7_2 : unsigned(31 downto 0);
signal s7_3 : unsigned(31 downto 0);
signal s8_1 : unsigned(31 downto 0);
signal s8_2 : unsigned(31 downto 0);
signal s8_3 : unsigned(31 downto 0);
component cf_cordic_v_32_32_32_49 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_49;
component cf_cordic_v_32_32_32_36 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_36;
component cf_cordic_v_32_32_32_34 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_34;
component cf_cordic_v_32_32_32_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_32;
component cf_cordic_v_32_32_32_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_30;
component cf_cordic_v_32_32_32_29 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_29;
component cf_cordic_v_32_32_32_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_28;
component cf_cordic_v_32_32_32_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_27;
begin
s1 : cf_cordic_v_32_32_32_49 port map (clock_c, i1, i2, s3_1, s3_2, s3_3, s1_1, s1_2, s1_3);
s2 : cf_cordic_v_32_32_32_36 port map (clock_c, i1, i2, s1_1, s1_2, s1_3, s2_1, s2_2, s2_3);
s3 : cf_cordic_v_32_32_32_34 port map (clock_c, i1, i2, s4_1, s4_2, s4_3, s3_1, s3_2, s3_3);
s4 : cf_cordic_v_32_32_32_32 port map (clock_c, i1, i2, s5_1, s5_2, s5_3, s4_1, s4_2, s4_3);
s5 : cf_cordic_v_32_32_32_30 port map (clock_c, i1, i2, s6_1, s6_2, s6_3, s5_1, s5_2, s5_3);
s6 : cf_cordic_v_32_32_32_29 port map (clock_c, i1, i2, s7_1, s7_2, s7_3, s6_1, s6_2, s6_3);
s7 : cf_cordic_v_32_32_32_28 port map (clock_c, i1, i2, s8_1, s8_2, s8_3, s7_1, s7_2, s7_3);
s8 : cf_cordic_v_32_32_32_27 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_25 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_25;
architecture rtl of cf_cordic_v_32_32_32_25 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(12 downto 0);
signal n6 : unsigned(13 downto 0);
signal n7 : unsigned(14 downto 0);
signal n8 : unsigned(16 downto 0);
signal n9 : unsigned(31 downto 0);
signal s10_1 : unsigned(8 downto 0);
component cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_v_32_32_32_54;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s10_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= n1 & n6;
n8 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15);
n9 <= n7 & n8;
s10 : cf_cordic_v_32_32_32_54 port map (n1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_24 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_24;
architecture rtl of cf_cordic_v_32_32_32_24 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_25 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_25;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000000101000101111101";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_25 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_25 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_23 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_23;
architecture rtl of cf_cordic_v_32_32_32_23 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(12 downto 0);
signal n6 : unsigned(13 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(31 downto 0);
signal s9_1 : unsigned(8 downto 0);
component cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_v_32_32_32_54;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s9_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14);
n8 <= n6 & n7;
s9 : cf_cordic_v_32_32_32_54 port map (n1, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_22;
architecture rtl of cf_cordic_v_32_32_32_22 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_23 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_23;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000001010001011111010";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_23 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_23 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_21 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_21;
architecture rtl of cf_cordic_v_32_32_32_21 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(12 downto 0);
signal n6 : unsigned(18 downto 0);
signal n7 : unsigned(31 downto 0);
signal s8_1 : unsigned(8 downto 0);
component cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_v_32_32_32_54;
begin
n1 <= i1(31 downto 31);
n2 <= n1 & s8_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13);
n7 <= n5 & n6;
s8 : cf_cordic_v_32_32_32_54 port map (n1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_20;
architecture rtl of cf_cordic_v_32_32_32_20 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_21 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_21;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000000000010100010111110011";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_21 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_21 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_19;
architecture rtl of cf_cordic_v_32_32_32_19 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(19 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0);
signal n10 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(9 downto 0);
signal n14 : unsigned(10 downto 0);
signal n15 : unsigned(11 downto 0);
signal n16 : unsigned(19 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s27_1 : unsigned(8 downto 0);
signal s28_1 : unsigned(8 downto 0);
signal s29_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_v_32_32_32_54;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s27_1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12);
n6 <= n4 & n5;
n7 <= i3 + n6;
n8 <= i3 - n6;
n9 <= n7 when s29_1 = "1" else n8;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n10 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
n11 <= not s29_1;
n12 <= i3(31 downto 31);
n13 <= n12 & s28_1;
n14 <= n12 & n13;
n15 <= n12 & n14;
n16 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12);
n17 <= n15 & n16;
n18 <= i4 + n17;
n19 <= i4 - n17;
n20 <= n18 when n11 = "1" else n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n21 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= "00000000000000101000101111100110";
n23 <= i5 + n22;
n24 <= i5 - n22;
n25 <= n23 when s29_1 = "1" else n24;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n26 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n26 <= n25;
    end if;
  end if;
end process;
s27 : cf_cordic_v_32_32_32_54 port map (n1, s27_1);
s28 : cf_cordic_v_32_32_32_54 port map (n12, s28_1);
s29 : cf_cordic_v_32_32_32_56 port map (i4, s29_1);
o3 <= n26;
o2 <= n21;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_18;
architecture rtl of cf_cordic_v_32_32_32_18 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(10 downto 0);
signal n4 : unsigned(20 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(9 downto 0);
signal n13 : unsigned(10 downto 0);
signal n14 : unsigned(20 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s25_1 : unsigned(8 downto 0);
signal s26_1 : unsigned(8 downto 0);
signal s27_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_v_32_32_32_54;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s25_1;
n3 <= n1 & n2;
n4 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11);
n5 <= n3 & n4;
n6 <= i3 + n5;
n7 <= i3 - n5;
n8 <= n6 when s27_1 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= not s27_1;
n11 <= i3(31 downto 31);
n12 <= n11 & s26_1;
n13 <= n11 & n12;
n14 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11);
n15 <= n13 & n14;
n16 <= i4 + n15;
n17 <= i4 - n15;
n18 <= n16 when n10 = "1" else n17;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n19 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= "00000000000001010001011111001100";
n21 <= i5 + n20;
n22 <= i5 - n20;
n23 <= n21 when s27_1 = "1" else n22;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n24 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
s25 : cf_cordic_v_32_32_32_54 port map (n1, s25_1);
s26 : cf_cordic_v_32_32_32_54 port map (n11, s26_1);
s27 : cf_cordic_v_32_32_32_56 port map (i4, s27_1);
o3 <= n24;
o2 <= n19;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_17;
architecture rtl of cf_cordic_v_32_32_32_17 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(21 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(9 downto 0);
signal n12 : unsigned(21 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s23_1 : unsigned(8 downto 0);
signal s24_1 : unsigned(8 downto 0);
signal s25_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_54 is
port (
i1 : in  unsigned(0 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_cordic_v_32_32_32_54;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & s23_1;
n3 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10);
n4 <= n2 & n3;
n5 <= i3 + n4;
n6 <= i3 - n4;
n7 <= n5 when s25_1 = "1" else n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n8 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
n9 <= not s25_1;
n10 <= i3(31 downto 31);
n11 <= n10 & s24_1;
n12 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10);
n13 <= n11 & n12;
n14 <= i4 + n13;
n15 <= i4 - n13;
n16 <= n14 when n9 = "1" else n15;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n17 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n17 <= n16;
    end if;
  end if;
end process;
n18 <= "00000000000010100010111110011000";
n19 <= i5 + n18;
n20 <= i5 - n18;
n21 <= n19 when s25_1 = "1" else n20;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n22 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n22 <= n21;
    end if;
  end if;
end process;
s23 : cf_cordic_v_32_32_32_54 port map (n1, s23_1);
s24 : cf_cordic_v_32_32_32_54 port map (n10, s24_1);
s25 : cf_cordic_v_32_32_32_56 port map (i4, s25_1);
o3 <= n22;
o2 <= n17;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_16;
architecture rtl of cf_cordic_v_32_32_32_16 is
signal s1_1 : unsigned(31 downto 0);
signal s1_2 : unsigned(31 downto 0);
signal s1_3 : unsigned(31 downto 0);
signal s2_1 : unsigned(31 downto 0);
signal s2_2 : unsigned(31 downto 0);
signal s2_3 : unsigned(31 downto 0);
signal s3_1 : unsigned(31 downto 0);
signal s3_2 : unsigned(31 downto 0);
signal s3_3 : unsigned(31 downto 0);
signal s4_1 : unsigned(31 downto 0);
signal s4_2 : unsigned(31 downto 0);
signal s4_3 : unsigned(31 downto 0);
signal s5_1 : unsigned(31 downto 0);
signal s5_2 : unsigned(31 downto 0);
signal s5_3 : unsigned(31 downto 0);
signal s6_1 : unsigned(31 downto 0);
signal s6_2 : unsigned(31 downto 0);
signal s6_3 : unsigned(31 downto 0);
signal s7_1 : unsigned(31 downto 0);
signal s7_2 : unsigned(31 downto 0);
signal s7_3 : unsigned(31 downto 0);
signal s8_1 : unsigned(31 downto 0);
signal s8_2 : unsigned(31 downto 0);
signal s8_3 : unsigned(31 downto 0);
component cf_cordic_v_32_32_32_51 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_51;
component cf_cordic_v_32_32_32_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_26;
component cf_cordic_v_32_32_32_24 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_24;
component cf_cordic_v_32_32_32_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_22;
component cf_cordic_v_32_32_32_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_20;
component cf_cordic_v_32_32_32_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_19;
component cf_cordic_v_32_32_32_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_18;
component cf_cordic_v_32_32_32_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_17;
begin
s1 : cf_cordic_v_32_32_32_51 port map (clock_c, i1, i2, s3_1, s3_2, s3_3, s1_1, s1_2, s1_3);
s2 : cf_cordic_v_32_32_32_26 port map (clock_c, i1, i2, s1_1, s1_2, s1_3, s2_1, s2_2, s2_3);
s3 : cf_cordic_v_32_32_32_24 port map (clock_c, i1, i2, s4_1, s4_2, s4_3, s3_1, s3_2, s3_3);
s4 : cf_cordic_v_32_32_32_22 port map (clock_c, i1, i2, s5_1, s5_2, s5_3, s4_1, s4_2, s4_3);
s5 : cf_cordic_v_32_32_32_20 port map (clock_c, i1, i2, s6_1, s6_2, s6_3, s5_1, s5_2, s5_3);
s6 : cf_cordic_v_32_32_32_19 port map (clock_c, i1, i2, s7_1, s7_2, s7_3, s6_1, s6_2, s6_3);
s7 : cf_cordic_v_32_32_32_18 port map (clock_c, i1, i2, s8_1, s8_2, s8_3, s7_1, s7_2, s7_3);
s8 : cf_cordic_v_32_32_32_17 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_15 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_15;
architecture rtl of cf_cordic_v_32_32_32_15 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(6 downto 0);
signal n8 : unsigned(7 downto 0);
signal n9 : unsigned(23 downto 0);
signal n10 : unsigned(31 downto 0);
begin
n1 <= i1(31 downto 31);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= n1 & n6;
n8 <= n1 & n7;
n9 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8);
n10 <= n8 & n9;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_14;
architecture rtl of cf_cordic_v_32_32_32_14 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_15 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_15;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000001010001011111001010011";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_15 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_15 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_13 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_13;
architecture rtl of cf_cordic_v_32_32_32_13 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(6 downto 0);
signal n8 : unsigned(24 downto 0);
signal n9 : unsigned(31 downto 0);
begin
n1 <= i1(31 downto 31);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= n1 & n6;
n8 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7);
n9 <= n7 & n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_12;
architecture rtl of cf_cordic_v_32_32_32_12 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_13 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_13;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000010100010111110001010101";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_13 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_13 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_11 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_11;
architecture rtl of cf_cordic_v_32_32_32_11 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(25 downto 0);
signal n8 : unsigned(31 downto 0);
begin
n1 <= i1(31 downto 31);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= n1 & n5;
n7 <= i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6);
n8 <= n6 & n7;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_10;
architecture rtl of cf_cordic_v_32_32_32_10 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s15_1 : unsigned(31 downto 0);
signal s16_1 : unsigned(31 downto 0);
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_11 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_11;
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i3 + s16_1;
n2 <= i3 - s16_1;
n3 <= n1 when s17_1 = "1" else n2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
n5 <= not s17_1;
n6 <= i4 + s15_1;
n7 <= i4 - s15_1;
n8 <= n6 when n5 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= "00000000101000101111011000011110";
n11 <= i5 + n10;
n12 <= i5 - n10;
n13 <= n11 when s17_1 = "1" else n12;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n14 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
s15 : cf_cordic_v_32_32_32_11 port map (i3, s15_1);
s16 : cf_cordic_v_32_32_32_11 port map (i4, s16_1);
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n14;
o2 <= n9;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_9;
architecture rtl of cf_cordic_v_32_32_32_9 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(26 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0);
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(1 downto 0);
signal n15 : unsigned(2 downto 0);
signal n16 : unsigned(3 downto 0);
signal n17 : unsigned(4 downto 0);
signal n18 : unsigned(26 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n24 : unsigned(31 downto 0);
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(31 downto 0);
signal n27 : unsigned(31 downto 0);
signal n28 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s29_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= n1 & n4;
n6 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5);
n7 <= n5 & n6;
n8 <= i3 + n7;
n9 <= i3 - n7;
n10 <= n8 when s29_1 = "1" else n9;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n11 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= not s29_1;
n13 <= i3(31 downto 31);
n14 <= n13 & n13;
n15 <= n13 & n14;
n16 <= n13 & n15;
n17 <= n13 & n16;
n18 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5);
n19 <= n17 & n18;
n20 <= i4 + n19;
n21 <= i4 - n19;
n22 <= n20 when n12 = "1" else n21;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n23 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n23 <= n22;
    end if;
  end if;
end process;
n24 <= "00000001010001011101011111100001";
n25 <= i5 + n24;
n26 <= i5 - n24;
n27 <= n25 when s29_1 = "1" else n26;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n28 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n28 <= n27;
    end if;
  end if;
end process;
s29 : cf_cordic_v_32_32_32_56 port map (i4, s29_1);
o3 <= n28;
o2 <= n23;
o1 <= n11;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_8;
architecture rtl of cf_cordic_v_32_32_32_8 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(27 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0);
signal n10 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(1 downto 0);
signal n14 : unsigned(2 downto 0);
signal n15 : unsigned(3 downto 0);
signal n16 : unsigned(27 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s27_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= n1 & n3;
n5 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4);
n6 <= n4 & n5;
n7 <= i3 + n6;
n8 <= i3 - n6;
n9 <= n7 when s27_1 = "1" else n8;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n10 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
n11 <= not s27_1;
n12 <= i3(31 downto 31);
n13 <= n12 & n12;
n14 <= n12 & n13;
n15 <= n12 & n14;
n16 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4);
n17 <= n15 & n16;
n18 <= i4 + n17;
n19 <= i4 - n17;
n20 <= n18 when n11 = "1" else n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n21 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= "00000010100010110000110101000011";
n23 <= i5 + n22;
n24 <= i5 - n22;
n25 <= n23 when s27_1 = "1" else n24;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n26 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n26 <= n25;
    end if;
  end if;
end process;
s27 : cf_cordic_v_32_32_32_56 port map (i4, s27_1);
o3 <= n26;
o2 <= n21;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_7;
architecture rtl of cf_cordic_v_32_32_32_7 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(28 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(1 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(28 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s25_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= n1 & n1;
n3 <= n1 & n2;
n4 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3);
n5 <= n3 & n4;
n6 <= i3 + n5;
n7 <= i3 - n5;
n8 <= n6 when s25_1 = "1" else n7;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= not s25_1;
n11 <= i3(31 downto 31);
n12 <= n11 & n11;
n13 <= n11 & n12;
n14 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3);
n15 <= n13 & n14;
n16 <= i4 + n15;
n17 <= i4 - n15;
n18 <= n16 when n10 = "1" else n17;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n19 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= "00000101000100010001000111010100";
n21 <= i5 + n20;
n22 <= i5 - n20;
n23 <= n21 when s25_1 = "1" else n22;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n24 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
s25 : cf_cordic_v_32_32_32_56 port map (i4, s25_1);
o3 <= n24;
o2 <= n19;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_6;
architecture rtl of cf_cordic_v_32_32_32_6 is
signal s1_1 : unsigned(31 downto 0);
signal s1_2 : unsigned(31 downto 0);
signal s1_3 : unsigned(31 downto 0);
signal s2_1 : unsigned(31 downto 0);
signal s2_2 : unsigned(31 downto 0);
signal s2_3 : unsigned(31 downto 0);
signal s3_1 : unsigned(31 downto 0);
signal s3_2 : unsigned(31 downto 0);
signal s3_3 : unsigned(31 downto 0);
signal s4_1 : unsigned(31 downto 0);
signal s4_2 : unsigned(31 downto 0);
signal s4_3 : unsigned(31 downto 0);
signal s5_1 : unsigned(31 downto 0);
signal s5_2 : unsigned(31 downto 0);
signal s5_3 : unsigned(31 downto 0);
signal s6_1 : unsigned(31 downto 0);
signal s6_2 : unsigned(31 downto 0);
signal s6_3 : unsigned(31 downto 0);
signal s7_1 : unsigned(31 downto 0);
signal s7_2 : unsigned(31 downto 0);
signal s7_3 : unsigned(31 downto 0);
signal s8_1 : unsigned(31 downto 0);
signal s8_2 : unsigned(31 downto 0);
signal s8_3 : unsigned(31 downto 0);
component cf_cordic_v_32_32_32_53 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_53;
component cf_cordic_v_32_32_32_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_16;
component cf_cordic_v_32_32_32_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_14;
component cf_cordic_v_32_32_32_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_12;
component cf_cordic_v_32_32_32_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_10;
component cf_cordic_v_32_32_32_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_9;
component cf_cordic_v_32_32_32_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_8;
component cf_cordic_v_32_32_32_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_7;
begin
s1 : cf_cordic_v_32_32_32_53 port map (clock_c, i1, i2, s3_1, s3_2, s3_3, s1_1, s1_2, s1_3);
s2 : cf_cordic_v_32_32_32_16 port map (clock_c, i1, i2, s1_1, s1_2, s1_3, s2_1, s2_2, s2_3);
s3 : cf_cordic_v_32_32_32_14 port map (clock_c, i1, i2, s4_1, s4_2, s4_3, s3_1, s3_2, s3_3);
s4 : cf_cordic_v_32_32_32_12 port map (clock_c, i1, i2, s5_1, s5_2, s5_3, s4_1, s4_2, s4_3);
s5 : cf_cordic_v_32_32_32_10 port map (clock_c, i1, i2, s6_1, s6_2, s6_3, s5_1, s5_2, s5_3);
s6 : cf_cordic_v_32_32_32_9 port map (clock_c, i1, i2, s7_1, s7_2, s7_3, s6_1, s6_2, s6_3);
s7 : cf_cordic_v_32_32_32_8 port map (clock_c, i1, i2, s8_1, s8_2, s8_3, s7_1, s7_2, s7_3);
s8 : cf_cordic_v_32_32_32_7 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_5;
architecture rtl of cf_cordic_v_32_32_32_5 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(30 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(30 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n16 : unsigned(31 downto 0);
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(31 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s21_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31);
n2 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3) &
  i4(2 downto 2) &
  i4(1 downto 1);
n3 <= n1 & n2;
n4 <= i3 + n3;
n5 <= i3 - n3;
n6 <= n4 when s21_1 = "1" else n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= not s21_1;
n9 <= i3(31 downto 31);
n10 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1);
n11 <= n9 & n10;
n12 <= i4 + n11;
n13 <= i4 - n11;
n14 <= n12 when n8 = "1" else n13;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n15 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
n16 <= "00010010111001000000010100011110";
n17 <= i5 + n16;
n18 <= i5 - n16;
n19 <= n17 when s21_1 = "1" else n18;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n20 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n20 <= n19;
    end if;
  end if;
end process;
s21 : cf_cordic_v_32_32_32_56 port map (i4, s21_1);
o3 <= n20;
o2 <= n15;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_4;
architecture rtl of cf_cordic_v_32_32_32_4 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0);
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(31 downto 0);
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(31 downto 0);
signal n16 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s17_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_56 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_56;
begin
n1 <= i4(31 downto 31) &
  i4(30 downto 30) &
  i4(29 downto 29) &
  i4(28 downto 28) &
  i4(27 downto 27) &
  i4(26 downto 26) &
  i4(25 downto 25) &
  i4(24 downto 24) &
  i4(23 downto 23) &
  i4(22 downto 22) &
  i4(21 downto 21) &
  i4(20 downto 20) &
  i4(19 downto 19) &
  i4(18 downto 18) &
  i4(17 downto 17) &
  i4(16 downto 16) &
  i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3) &
  i4(2 downto 2) &
  i4(1 downto 1) &
  i4(0 downto 0);
n2 <= i3 + n1;
n3 <= i3 - n1;
n4 <= n2 when s17_1 = "1" else n3;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n5 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
n6 <= not s17_1;
n7 <= i3(31 downto 31) &
  i3(30 downto 30) &
  i3(29 downto 29) &
  i3(28 downto 28) &
  i3(27 downto 27) &
  i3(26 downto 26) &
  i3(25 downto 25) &
  i3(24 downto 24) &
  i3(23 downto 23) &
  i3(22 downto 22) &
  i3(21 downto 21) &
  i3(20 downto 20) &
  i3(19 downto 19) &
  i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= i4 + n7;
n9 <= i4 - n7;
n10 <= n8 when n6 = "1" else n9;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n11 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= "00100000000000000000000000000000";
n13 <= i5 + n12;
n14 <= i5 - n12;
n15 <= n13 when s17_1 = "1" else n14;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n16 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
s17 : cf_cordic_v_32_32_32_56 port map (i4, s17_1);
o3 <= n16;
o2 <= n11;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_3;
architecture rtl of cf_cordic_v_32_32_32_3 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(31 downto 0);
signal n6 : unsigned(31 downto 0);
signal n7 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(31 downto 0);
begin
n1 <= "00000000000000000000000000000000";
n2 <= n1 - i3;
n3 <= "00000000000000000000000000000000";
n4 <= n3 - i4;
n5 <= i5 - n12;
n6 <= n2 when i6 = "1" else i3;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n7 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n7 <= n6;
    end if;
  end if;
end process;
n8 <= n4 when i6 = "1" else i4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n9 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
n10 <= n5 when i6 = "1" else i5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n11 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= "10000000000000000000000000000000";
o3 <= n11;
o2 <= n9;
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_2 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_cordic_v_32_32_32_2;
architecture rtl of cf_cordic_v_32_32_32_2 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(30 downto 0);
signal n4 : unsigned(31 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(32 downto 0);
signal n7 : unsigned(32 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(32 downto 0);
begin
n1 <= i1(31 downto 31);
n2 <= not n1;
n3 <= i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n4 <= n2 & n3;
n5 <= "0";
n6 <= n5 & n4;
n7 <= n6 - n9;
n8 <= n7(32 downto 32);
n9 <= "010000000000000000000000000000000";
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32_1;
architecture rtl of cf_cordic_v_32_32_32_1 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n3 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal s4_1 : unsigned(31 downto 0);
signal s4_2 : unsigned(31 downto 0);
signal s4_3 : unsigned(31 downto 0);
signal s5_1 : unsigned(31 downto 0);
signal s5_2 : unsigned(31 downto 0);
signal s5_3 : unsigned(31 downto 0);
signal s6_1 : unsigned(31 downto 0);
signal s6_2 : unsigned(31 downto 0);
signal s6_3 : unsigned(31 downto 0);
signal s7_1 : unsigned(31 downto 0);
signal s7_2 : unsigned(31 downto 0);
signal s7_3 : unsigned(31 downto 0);
signal s8_1 : unsigned(31 downto 0);
signal s8_2 : unsigned(31 downto 0);
signal s8_3 : unsigned(31 downto 0);
signal s9_1 : unsigned(0 downto 0);
component cf_cordic_v_32_32_32_55 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_55;
component cf_cordic_v_32_32_32_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_6;
component cf_cordic_v_32_32_32_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_5;
component cf_cordic_v_32_32_32_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_4;
component cf_cordic_v_32_32_32_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_3;
component cf_cordic_v_32_32_32_2 is
port (
i1 : in  unsigned(31 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_cordic_v_32_32_32_2;
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n1 <= i3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n2 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n2 <= i4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i2 = "1" then
      n3 <= "00000000000000000000000000000000";
    elsif i1 = "1" then
      n3 <= i5;
    end if;
  end if;
end process;
s4 : cf_cordic_v_32_32_32_55 port map (clock_c, i1, i2, s6_1, s6_2, s6_3, s4_1, s4_2, s4_3);
s5 : cf_cordic_v_32_32_32_6 port map (clock_c, i1, i2, s4_1, s4_2, s4_3, s5_1, s5_2, s5_3);
s6 : cf_cordic_v_32_32_32_5 port map (clock_c, i1, i2, s7_1, s7_2, s7_3, s6_1, s6_2, s6_3);
s7 : cf_cordic_v_32_32_32_4 port map (clock_c, i1, i2, s8_1, s8_2, s8_3, s7_1, s7_2, s7_3);
s8 : cf_cordic_v_32_32_32_3 port map (clock_c, i1, i2, n1, n2, n3, s9_1, s8_1, s8_2, s8_3);
s9 : cf_cordic_v_32_32_32_2 port map (n1, s9_1);
o3 <= s5_3;
o2 <= s5_2;
o1 <= s5_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_cordic_v_32_32_32 is
port(
signal clock_c : in std_logic;
signal enable_i : in unsigned(0 downto 0);
signal reset_i : in unsigned(0 downto 0);
signal real_i : in unsigned(31 downto 0);
signal imag_i : in unsigned(31 downto 0);
signal ang_i : in unsigned(31 downto 0);
signal real_o : out unsigned(31 downto 0);
signal imag_o : out unsigned(31 downto 0);
signal ang_o : out unsigned(31 downto 0));
end entity cf_cordic_v_32_32_32;
architecture rtl of cf_cordic_v_32_32_32 is
component cf_cordic_v_32_32_32_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(31 downto 0);
i5 : in  unsigned(31 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_cordic_v_32_32_32_1;
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
begin
s1 : cf_cordic_v_32_32_32_1 port map (clock_c, enable_i, reset_i, real_i, imag_i, ang_i, n1, n2, n3);
real_o <= n1;
imag_o <= n2;
ang_o <= n3;
end architecture rtl;


